library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;
library work;

package config is

  -- LLR bit-widths
  constant QLLR : integer := 3;
  constant QCh : integer := 4;

  -- Variable node degree
  constant VNodeDegree : integer := 5;

  -- Channel LLR
  subtype ChLLRType is integer range 0 to 2**QCh-1;

  -- Internal LLR
  subtype IntLLRSubType is integer range 0 to 2**QLLR-1;
  type IntLLRType is array (0 to VNodeDegree-1) of IntLLRSubType;
  
  -- LUT definition
  constant LUTSize : integer := 2**(QCh + (VNodeDegree-1)*QLLR);  
  type LUTType is array (0 to LUTSize-1) of integer range 0 to 2**QLLR-1;
  -- LUT for VNodeDegree 3
  --constant LUT : LUTType := (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,0,0,0,0,0,0,0,0,0,1,1,1,1,1,2,2,0,0,0,0,0,0,1,1,1,1,1,1,1,2,2,3,0,0,0,1,1,1,1,1,1,2,2,2,2,3,4,5,1,1,2,2,2,3,3,3,4,4,4,5,5,5,6,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,0,0,0,0,0,0,1,1,1,1,1,1,1,2,2,3,0,0,0,0,1,1,1,1,1,1,1,2,2,2,3,4,0,0,1,1,1,1,1,1,2,2,2,2,3,3,4,5,0,1,1,1,1,2,2,2,2,3,3,3,4,4,5,6,1,1,2,2,2,3,3,3,4,4,4,5,5,5,6,6,2,3,4,5,5,5,5,6,6,6,6,6,6,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,1,1,1,1,1,1,1,2,2,3,0,0,0,1,1,1,1,1,1,2,2,2,2,3,4,5,0,1,1,1,1,1,2,2,2,2,2,3,3,4,4,5,0,1,1,1,2,2,2,2,3,3,3,4,4,5,5,6,1,1,2,2,2,3,3,3,4,4,4,5,5,5,6,6,1,2,3,3,4,4,4,5,5,5,5,6,6,6,6,7,4,5,5,6,6,6,6,6,6,6,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,0,0,0,0,1,1,1,1,1,1,1,2,2,2,3,4,0,1,1,1,1,1,2,2,2,2,2,3,3,4,4,5,0,1,1,1,2,2,2,2,3,3,3,4,4,5,5,6,1,1,2,2,2,3,3,3,4,4,4,5,5,5,6,6,1,2,2,3,3,4,4,4,5,5,5,5,6,6,6,7,2,3,4,4,5,5,5,5,6,6,6,6,6,6,7,7,5,5,6,6,6,6,6,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,1,1,1,1,1,2,2,0,0,1,1,1,1,1,1,2,2,2,2,3,3,4,5,0,1,1,1,2,2,2,2,3,3,3,4,4,5,5,6,1,1,2,2,2,3,3,3,4,4,4,5,5,5,6,6,1,2,2,3,3,4,4,4,5,5,5,5,6,6,6,7,2,3,3,4,4,5,5,5,5,5,6,6,6,6,6,7,3,4,5,5,5,6,6,6,6,6,6,6,7,7,7,7,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,1,1,1,1,1,1,1,2,2,3,0,1,1,1,1,2,2,2,2,3,3,3,4,4,5,6,1,1,2,2,2,3,3,3,4,4,4,5,5,5,6,6,1,2,2,3,3,4,4,4,5,5,5,5,6,6,6,7,2,3,3,4,4,5,5,5,5,5,6,6,6,6,6,7,2,3,4,5,5,5,5,6,6,6,6,6,6,7,7,7,4,5,5,6,6,6,6,6,6,6,7,7,7,7,7,7,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,1,1,1,1,1,1,2,2,2,2,3,4,5,1,1,2,2,2,3,3,3,4,4,4,5,5,5,6,6,1,2,3,3,4,4,4,5,5,5,5,6,6,6,6,7,2,3,4,4,5,5,5,5,6,6,6,6,6,6,7,7,3,4,5,5,5,6,6,6,6,6,6,6,7,7,7,7,4,5,5,6,6,6,6,6,6,6,7,7,7,7,7,7,5,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,1,2,2,2,3,3,3,4,4,4,5,5,5,6,6,2,3,4,5,5,5,5,6,6,6,6,6,6,7,7,7,4,5,5,6,6,6,6,6,6,6,7,7,7,7,7,7,5,5,6,6,6,6,6,7,7,7,7,7,7,7,7,7,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7);
  -- LUT for VNodeDegree 4
  --constant LUT : LUTType := (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,3,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,0,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,4,4,5,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,1,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,3,3,3,4,5,5,6,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,6,0,0,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,6,0,0,0,0,1,1,1,1,2,2,3,3,4,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,7,7,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,6,0,0,0,0,1,1,1,1,2,2,3,3,4,4,5,6,0,0,0,1,1,1,2,2,2,3,3,4,4,5,6,7,0,1,1,1,2,2,3,3,4,4,4,5,5,6,6,7,0,1,2,2,3,4,4,4,5,5,6,6,6,6,7,7,0,0,0,0,0,0,0,0,0,0,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,1,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,1,2,2,3,3,4,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,3,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,4,4,5,6,0,0,1,1,1,1,2,2,3,3,3,4,5,5,6,7,0,0,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,7,7,0,1,2,2,3,4,4,4,5,5,6,6,6,6,7,7,1,2,3,3,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,4,4,5,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,5,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,0,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,4,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,0,1,1,1,2,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,4,4,5,6,0,0,1,1,1,1,2,2,3,3,3,4,5,5,6,7,0,1,1,2,2,3,3,3,4,4,5,5,6,6,6,7,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,6,0,0,0,0,1,1,1,1,2,2,2,3,4,4,5,6,0,0,0,1,1,1,2,2,2,3,3,4,4,5,6,7,0,0,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,4,4,5,6,0,0,0,1,1,1,2,2,2,3,3,4,4,5,6,7,0,0,1,1,1,2,2,3,3,3,4,4,5,6,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,7,7,1,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,5,0,0,0,0,0,0,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,4,4,5,6,0,0,0,1,1,1,2,2,2,3,3,4,4,5,6,7,0,0,1,1,1,2,2,3,3,3,4,4,5,6,6,7,0,1,1,2,2,3,3,3,4,4,5,5,6,6,6,7,0,1,2,2,3,4,4,4,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,6,6,6,6,6,7,7,7,7,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,4,4,5,6,0,0,1,1,1,1,2,2,3,3,3,4,5,5,6,7,0,0,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,7,7,0,1,2,2,3,4,4,4,5,5,6,6,6,6,7,7,1,2,3,3,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,4,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,3,4,4,5,5,6,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,6,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,1,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,3,3,3,4,5,5,6,7,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,0,1,1,1,2,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,4,4,5,6,0,0,1,1,1,1,2,2,3,3,3,4,5,5,6,7,0,1,1,2,2,3,3,3,4,4,5,5,6,6,6,7,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,1,1,1,2,2,3,5,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,6,0,0,0,0,0,1,1,1,1,2,2,3,3,4,5,6,0,0,0,0,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,1,2,2,3,3,3,4,5,5,6,7,0,1,1,1,2,2,3,3,4,4,4,5,5,6,6,7,0,1,2,3,3,4,4,5,5,5,6,6,6,7,7,7,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,1,2,2,3,3,3,4,5,5,6,7,0,0,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,1,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,3,3,4,4,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,1,2,2,3,3,3,4,5,5,6,7,0,0,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,7,7,0,1,2,3,3,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,4,4,5,6,0,0,1,1,1,1,2,2,3,3,3,4,5,5,6,7,0,0,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,7,7,0,1,2,2,3,4,4,4,5,5,6,6,6,6,7,7,1,2,3,3,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,0,0,0,0,1,1,1,1,1,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,3,3,3,4,5,5,6,7,0,1,1,1,2,2,3,3,4,4,4,5,5,6,6,7,0,1,1,2,3,3,4,4,4,5,5,6,6,6,7,7,0,1,2,3,3,4,4,5,5,5,6,6,6,7,7,7,1,2,3,3,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,7,7,7,7,7,7,2,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,0,0,1,1,1,1,2,2,3,3,3,4,5,5,6,7,0,1,1,2,2,3,3,3,4,4,5,5,6,6,6,7,0,1,2,3,3,4,4,5,5,5,6,6,6,7,7,7,1,2,3,3,4,4,5,5,6,6,6,6,7,7,7,7,1,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,6,0,0,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,6,0,0,0,0,1,1,1,1,2,2,2,3,4,4,5,6,0,0,0,1,1,1,2,2,2,3,3,4,4,5,6,7,0,0,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,1,2,2,3,3,3,4,5,5,6,7,0,0,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,1,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,3,3,4,4,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,0,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,7,7,0,1,2,3,3,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,4,4,5,6,0,0,1,1,1,1,2,2,3,3,3,4,5,5,6,7,0,0,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,7,7,0,1,2,2,3,4,4,4,5,5,6,6,6,6,7,7,1,2,3,3,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,4,4,5,6,7,0,0,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,7,7,0,1,2,2,3,4,4,4,5,5,6,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,6,0,0,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,1,2,3,3,4,4,4,5,5,6,6,6,7,7,0,1,2,3,3,4,4,5,5,5,6,6,6,7,7,7,1,2,3,3,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,0,0,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,3,4,4,5,5,6,6,6,6,7,7,7,7,1,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,6,0,0,0,0,1,1,1,1,2,2,3,3,4,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,7,7,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,4,4,5,6,0,0,0,1,1,1,2,2,2,3,3,4,4,5,6,7,0,0,1,1,1,2,2,3,3,3,4,4,5,6,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,7,7,1,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,1,2,2,3,3,3,4,5,5,6,7,0,0,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,7,7,0,1,2,3,3,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,4,4,5,6,0,0,1,1,1,1,2,2,3,3,3,4,5,5,6,7,0,0,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,7,7,0,1,2,2,3,4,4,4,5,5,6,6,6,6,7,7,1,2,3,3,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,4,4,5,6,7,0,0,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,7,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,3,3,4,4,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,6,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,7,7,0,1,2,2,3,4,4,4,5,5,6,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,7,7,0,1,2,3,3,4,4,5,5,5,6,6,6,7,7,7,1,2,3,3,4,5,5,5,6,6,6,6,7,7,7,7,1,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,7,7,1,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,6,0,0,0,0,1,1,1,1,2,2,3,3,4,4,5,6,0,0,0,1,1,1,2,2,2,3,3,4,4,5,6,7,0,1,1,1,2,2,3,3,4,4,4,5,5,6,6,7,0,1,2,2,3,4,4,4,5,5,6,6,6,6,7,7,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,5,0,0,0,0,0,0,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,4,4,5,6,0,0,0,1,1,1,2,2,2,3,3,4,4,5,6,7,0,0,1,1,1,2,2,3,3,3,4,4,5,6,6,7,0,1,1,2,2,3,3,3,4,4,5,5,6,6,6,7,0,1,2,2,3,4,4,4,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,6,6,6,6,6,7,7,7,7,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,4,4,5,6,0,0,1,1,1,1,2,2,3,3,3,4,5,5,6,7,0,0,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,7,7,0,1,2,2,3,4,4,4,5,5,6,6,6,6,7,7,1,2,3,3,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,4,4,5,6,7,0,0,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,7,7,0,1,2,2,3,4,4,4,5,5,6,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,3,3,4,4,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,6,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,7,7,0,1,2,2,3,4,4,4,5,5,6,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,0,0,0,1,1,1,2,2,2,3,3,4,4,5,6,7,0,1,1,2,2,3,3,3,4,4,5,5,6,6,6,7,0,1,2,2,3,4,4,4,5,5,6,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,7,7,7,7,1,2,3,4,4,5,5,6,6,6,6,7,7,7,7,7,1,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,2,4,5,5,6,6,6,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,0,1,1,1,2,2,3,3,4,4,4,5,5,6,6,7,0,1,2,2,3,4,4,4,5,5,6,6,6,6,7,7,1,2,3,3,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,5,6,6,6,7,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,0,1,2,2,3,4,4,4,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,6,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,1,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,1,2,2,3,3,4,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,3,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,4,4,5,6,0,0,1,1,1,1,2,2,3,3,3,4,5,5,6,7,0,0,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,7,7,0,1,2,2,3,4,4,4,5,5,6,6,6,6,7,7,1,2,3,3,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,0,0,0,0,1,1,1,1,1,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,3,3,3,4,5,5,6,7,0,1,1,1,2,2,3,3,4,4,4,5,5,6,6,7,0,1,1,2,3,3,4,4,4,5,5,6,6,6,7,7,0,1,2,3,3,4,4,5,5,5,6,6,6,7,7,7,1,2,3,3,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,7,7,7,7,7,7,2,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,6,0,0,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,1,2,3,3,4,4,4,5,5,6,6,6,7,7,0,1,2,3,3,4,4,5,5,5,6,6,6,7,7,7,1,2,3,3,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,7,7,0,1,2,3,3,4,4,5,5,5,6,6,6,7,7,7,1,2,3,3,4,5,5,5,6,6,6,6,7,7,7,7,1,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,0,1,1,1,2,2,3,3,4,4,4,5,5,6,6,7,0,1,2,2,3,4,4,4,5,5,6,6,6,6,7,7,1,2,3,3,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,5,6,6,6,7,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,3,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,7,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,2,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,2,3,3,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,4,4,5,6,0,0,1,1,1,1,2,2,3,3,3,4,5,5,6,7,0,0,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,7,7,0,1,2,2,3,4,4,4,5,5,6,6,6,6,7,7,1,2,3,3,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,4,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,3,4,4,5,5,6,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,6,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,7,7,7,7,7,7,7,7,7,7,0,0,1,1,1,1,2,2,3,3,3,4,5,5,6,7,0,1,1,2,2,3,3,3,4,4,5,5,6,6,6,7,0,1,2,3,3,4,4,5,5,5,6,6,6,7,7,7,1,2,3,3,4,4,5,5,6,6,6,6,7,7,7,7,1,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,0,0,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,3,4,4,5,5,6,6,6,6,7,7,7,7,1,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,7,7,1,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,1,2,2,3,4,4,4,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,6,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,2,3,3,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,7,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,4,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7);
  -- LUT for VNodeDegree 5
  constant LUT : LUTType := (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,3,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,4,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,3,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,1,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,0,1,1,1,1,2,2,4,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,3,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,1,2,2,2,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,3,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,1,2,2,2,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,1,2,2,2,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,0,0,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,1,2,2,2,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,6,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,0,1,1,1,1,2,2,4,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,1,1,1,1,2,2,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,4,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,4,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,0,0,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,4,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,3,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,1,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,3,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,1,2,2,2,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,1,2,2,2,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,6,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,0,0,0,0,1,1,1,1,1,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,6,7,0,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,5,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,0,1,1,1,1,2,2,4,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,2,2,2,3,3,4,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,3,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,3,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,1,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,3,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,2,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,7,0,1,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,6,6,6,6,6,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,3,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,3,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,1,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,7,7,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,3,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,7,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,3,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,0,1,1,1,1,2,2,4,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,1,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,1,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,7,7,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,0,0,0,0,0,0,0,0,0,1,1,1,1,2,2,4,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,1,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,3,4,4,5,6,7,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,5,5,5,6,6,6,6,6,7,7,7,7,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,1,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,5,5,5,6,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,3,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,5,5,5,6,6,6,6,6,7,7,7,7,0,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,6,7,0,1,2,3,3,4,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,5,5,5,6,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,4,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,2,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,7,0,1,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,6,6,6,6,6,7,7,7,7,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,1,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,5,5,5,6,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,5,5,5,6,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,4,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,6,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,4,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,3,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,1,2,2,2,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,3,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,1,2,2,2,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,3,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,3,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,1,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,7,7,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,3,4,4,5,6,7,0,1,1,2,2,3,3,3,4,4,5,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,2,2,2,3,4,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,4,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,7,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,3,4,4,5,6,7,0,1,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,1,2,2,2,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,3,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,2,2,2,3,4,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,3,5,0,0,0,0,0,1,1,1,1,2,2,2,3,4,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,7,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,0,0,0,0,1,1,1,1,1,2,2,2,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,3,5,6,6,6,6,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,1,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,7,7,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,4,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,7,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,0,0,1,1,1,1,2,2,3,3,5,0,0,0,0,1,1,1,1,1,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,7,7,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,3,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,1,2,2,2,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,3,4,4,5,6,7,0,1,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,7,0,0,0,0,1,1,1,1,1,2,2,2,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,6,7,7,7,7,7,7,7,7,7,7,4,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,3,5,6,6,6,6,7,7,7,7,7,7,7,7,7,7,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,7,7,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,3,5,6,6,6,6,7,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,1,2,2,2,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,0,0,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,1,2,2,2,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,6,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,3,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,7,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,3,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,1,2,2,2,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,3,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,2,2,2,3,4,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,3,5,0,0,0,0,0,1,1,1,1,2,2,2,3,4,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,7,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,0,0,0,0,1,1,1,1,1,2,2,2,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,3,5,6,6,6,6,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,3,5,0,0,0,0,0,1,1,1,1,2,2,2,3,4,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,7,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,3,4,4,5,5,5,6,6,7,0,1,2,3,3,4,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,6,6,6,6,6,7,7,7,7,2,4,4,5,5,6,6,6,6,7,7,7,7,7,7,7,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,0,1,2,3,3,4,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,6,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,3,5,5,6,6,6,6,7,7,7,7,7,7,7,7,7,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,5,5,6,6,6,6,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,0,0,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,6,6,6,6,6,7,7,7,7,2,4,4,5,5,6,6,6,6,7,7,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,0,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,3,5,6,6,6,6,7,7,7,7,7,7,7,7,7,7,0,0,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,6,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,6,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,1,2,2,2,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,6,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,0,0,0,0,1,1,1,1,1,2,2,2,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,0,1,2,3,3,4,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,6,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,3,5,5,6,6,6,6,7,7,7,7,7,7,7,7,7,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,0,0,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,6,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,6,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,3,5,5,6,6,6,6,7,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,3,5,6,6,6,6,7,7,7,7,7,7,7,7,7,7,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,5,5,6,6,6,6,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,6,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,3,5,5,6,6,6,6,7,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,6,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,0,1,1,1,1,2,2,4,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,1,1,1,1,2,2,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,4,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,0,1,1,1,1,2,2,4,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,1,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,1,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,7,7,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,0,0,0,0,0,0,0,0,0,1,1,1,1,2,2,4,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,1,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,3,4,4,5,6,7,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,5,5,5,6,6,6,6,6,7,7,7,7,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,1,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,5,5,5,6,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,1,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,7,7,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,4,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,7,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,0,0,1,1,1,1,2,2,3,3,5,0,0,0,0,1,1,1,1,1,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,7,7,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,3,0,0,0,0,0,0,0,0,0,1,1,1,1,2,2,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,0,0,0,0,0,0,0,0,0,1,1,1,1,2,2,4,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,1,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,3,4,4,5,6,7,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,0,0,0,0,0,0,0,1,1,1,1,2,2,3,3,5,0,0,0,0,1,1,1,1,1,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,3,4,4,5,6,7,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,0,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,3,4,5,5,5,6,6,6,6,7,7,7,7,7,2,4,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,4,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,5,5,5,6,6,6,6,6,7,7,7,7,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,0,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,3,4,5,5,5,6,6,6,6,7,7,7,7,7,2,4,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,3,4,5,5,5,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,3,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,4,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,5,5,5,6,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,3,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,4,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,0,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,4,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,1,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,5,5,5,6,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,7,7,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,5,5,5,6,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,4,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,0,0,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,4,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,2,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,3,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,3,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,5,5,5,6,6,6,6,6,7,7,7,7,0,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,6,7,0,1,2,3,3,4,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,5,5,5,6,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,4,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,0,0,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,6,6,6,6,6,7,7,7,7,2,4,4,5,5,6,6,6,6,7,7,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,0,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,3,5,6,6,6,6,7,7,7,7,7,7,7,7,7,7,0,0,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,6,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,6,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,1,1,1,1,2,4,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,0,0,0,0,0,0,0,1,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,5,5,5,6,6,6,6,6,7,7,7,7,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,0,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,3,4,5,5,5,6,6,6,6,7,7,7,7,7,2,4,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,3,4,5,5,5,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,3,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,4,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,5,5,5,6,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,1,1,1,1,2,3,4,0,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,0,1,1,1,1,2,2,2,3,4,5,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,6,7,0,1,2,3,3,4,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,0,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,3,5,6,6,6,6,7,7,7,7,7,7,7,7,7,7,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,3,4,5,5,5,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,0,1,2,3,3,4,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,6,7,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,0,0,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,6,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,3,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,4,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,4,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,5,5,5,6,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,4,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,6,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,5,5,5,6,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,6,7,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,4,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,3,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,1,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,3,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,1,2,2,2,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,1,2,2,2,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,6,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,0,0,0,0,1,1,1,1,1,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,6,7,0,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,5,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,3,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,1,2,2,2,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,3,4,4,5,6,7,0,1,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,7,0,0,0,0,1,1,1,1,1,2,2,2,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,6,7,7,7,7,7,7,7,7,7,7,4,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,1,1,1,2,2,4,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,1,2,2,2,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,6,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,0,0,0,0,1,1,1,1,1,2,2,2,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,0,1,2,3,3,4,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,6,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,3,5,5,6,6,6,6,7,7,7,7,7,7,7,7,7,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,0,0,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,6,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,6,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,3,5,5,6,6,6,6,7,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,3,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,4,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,0,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,4,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,1,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,0,0,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,6,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,3,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,4,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,4,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,1,1,1,1,1,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,6,7,0,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,5,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,0,1,1,1,2,2,3,3,3,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,6,7,7,7,7,7,7,7,7,7,7,4,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,6,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,4,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,4,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,3,4,4,5,5,5,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,6,7,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,3,5,5,6,6,6,6,7,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,2,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,0,0,0,1,1,1,2,4,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,0,0,0,0,0,0,0,0,1,1,1,1,2,2,3,5,0,0,0,0,0,1,1,1,1,2,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,7,0,1,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,6,6,6,6,6,7,7,7,7,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,1,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,5,5,5,6,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,5,5,5,6,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,4,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,6,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,4,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,0,1,1,1,1,1,2,3,5,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,0,0,0,0,0,1,1,1,1,1,2,2,2,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,3,5,6,6,6,6,7,7,7,7,7,7,7,7,7,7,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,7,7,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,3,5,6,6,6,6,7,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,0,0,1,1,1,1,2,2,3,4,5,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,3,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,4,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,3,5,6,6,6,6,7,7,7,7,7,7,7,7,7,7,0,0,1,1,2,2,2,3,3,3,4,4,5,5,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,2,2,3,4,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,5,5,6,6,6,6,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,6,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,3,5,5,6,6,6,6,7,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,6,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,0,1,1,1,1,1,2,2,3,3,4,6,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,0,0,0,1,1,1,1,2,2,2,3,3,4,5,5,6,0,1,1,1,2,2,2,3,3,4,4,5,5,6,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,5,5,5,6,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,0,0,1,1,1,2,2,3,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,5,5,5,6,6,7,7,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,0,1,2,2,3,3,4,4,4,5,5,5,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,5,5,5,6,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,0,0,1,1,1,1,2,2,2,3,3,4,5,6,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,0,0,1,1,1,2,2,2,3,3,4,4,5,5,6,7,0,1,1,2,2,3,3,4,4,4,5,5,6,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,5,5,5,6,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,4,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,0,1,2,2,3,3,4,4,4,5,5,6,6,6,7,7,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,6,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,5,5,5,6,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,6,7,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,4,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,0,1,1,1,1,2,2,2,3,3,4,4,5,6,6,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,0,1,2,2,3,3,4,4,5,5,5,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,5,6,6,6,6,7,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,2,2,3,4,4,5,5,5,6,6,6,6,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,6,7,7,7,7,7,7,7,3,5,5,6,6,6,6,7,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,3,4,5,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,4,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,0,1,1,2,2,2,3,3,4,4,5,5,5,6,6,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,1,1,2,3,3,4,4,5,5,5,6,6,6,6,7,7,1,2,3,4,4,5,5,6,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,4,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,2,3,4,4,5,5,5,6,6,6,6,7,7,7,7,2,3,4,5,5,6,6,6,6,6,7,7,7,7,7,7,3,4,5,6,6,6,6,7,7,7,7,7,7,7,7,7,3,5,6,6,6,6,7,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,1,3,4,4,5,5,6,6,6,6,6,7,7,7,7,7,2,4,5,5,6,6,6,6,7,7,7,7,7,7,7,7,3,5,6,6,6,6,7,7,7,7,7,7,7,7,7,7,4,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,2,3,4,5,5,6,6,6,6,7,7,7,7,7,7,7,3,5,5,6,6,6,7,7,7,7,7,7,7,7,7,7,4,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,2,4,5,6,6,6,6,6,7,7,7,7,7,7,7,7,4,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,3,5,6,6,6,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,5,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7);
  
  -- LUT address types
  subtype LUTAddr is integer range 0 to LUTSize-1;
  type LUTAddrType is array (0 to VNodeDegree-1) of LUTAddr;
  subtype LUTAddrSLV is std_logic_vector(0 to integer(ceil(log2(real(LUTSize))))-1);
  type LUTAddrSLVType is array (0 to VNodeDegree-1) of LUTAddrSLV;
  
end config;

package body config is

end config;
