library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
use work.config.all;

entity TopLevelDecoder is
  port (
    ChLLRxDI       : in ChLLRTypeStage;
    ClkxCI         : in std_logic;
    RstxRBI        : in std_logic;
    DecodedBitsxDO : out std_logic_vector(N-1 downto 0)
  );
end TopLevelDecoder;

architecture arch of TopLevelDecoder is

  component CNStage is
    port (
      ClkxCI           : in std_logic;
      RstxRBI          : in std_logic;
      IntLLRCNStagexDI : in IntLLRTypeCNStage;
      ChLLRCNStagexDI  : in ChLLRTypeStage;
      IntLLRCNStagexDO : out IntLLRTypeCNStage;
      ChLLRCNStagexDO  : out ChLLRTypeStage
  );
  end component;

  component VNStage_S0 is
    port (
      ClkxCI           : in std_logic;
      RstxRBI          : in std_logic;
      IntLLRVNStagexDI : in IntLLRTypeVNStage;
      ChLLRVNStagexDI  : in ChLLRTypeStage;
      IntLLRVNStagexDO : out IntLLRTypeVNStage;
      ChLLRVNStagexDO  : out ChLLRTypeStage
  );
  end component;

  component VNStage_S1 is
    port (
      ClkxCI           : in std_logic;
      RstxRBI          : in std_logic;
      IntLLRVNStagexDI : in IntLLRTypeVNStage;
      ChLLRVNStagexDI  : in ChLLRTypeStage;
      IntLLRVNStagexDO : out IntLLRTypeVNStage;
      ChLLRVNStagexDO  : out ChLLRTypeStage
  );
  end component;

  component VNStage_S2 is
    port (
      ClkxCI           : in std_logic;
      RstxRBI          : in std_logic;
      IntLLRVNStagexDI : in IntLLRTypeVNStage;
      ChLLRVNStagexDI  : in ChLLRTypeStage;
      IntLLRVNStagexDO : out IntLLRTypeVNStage;
      ChLLRVNStagexDO  : out ChLLRTypeStage
  );
  end component;

  component VNStage_S3 is
    port (
      ClkxCI           : in std_logic;
      RstxRBI          : in std_logic;
      IntLLRVNStagexDI : in IntLLRTypeVNStage;
      ChLLRVNStagexDI  : in ChLLRTypeStage;
      IntLLRVNStagexDO : out IntLLRTypeVNStage;
      ChLLRVNStagexDO  : out ChLLRTypeStage
  );
  end component;

  component VNStage_S4 is
    port (
      ClkxCI           : in std_logic;
      RstxRBI          : in std_logic;
      IntLLRVNStagexDI : in IntLLRTypeVNStage;
      ChLLRVNStagexDI  : in ChLLRTypeStage;
      IntLLRVNStagexDO : out IntLLRTypeVNStage;
      ChLLRVNStagexDO  : out ChLLRTypeStage
  );
  end component;

  component VNStage_S5 is
    port (
      ClkxCI           : in std_logic;
      RstxRBI          : in std_logic;
      IntLLRVNStagexDI : in IntLLRTypeVNStage;
      ChLLRVNStagexDI  : in ChLLRTypeStage;
      IntLLRVNStagexDO : out IntLLRTypeVNStage;
      ChLLRVNStagexDO  : out ChLLRTypeStage
  );
  end component;

  component VNStage_S6 is
    port (
      ClkxCI           : in std_logic;
      RstxRBI          : in std_logic;
      IntLLRVNStagexDI : in IntLLRTypeVNStage;
      ChLLRVNStagexDI  : in ChLLRTypeStage;
      IntLLRVNStagexDO : out IntLLRTypeVNStage;
      ChLLRVNStagexDO  : out ChLLRTypeStage
  );
  end component;

  component VNStage_S7 is
    port (
      ClkxCI           : in std_logic;
      RstxRBI          : in std_logic;
      IntLLRVNStagexDI : in IntLLRTypeVNStage;
      ChLLRVNStagexDI  : in ChLLRTypeStage;
      IntLLRVNStagexDO : out std_logic_vector(N-1 downto 0)
  );
  end component;

  -- VN Stage input signals
  signal VNStageIntLLRInputS0xD, VNStageIntLLRInputS1xD, VNStageIntLLRInputS2xD, VNStageIntLLRInputS3xD, VNStageIntLLRInputS4xD, VNStageIntLLRInputS5xD, VNStageIntLLRInputS6xD, VNStageIntLLRInputS7xD : IntLLRTypeVNStage;
  signal VNStageChLLRInputS0xD, VNStageChLLRInputS1xD, VNStageChLLRInputS2xD, VNStageChLLRInputS3xD, VNStageChLLRInputS4xD, VNStageChLLRInputS5xD, VNStageChLLRInputS6xD, VNStageChLLRInputS7xD : ChLLRTypeStage;

  -- VN Stage output signals
  signal VNStageIntLLROutputS0xD, VNStageIntLLROutputS1xD, VNStageIntLLROutputS2xD, VNStageIntLLROutputS3xD, VNStageIntLLROutputS4xD, VNStageIntLLROutputS5xD, VNStageIntLLROutputS6xD : IntLLRTypeVNStage;
  signal VNStageIntLLROutputS7xD : std_logic_vector(N-1 downto 0);
  signal VNStageChLLROutputS0xD, VNStageChLLROutputS1xD, VNStageChLLROutputS2xD, VNStageChLLROutputS3xD, VNStageChLLROutputS4xD, VNStageChLLROutputS5xD, VNStageChLLROutputS6xD : ChLLRTypeStage;

  -- CN Stage input signals
  signal CNStageIntLLRInputS0xD, CNStageIntLLRInputS1xD, CNStageIntLLRInputS2xD, CNStageIntLLRInputS3xD, CNStageIntLLRInputS4xD, CNStageIntLLRInputS5xD, CNStageIntLLRInputS6xD, CNStageIntLLRInputS7xD : IntLLRTypeCNStage;
  signal CNStageChLLRInputS0xD, CNStageChLLRInputS1xD, CNStageChLLRInputS2xD, CNStageChLLRInputS3xD, CNStageChLLRInputS4xD, CNStageChLLRInputS5xD, CNStageChLLRInputS6xD, CNStageChLLRInputS7xD : ChLLRTypeStage;

  -- CN Stage output signals
  signal CNStageIntLLROutputS0xD, CNStageIntLLROutputS1xD, CNStageIntLLROutputS2xD, CNStageIntLLROutputS3xD, CNStageIntLLROutputS4xD, CNStageIntLLROutputS5xD, CNStageIntLLROutputS6xD, CNStageIntLLROutputS7xD : IntLLRTypeCNStage;
  signal CNStageChLLROutputS0xD, CNStageChLLROutputS1xD, CNStageChLLROutputS2xD, CNStageChLLROutputS3xD, CNStageChLLROutputS4xD, CNStageChLLROutputS5xD, CNStageChLLROutputS6xD, CNStageChLLROutputS7xD : ChLLRTypeStage;

begin

  -- Instantiate CN and VN stages
  CNStage_0: CNStage port map(
    ClkxCI => ClkxCI,
    RstxRBI => RstxRBI,
    IntLLRCNStagexDI => CNStageIntLLRInputS0xD,
    ChLLRCNStagexDI => CNStageChLLRInputS0xD,
    IntLLRCNStagexDO => CNStageIntLLROutputS0xD,
    ChLLRCNStagexDO => CNStageChLLROutputS0xD
  );

  VNStage_0: VNStage_S0 port map(
    ClkxCI => ClkxCI,
    RstxRBI => RstxRBI,
    IntLLRVNStagexDI => VNStageIntLLRInputS0xD,
    ChLLRVNStagexDI => VNStageChLLRInputS0xD,
    IntLLRVNStagexDO => VNStageIntLLROutputS0xD,
    ChLLRVNStagexDO => VNStageChLLROutputS0xD
  );

  CNStage_1: CNStage port map(
    ClkxCI => ClkxCI,
    RstxRBI => RstxRBI,
    IntLLRCNStagexDI => CNStageIntLLRInputS1xD,
    ChLLRCNStagexDI => CNStageChLLRInputS1xD,
    IntLLRCNStagexDO => CNStageIntLLROutputS1xD,
    ChLLRCNStagexDO => CNStageChLLROutputS1xD
  );

  VNStage_1: VNStage_S1 port map(
    ClkxCI => ClkxCI,
    RstxRBI => RstxRBI,
    IntLLRVNStagexDI => VNStageIntLLRInputS1xD,
    ChLLRVNStagexDI => VNStageChLLRInputS1xD,
    IntLLRVNStagexDO => VNStageIntLLROutputS1xD,
    ChLLRVNStagexDO => VNStageChLLROutputS1xD
  );

  CNStage_2: CNStage port map(
    ClkxCI => ClkxCI,
    RstxRBI => RstxRBI,
    IntLLRCNStagexDI => CNStageIntLLRInputS2xD,
    ChLLRCNStagexDI => CNStageChLLRInputS2xD,
    IntLLRCNStagexDO => CNStageIntLLROutputS2xD,
    ChLLRCNStagexDO => CNStageChLLROutputS2xD
  );

  VNStage_2: VNStage_S2 port map(
    ClkxCI => ClkxCI,
    RstxRBI => RstxRBI,
    IntLLRVNStagexDI => VNStageIntLLRInputS2xD,
    ChLLRVNStagexDI => VNStageChLLRInputS2xD,
    IntLLRVNStagexDO => VNStageIntLLROutputS2xD,
    ChLLRVNStagexDO => VNStageChLLROutputS2xD
  );

  CNStage_3: CNStage port map(
    ClkxCI => ClkxCI,
    RstxRBI => RstxRBI,
    IntLLRCNStagexDI => CNStageIntLLRInputS3xD,
    ChLLRCNStagexDI => CNStageChLLRInputS3xD,
    IntLLRCNStagexDO => CNStageIntLLROutputS3xD,
    ChLLRCNStagexDO => CNStageChLLROutputS3xD
  );

  VNStage_3: VNStage_S3 port map(
    ClkxCI => ClkxCI,
    RstxRBI => RstxRBI,
    IntLLRVNStagexDI => VNStageIntLLRInputS3xD,
    ChLLRVNStagexDI => VNStageChLLRInputS3xD,
    IntLLRVNStagexDO => VNStageIntLLROutputS3xD,
    ChLLRVNStagexDO => VNStageChLLROutputS3xD
  );

  CNStage_4: CNStage port map(
    ClkxCI => ClkxCI,
    RstxRBI => RstxRBI,
    IntLLRCNStagexDI => CNStageIntLLRInputS4xD,
    ChLLRCNStagexDI => CNStageChLLRInputS4xD,
    IntLLRCNStagexDO => CNStageIntLLROutputS4xD,
    ChLLRCNStagexDO => CNStageChLLROutputS4xD
  );

  VNStage_4: VNStage_S4 port map(
    ClkxCI => ClkxCI,
    RstxRBI => RstxRBI,
    IntLLRVNStagexDI => VNStageIntLLRInputS4xD,
    ChLLRVNStagexDI => VNStageChLLRInputS4xD,
    IntLLRVNStagexDO => VNStageIntLLROutputS4xD,
    ChLLRVNStagexDO => VNStageChLLROutputS4xD
  );

  CNStage_5: CNStage port map(
    ClkxCI => ClkxCI,
    RstxRBI => RstxRBI,
    IntLLRCNStagexDI => CNStageIntLLRInputS5xD,
    ChLLRCNStagexDI => CNStageChLLRInputS5xD,
    IntLLRCNStagexDO => CNStageIntLLROutputS5xD,
    ChLLRCNStagexDO => CNStageChLLROutputS5xD
  );

  VNStage_5: VNStage_S5 port map(
    ClkxCI => ClkxCI,
    RstxRBI => RstxRBI,
    IntLLRVNStagexDI => VNStageIntLLRInputS5xD,
    ChLLRVNStagexDI => VNStageChLLRInputS5xD,
    IntLLRVNStagexDO => VNStageIntLLROutputS5xD,
    ChLLRVNStagexDO => VNStageChLLROutputS5xD
  );

  CNStage_6: CNStage port map(
    ClkxCI => ClkxCI,
    RstxRBI => RstxRBI,
    IntLLRCNStagexDI => CNStageIntLLRInputS6xD,
    ChLLRCNStagexDI => CNStageChLLRInputS6xD,
    IntLLRCNStagexDO => CNStageIntLLROutputS6xD,
    ChLLRCNStagexDO => CNStageChLLROutputS6xD
  );

  VNStage_6: VNStage_S6 port map(
    ClkxCI => ClkxCI,
    RstxRBI => RstxRBI,
    IntLLRVNStagexDI => VNStageIntLLRInputS6xD,
    ChLLRVNStagexDI => VNStageChLLRInputS6xD,
    IntLLRVNStagexDO => VNStageIntLLROutputS6xD,
    ChLLRVNStagexDO => VNStageChLLROutputS6xD
  );

  CNStage_7: CNStage port map(
    ClkxCI => ClkxCI,
    RstxRBI => RstxRBI,
    IntLLRCNStagexDI => CNStageIntLLRInputS7xD,
    ChLLRCNStagexDI => CNStageChLLRInputS7xD,
    IntLLRCNStagexDO => CNStageIntLLROutputS7xD,
    ChLLRCNStagexDO => CNStageChLLROutputS7xD
  );

  VNStage_7: VNStage_S7 port map(
    ClkxCI => ClkxCI,
    RstxRBI => RstxRBI,
    IntLLRVNStagexDI => VNStageIntLLRInputS7xD,
    ChLLRVNStagexDI => VNStageChLLRInputS7xD,
    IntLLRVNStagexDO => VNStageIntLLROutputS7xD
  );

  -- Connect input channel LLRS to first CN stage
  CNStageIntLLRInputS0xD(53)(0) <= LUT_4bit_to_3bit(ChLLRxDI(0));
  CNStageIntLLRInputS0xD(110)(0) <= LUT_4bit_to_3bit(ChLLRxDI(0));
  CNStageIntLLRInputS0xD(170)(0) <= LUT_4bit_to_3bit(ChLLRxDI(0));
  CNStageIntLLRInputS0xD(224)(0) <= LUT_4bit_to_3bit(ChLLRxDI(0));
  CNStageIntLLRInputS0xD(279)(0) <= LUT_4bit_to_3bit(ChLLRxDI(0));
  CNStageIntLLRInputS0xD(332)(0) <= LUT_4bit_to_3bit(ChLLRxDI(0));
  CNStageIntLLRInputS0xD(51)(0) <= LUT_4bit_to_3bit(ChLLRxDI(1));
  CNStageIntLLRInputS0xD(139)(0) <= LUT_4bit_to_3bit(ChLLRxDI(1));
  CNStageIntLLRInputS0xD(223)(0) <= LUT_4bit_to_3bit(ChLLRxDI(1));
  CNStageIntLLRInputS0xD(241)(0) <= LUT_4bit_to_3bit(ChLLRxDI(1));
  CNStageIntLLRInputS0xD(307)(0) <= LUT_4bit_to_3bit(ChLLRxDI(1));
  CNStageIntLLRInputS0xD(356)(0) <= LUT_4bit_to_3bit(ChLLRxDI(1));
  CNStageIntLLRInputS0xD(50)(0) <= LUT_4bit_to_3bit(ChLLRxDI(2));
  CNStageIntLLRInputS0xD(92)(0) <= LUT_4bit_to_3bit(ChLLRxDI(2));
  CNStageIntLLRInputS0xD(138)(0) <= LUT_4bit_to_3bit(ChLLRxDI(2));
  CNStageIntLLRInputS0xD(222)(0) <= LUT_4bit_to_3bit(ChLLRxDI(2));
  CNStageIntLLRInputS0xD(240)(0) <= LUT_4bit_to_3bit(ChLLRxDI(2));
  CNStageIntLLRInputS0xD(306)(0) <= LUT_4bit_to_3bit(ChLLRxDI(2));
  CNStageIntLLRInputS0xD(355)(0) <= LUT_4bit_to_3bit(ChLLRxDI(2));
  CNStageIntLLRInputS0xD(91)(0) <= LUT_4bit_to_3bit(ChLLRxDI(3));
  CNStageIntLLRInputS0xD(137)(0) <= LUT_4bit_to_3bit(ChLLRxDI(3));
  CNStageIntLLRInputS0xD(221)(0) <= LUT_4bit_to_3bit(ChLLRxDI(3));
  CNStageIntLLRInputS0xD(239)(0) <= LUT_4bit_to_3bit(ChLLRxDI(3));
  CNStageIntLLRInputS0xD(305)(0) <= LUT_4bit_to_3bit(ChLLRxDI(3));
  CNStageIntLLRInputS0xD(49)(0) <= LUT_4bit_to_3bit(ChLLRxDI(4));
  CNStageIntLLRInputS0xD(90)(0) <= LUT_4bit_to_3bit(ChLLRxDI(4));
  CNStageIntLLRInputS0xD(220)(0) <= LUT_4bit_to_3bit(ChLLRxDI(4));
  CNStageIntLLRInputS0xD(238)(0) <= LUT_4bit_to_3bit(ChLLRxDI(4));
  CNStageIntLLRInputS0xD(304)(0) <= LUT_4bit_to_3bit(ChLLRxDI(4));
  CNStageIntLLRInputS0xD(354)(0) <= LUT_4bit_to_3bit(ChLLRxDI(4));
  CNStageIntLLRInputS0xD(48)(0) <= LUT_4bit_to_3bit(ChLLRxDI(5));
  CNStageIntLLRInputS0xD(89)(0) <= LUT_4bit_to_3bit(ChLLRxDI(5));
  CNStageIntLLRInputS0xD(136)(0) <= LUT_4bit_to_3bit(ChLLRxDI(5));
  CNStageIntLLRInputS0xD(219)(0) <= LUT_4bit_to_3bit(ChLLRxDI(5));
  CNStageIntLLRInputS0xD(237)(0) <= LUT_4bit_to_3bit(ChLLRxDI(5));
  CNStageIntLLRInputS0xD(303)(0) <= LUT_4bit_to_3bit(ChLLRxDI(5));
  CNStageIntLLRInputS0xD(353)(0) <= LUT_4bit_to_3bit(ChLLRxDI(5));
  CNStageIntLLRInputS0xD(47)(0) <= LUT_4bit_to_3bit(ChLLRxDI(6));
  CNStageIntLLRInputS0xD(88)(0) <= LUT_4bit_to_3bit(ChLLRxDI(6));
  CNStageIntLLRInputS0xD(135)(0) <= LUT_4bit_to_3bit(ChLLRxDI(6));
  CNStageIntLLRInputS0xD(218)(0) <= LUT_4bit_to_3bit(ChLLRxDI(6));
  CNStageIntLLRInputS0xD(236)(0) <= LUT_4bit_to_3bit(ChLLRxDI(6));
  CNStageIntLLRInputS0xD(302)(0) <= LUT_4bit_to_3bit(ChLLRxDI(6));
  CNStageIntLLRInputS0xD(352)(0) <= LUT_4bit_to_3bit(ChLLRxDI(6));
  CNStageIntLLRInputS0xD(46)(0) <= LUT_4bit_to_3bit(ChLLRxDI(7));
  CNStageIntLLRInputS0xD(87)(0) <= LUT_4bit_to_3bit(ChLLRxDI(7));
  CNStageIntLLRInputS0xD(134)(0) <= LUT_4bit_to_3bit(ChLLRxDI(7));
  CNStageIntLLRInputS0xD(217)(0) <= LUT_4bit_to_3bit(ChLLRxDI(7));
  CNStageIntLLRInputS0xD(235)(0) <= LUT_4bit_to_3bit(ChLLRxDI(7));
  CNStageIntLLRInputS0xD(301)(0) <= LUT_4bit_to_3bit(ChLLRxDI(7));
  CNStageIntLLRInputS0xD(351)(0) <= LUT_4bit_to_3bit(ChLLRxDI(7));
  CNStageIntLLRInputS0xD(45)(0) <= LUT_4bit_to_3bit(ChLLRxDI(8));
  CNStageIntLLRInputS0xD(133)(0) <= LUT_4bit_to_3bit(ChLLRxDI(8));
  CNStageIntLLRInputS0xD(216)(0) <= LUT_4bit_to_3bit(ChLLRxDI(8));
  CNStageIntLLRInputS0xD(44)(0) <= LUT_4bit_to_3bit(ChLLRxDI(9));
  CNStageIntLLRInputS0xD(86)(0) <= LUT_4bit_to_3bit(ChLLRxDI(9));
  CNStageIntLLRInputS0xD(132)(0) <= LUT_4bit_to_3bit(ChLLRxDI(9));
  CNStageIntLLRInputS0xD(215)(0) <= LUT_4bit_to_3bit(ChLLRxDI(9));
  CNStageIntLLRInputS0xD(234)(0) <= LUT_4bit_to_3bit(ChLLRxDI(9));
  CNStageIntLLRInputS0xD(300)(0) <= LUT_4bit_to_3bit(ChLLRxDI(9));
  CNStageIntLLRInputS0xD(350)(0) <= LUT_4bit_to_3bit(ChLLRxDI(9));
  CNStageIntLLRInputS0xD(43)(0) <= LUT_4bit_to_3bit(ChLLRxDI(10));
  CNStageIntLLRInputS0xD(85)(0) <= LUT_4bit_to_3bit(ChLLRxDI(10));
  CNStageIntLLRInputS0xD(131)(0) <= LUT_4bit_to_3bit(ChLLRxDI(10));
  CNStageIntLLRInputS0xD(233)(0) <= LUT_4bit_to_3bit(ChLLRxDI(10));
  CNStageIntLLRInputS0xD(349)(0) <= LUT_4bit_to_3bit(ChLLRxDI(10));
  CNStageIntLLRInputS0xD(42)(0) <= LUT_4bit_to_3bit(ChLLRxDI(11));
  CNStageIntLLRInputS0xD(84)(0) <= LUT_4bit_to_3bit(ChLLRxDI(11));
  CNStageIntLLRInputS0xD(130)(0) <= LUT_4bit_to_3bit(ChLLRxDI(11));
  CNStageIntLLRInputS0xD(214)(0) <= LUT_4bit_to_3bit(ChLLRxDI(11));
  CNStageIntLLRInputS0xD(232)(0) <= LUT_4bit_to_3bit(ChLLRxDI(11));
  CNStageIntLLRInputS0xD(348)(0) <= LUT_4bit_to_3bit(ChLLRxDI(11));
  CNStageIntLLRInputS0xD(41)(0) <= LUT_4bit_to_3bit(ChLLRxDI(12));
  CNStageIntLLRInputS0xD(83)(0) <= LUT_4bit_to_3bit(ChLLRxDI(12));
  CNStageIntLLRInputS0xD(129)(0) <= LUT_4bit_to_3bit(ChLLRxDI(12));
  CNStageIntLLRInputS0xD(213)(0) <= LUT_4bit_to_3bit(ChLLRxDI(12));
  CNStageIntLLRInputS0xD(231)(0) <= LUT_4bit_to_3bit(ChLLRxDI(12));
  CNStageIntLLRInputS0xD(299)(0) <= LUT_4bit_to_3bit(ChLLRxDI(12));
  CNStageIntLLRInputS0xD(347)(0) <= LUT_4bit_to_3bit(ChLLRxDI(12));
  CNStageIntLLRInputS0xD(82)(0) <= LUT_4bit_to_3bit(ChLLRxDI(13));
  CNStageIntLLRInputS0xD(128)(0) <= LUT_4bit_to_3bit(ChLLRxDI(13));
  CNStageIntLLRInputS0xD(212)(0) <= LUT_4bit_to_3bit(ChLLRxDI(13));
  CNStageIntLLRInputS0xD(230)(0) <= LUT_4bit_to_3bit(ChLLRxDI(13));
  CNStageIntLLRInputS0xD(298)(0) <= LUT_4bit_to_3bit(ChLLRxDI(13));
  CNStageIntLLRInputS0xD(346)(0) <= LUT_4bit_to_3bit(ChLLRxDI(13));
  CNStageIntLLRInputS0xD(40)(0) <= LUT_4bit_to_3bit(ChLLRxDI(14));
  CNStageIntLLRInputS0xD(81)(0) <= LUT_4bit_to_3bit(ChLLRxDI(14));
  CNStageIntLLRInputS0xD(127)(0) <= LUT_4bit_to_3bit(ChLLRxDI(14));
  CNStageIntLLRInputS0xD(211)(0) <= LUT_4bit_to_3bit(ChLLRxDI(14));
  CNStageIntLLRInputS0xD(229)(0) <= LUT_4bit_to_3bit(ChLLRxDI(14));
  CNStageIntLLRInputS0xD(297)(0) <= LUT_4bit_to_3bit(ChLLRxDI(14));
  CNStageIntLLRInputS0xD(345)(0) <= LUT_4bit_to_3bit(ChLLRxDI(14));
  CNStageIntLLRInputS0xD(39)(0) <= LUT_4bit_to_3bit(ChLLRxDI(15));
  CNStageIntLLRInputS0xD(80)(0) <= LUT_4bit_to_3bit(ChLLRxDI(15));
  CNStageIntLLRInputS0xD(126)(0) <= LUT_4bit_to_3bit(ChLLRxDI(15));
  CNStageIntLLRInputS0xD(210)(0) <= LUT_4bit_to_3bit(ChLLRxDI(15));
  CNStageIntLLRInputS0xD(228)(0) <= LUT_4bit_to_3bit(ChLLRxDI(15));
  CNStageIntLLRInputS0xD(296)(0) <= LUT_4bit_to_3bit(ChLLRxDI(15));
  CNStageIntLLRInputS0xD(344)(0) <= LUT_4bit_to_3bit(ChLLRxDI(15));
  CNStageIntLLRInputS0xD(38)(0) <= LUT_4bit_to_3bit(ChLLRxDI(16));
  CNStageIntLLRInputS0xD(125)(0) <= LUT_4bit_to_3bit(ChLLRxDI(16));
  CNStageIntLLRInputS0xD(209)(0) <= LUT_4bit_to_3bit(ChLLRxDI(16));
  CNStageIntLLRInputS0xD(227)(0) <= LUT_4bit_to_3bit(ChLLRxDI(16));
  CNStageIntLLRInputS0xD(295)(0) <= LUT_4bit_to_3bit(ChLLRxDI(16));
  CNStageIntLLRInputS0xD(343)(0) <= LUT_4bit_to_3bit(ChLLRxDI(16));
  CNStageIntLLRInputS0xD(37)(0) <= LUT_4bit_to_3bit(ChLLRxDI(17));
  CNStageIntLLRInputS0xD(79)(0) <= LUT_4bit_to_3bit(ChLLRxDI(17));
  CNStageIntLLRInputS0xD(124)(0) <= LUT_4bit_to_3bit(ChLLRxDI(17));
  CNStageIntLLRInputS0xD(208)(0) <= LUT_4bit_to_3bit(ChLLRxDI(17));
  CNStageIntLLRInputS0xD(226)(0) <= LUT_4bit_to_3bit(ChLLRxDI(17));
  CNStageIntLLRInputS0xD(294)(0) <= LUT_4bit_to_3bit(ChLLRxDI(17));
  CNStageIntLLRInputS0xD(342)(0) <= LUT_4bit_to_3bit(ChLLRxDI(17));
  CNStageIntLLRInputS0xD(36)(0) <= LUT_4bit_to_3bit(ChLLRxDI(18));
  CNStageIntLLRInputS0xD(78)(0) <= LUT_4bit_to_3bit(ChLLRxDI(18));
  CNStageIntLLRInputS0xD(123)(0) <= LUT_4bit_to_3bit(ChLLRxDI(18));
  CNStageIntLLRInputS0xD(207)(0) <= LUT_4bit_to_3bit(ChLLRxDI(18));
  CNStageIntLLRInputS0xD(225)(0) <= LUT_4bit_to_3bit(ChLLRxDI(18));
  CNStageIntLLRInputS0xD(293)(0) <= LUT_4bit_to_3bit(ChLLRxDI(18));
  CNStageIntLLRInputS0xD(341)(0) <= LUT_4bit_to_3bit(ChLLRxDI(18));
  CNStageIntLLRInputS0xD(35)(0) <= LUT_4bit_to_3bit(ChLLRxDI(19));
  CNStageIntLLRInputS0xD(77)(0) <= LUT_4bit_to_3bit(ChLLRxDI(19));
  CNStageIntLLRInputS0xD(122)(0) <= LUT_4bit_to_3bit(ChLLRxDI(19));
  CNStageIntLLRInputS0xD(278)(0) <= LUT_4bit_to_3bit(ChLLRxDI(19));
  CNStageIntLLRInputS0xD(340)(0) <= LUT_4bit_to_3bit(ChLLRxDI(19));
  CNStageIntLLRInputS0xD(34)(0) <= LUT_4bit_to_3bit(ChLLRxDI(20));
  CNStageIntLLRInputS0xD(76)(0) <= LUT_4bit_to_3bit(ChLLRxDI(20));
  CNStageIntLLRInputS0xD(277)(0) <= LUT_4bit_to_3bit(ChLLRxDI(20));
  CNStageIntLLRInputS0xD(292)(0) <= LUT_4bit_to_3bit(ChLLRxDI(20));
  CNStageIntLLRInputS0xD(339)(0) <= LUT_4bit_to_3bit(ChLLRxDI(20));
  CNStageIntLLRInputS0xD(33)(0) <= LUT_4bit_to_3bit(ChLLRxDI(21));
  CNStageIntLLRInputS0xD(75)(0) <= LUT_4bit_to_3bit(ChLLRxDI(21));
  CNStageIntLLRInputS0xD(121)(0) <= LUT_4bit_to_3bit(ChLLRxDI(21));
  CNStageIntLLRInputS0xD(206)(0) <= LUT_4bit_to_3bit(ChLLRxDI(21));
  CNStageIntLLRInputS0xD(276)(0) <= LUT_4bit_to_3bit(ChLLRxDI(21));
  CNStageIntLLRInputS0xD(291)(0) <= LUT_4bit_to_3bit(ChLLRxDI(21));
  CNStageIntLLRInputS0xD(338)(0) <= LUT_4bit_to_3bit(ChLLRxDI(21));
  CNStageIntLLRInputS0xD(32)(0) <= LUT_4bit_to_3bit(ChLLRxDI(22));
  CNStageIntLLRInputS0xD(74)(0) <= LUT_4bit_to_3bit(ChLLRxDI(22));
  CNStageIntLLRInputS0xD(120)(0) <= LUT_4bit_to_3bit(ChLLRxDI(22));
  CNStageIntLLRInputS0xD(205)(0) <= LUT_4bit_to_3bit(ChLLRxDI(22));
  CNStageIntLLRInputS0xD(275)(0) <= LUT_4bit_to_3bit(ChLLRxDI(22));
  CNStageIntLLRInputS0xD(290)(0) <= LUT_4bit_to_3bit(ChLLRxDI(22));
  CNStageIntLLRInputS0xD(337)(0) <= LUT_4bit_to_3bit(ChLLRxDI(22));
  CNStageIntLLRInputS0xD(31)(0) <= LUT_4bit_to_3bit(ChLLRxDI(23));
  CNStageIntLLRInputS0xD(73)(0) <= LUT_4bit_to_3bit(ChLLRxDI(23));
  CNStageIntLLRInputS0xD(119)(0) <= LUT_4bit_to_3bit(ChLLRxDI(23));
  CNStageIntLLRInputS0xD(204)(0) <= LUT_4bit_to_3bit(ChLLRxDI(23));
  CNStageIntLLRInputS0xD(274)(0) <= LUT_4bit_to_3bit(ChLLRxDI(23));
  CNStageIntLLRInputS0xD(289)(0) <= LUT_4bit_to_3bit(ChLLRxDI(23));
  CNStageIntLLRInputS0xD(336)(0) <= LUT_4bit_to_3bit(ChLLRxDI(23));
  CNStageIntLLRInputS0xD(30)(0) <= LUT_4bit_to_3bit(ChLLRxDI(24));
  CNStageIntLLRInputS0xD(72)(0) <= LUT_4bit_to_3bit(ChLLRxDI(24));
  CNStageIntLLRInputS0xD(118)(0) <= LUT_4bit_to_3bit(ChLLRxDI(24));
  CNStageIntLLRInputS0xD(203)(0) <= LUT_4bit_to_3bit(ChLLRxDI(24));
  CNStageIntLLRInputS0xD(273)(0) <= LUT_4bit_to_3bit(ChLLRxDI(24));
  CNStageIntLLRInputS0xD(288)(0) <= LUT_4bit_to_3bit(ChLLRxDI(24));
  CNStageIntLLRInputS0xD(335)(0) <= LUT_4bit_to_3bit(ChLLRxDI(24));
  CNStageIntLLRInputS0xD(29)(0) <= LUT_4bit_to_3bit(ChLLRxDI(25));
  CNStageIntLLRInputS0xD(71)(0) <= LUT_4bit_to_3bit(ChLLRxDI(25));
  CNStageIntLLRInputS0xD(117)(0) <= LUT_4bit_to_3bit(ChLLRxDI(25));
  CNStageIntLLRInputS0xD(202)(0) <= LUT_4bit_to_3bit(ChLLRxDI(25));
  CNStageIntLLRInputS0xD(287)(0) <= LUT_4bit_to_3bit(ChLLRxDI(25));
  CNStageIntLLRInputS0xD(28)(0) <= LUT_4bit_to_3bit(ChLLRxDI(26));
  CNStageIntLLRInputS0xD(70)(0) <= LUT_4bit_to_3bit(ChLLRxDI(26));
  CNStageIntLLRInputS0xD(116)(0) <= LUT_4bit_to_3bit(ChLLRxDI(26));
  CNStageIntLLRInputS0xD(201)(0) <= LUT_4bit_to_3bit(ChLLRxDI(26));
  CNStageIntLLRInputS0xD(272)(0) <= LUT_4bit_to_3bit(ChLLRxDI(26));
  CNStageIntLLRInputS0xD(286)(0) <= LUT_4bit_to_3bit(ChLLRxDI(26));
  CNStageIntLLRInputS0xD(334)(0) <= LUT_4bit_to_3bit(ChLLRxDI(26));
  CNStageIntLLRInputS0xD(27)(0) <= LUT_4bit_to_3bit(ChLLRxDI(27));
  CNStageIntLLRInputS0xD(69)(0) <= LUT_4bit_to_3bit(ChLLRxDI(27));
  CNStageIntLLRInputS0xD(115)(0) <= LUT_4bit_to_3bit(ChLLRxDI(27));
  CNStageIntLLRInputS0xD(200)(0) <= LUT_4bit_to_3bit(ChLLRxDI(27));
  CNStageIntLLRInputS0xD(285)(0) <= LUT_4bit_to_3bit(ChLLRxDI(27));
  CNStageIntLLRInputS0xD(26)(0) <= LUT_4bit_to_3bit(ChLLRxDI(28));
  CNStageIntLLRInputS0xD(68)(0) <= LUT_4bit_to_3bit(ChLLRxDI(28));
  CNStageIntLLRInputS0xD(114)(0) <= LUT_4bit_to_3bit(ChLLRxDI(28));
  CNStageIntLLRInputS0xD(199)(0) <= LUT_4bit_to_3bit(ChLLRxDI(28));
  CNStageIntLLRInputS0xD(271)(0) <= LUT_4bit_to_3bit(ChLLRxDI(28));
  CNStageIntLLRInputS0xD(333)(0) <= LUT_4bit_to_3bit(ChLLRxDI(28));
  CNStageIntLLRInputS0xD(25)(0) <= LUT_4bit_to_3bit(ChLLRxDI(29));
  CNStageIntLLRInputS0xD(67)(0) <= LUT_4bit_to_3bit(ChLLRxDI(29));
  CNStageIntLLRInputS0xD(113)(0) <= LUT_4bit_to_3bit(ChLLRxDI(29));
  CNStageIntLLRInputS0xD(270)(0) <= LUT_4bit_to_3bit(ChLLRxDI(29));
  CNStageIntLLRInputS0xD(24)(0) <= LUT_4bit_to_3bit(ChLLRxDI(30));
  CNStageIntLLRInputS0xD(66)(0) <= LUT_4bit_to_3bit(ChLLRxDI(30));
  CNStageIntLLRInputS0xD(112)(0) <= LUT_4bit_to_3bit(ChLLRxDI(30));
  CNStageIntLLRInputS0xD(198)(0) <= LUT_4bit_to_3bit(ChLLRxDI(30));
  CNStageIntLLRInputS0xD(269)(0) <= LUT_4bit_to_3bit(ChLLRxDI(30));
  CNStageIntLLRInputS0xD(284)(0) <= LUT_4bit_to_3bit(ChLLRxDI(30));
  CNStageIntLLRInputS0xD(23)(0) <= LUT_4bit_to_3bit(ChLLRxDI(31));
  CNStageIntLLRInputS0xD(65)(0) <= LUT_4bit_to_3bit(ChLLRxDI(31));
  CNStageIntLLRInputS0xD(197)(0) <= LUT_4bit_to_3bit(ChLLRxDI(31));
  CNStageIntLLRInputS0xD(283)(0) <= LUT_4bit_to_3bit(ChLLRxDI(31));
  CNStageIntLLRInputS0xD(22)(0) <= LUT_4bit_to_3bit(ChLLRxDI(32));
  CNStageIntLLRInputS0xD(64)(0) <= LUT_4bit_to_3bit(ChLLRxDI(32));
  CNStageIntLLRInputS0xD(111)(0) <= LUT_4bit_to_3bit(ChLLRxDI(32));
  CNStageIntLLRInputS0xD(268)(0) <= LUT_4bit_to_3bit(ChLLRxDI(32));
  CNStageIntLLRInputS0xD(21)(0) <= LUT_4bit_to_3bit(ChLLRxDI(33));
  CNStageIntLLRInputS0xD(63)(0) <= LUT_4bit_to_3bit(ChLLRxDI(33));
  CNStageIntLLRInputS0xD(169)(0) <= LUT_4bit_to_3bit(ChLLRxDI(33));
  CNStageIntLLRInputS0xD(196)(0) <= LUT_4bit_to_3bit(ChLLRxDI(33));
  CNStageIntLLRInputS0xD(267)(0) <= LUT_4bit_to_3bit(ChLLRxDI(33));
  CNStageIntLLRInputS0xD(282)(0) <= LUT_4bit_to_3bit(ChLLRxDI(33));
  CNStageIntLLRInputS0xD(20)(0) <= LUT_4bit_to_3bit(ChLLRxDI(34));
  CNStageIntLLRInputS0xD(62)(0) <= LUT_4bit_to_3bit(ChLLRxDI(34));
  CNStageIntLLRInputS0xD(168)(0) <= LUT_4bit_to_3bit(ChLLRxDI(34));
  CNStageIntLLRInputS0xD(195)(0) <= LUT_4bit_to_3bit(ChLLRxDI(34));
  CNStageIntLLRInputS0xD(266)(0) <= LUT_4bit_to_3bit(ChLLRxDI(34));
  CNStageIntLLRInputS0xD(281)(0) <= LUT_4bit_to_3bit(ChLLRxDI(34));
  CNStageIntLLRInputS0xD(19)(0) <= LUT_4bit_to_3bit(ChLLRxDI(35));
  CNStageIntLLRInputS0xD(61)(0) <= LUT_4bit_to_3bit(ChLLRxDI(35));
  CNStageIntLLRInputS0xD(167)(0) <= LUT_4bit_to_3bit(ChLLRxDI(35));
  CNStageIntLLRInputS0xD(194)(0) <= LUT_4bit_to_3bit(ChLLRxDI(35));
  CNStageIntLLRInputS0xD(265)(0) <= LUT_4bit_to_3bit(ChLLRxDI(35));
  CNStageIntLLRInputS0xD(280)(0) <= LUT_4bit_to_3bit(ChLLRxDI(35));
  CNStageIntLLRInputS0xD(18)(0) <= LUT_4bit_to_3bit(ChLLRxDI(36));
  CNStageIntLLRInputS0xD(60)(0) <= LUT_4bit_to_3bit(ChLLRxDI(36));
  CNStageIntLLRInputS0xD(166)(0) <= LUT_4bit_to_3bit(ChLLRxDI(36));
  CNStageIntLLRInputS0xD(264)(0) <= LUT_4bit_to_3bit(ChLLRxDI(36));
  CNStageIntLLRInputS0xD(17)(0) <= LUT_4bit_to_3bit(ChLLRxDI(37));
  CNStageIntLLRInputS0xD(59)(0) <= LUT_4bit_to_3bit(ChLLRxDI(37));
  CNStageIntLLRInputS0xD(165)(0) <= LUT_4bit_to_3bit(ChLLRxDI(37));
  CNStageIntLLRInputS0xD(193)(0) <= LUT_4bit_to_3bit(ChLLRxDI(37));
  CNStageIntLLRInputS0xD(263)(0) <= LUT_4bit_to_3bit(ChLLRxDI(37));
  CNStageIntLLRInputS0xD(331)(0) <= LUT_4bit_to_3bit(ChLLRxDI(37));
  CNStageIntLLRInputS0xD(383)(0) <= LUT_4bit_to_3bit(ChLLRxDI(37));
  CNStageIntLLRInputS0xD(16)(0) <= LUT_4bit_to_3bit(ChLLRxDI(38));
  CNStageIntLLRInputS0xD(58)(0) <= LUT_4bit_to_3bit(ChLLRxDI(38));
  CNStageIntLLRInputS0xD(164)(0) <= LUT_4bit_to_3bit(ChLLRxDI(38));
  CNStageIntLLRInputS0xD(192)(0) <= LUT_4bit_to_3bit(ChLLRxDI(38));
  CNStageIntLLRInputS0xD(262)(0) <= LUT_4bit_to_3bit(ChLLRxDI(38));
  CNStageIntLLRInputS0xD(330)(0) <= LUT_4bit_to_3bit(ChLLRxDI(38));
  CNStageIntLLRInputS0xD(382)(0) <= LUT_4bit_to_3bit(ChLLRxDI(38));
  CNStageIntLLRInputS0xD(15)(0) <= LUT_4bit_to_3bit(ChLLRxDI(39));
  CNStageIntLLRInputS0xD(57)(0) <= LUT_4bit_to_3bit(ChLLRxDI(39));
  CNStageIntLLRInputS0xD(163)(0) <= LUT_4bit_to_3bit(ChLLRxDI(39));
  CNStageIntLLRInputS0xD(191)(0) <= LUT_4bit_to_3bit(ChLLRxDI(39));
  CNStageIntLLRInputS0xD(261)(0) <= LUT_4bit_to_3bit(ChLLRxDI(39));
  CNStageIntLLRInputS0xD(329)(0) <= LUT_4bit_to_3bit(ChLLRxDI(39));
  CNStageIntLLRInputS0xD(381)(0) <= LUT_4bit_to_3bit(ChLLRxDI(39));
  CNStageIntLLRInputS0xD(14)(0) <= LUT_4bit_to_3bit(ChLLRxDI(40));
  CNStageIntLLRInputS0xD(56)(0) <= LUT_4bit_to_3bit(ChLLRxDI(40));
  CNStageIntLLRInputS0xD(162)(0) <= LUT_4bit_to_3bit(ChLLRxDI(40));
  CNStageIntLLRInputS0xD(260)(0) <= LUT_4bit_to_3bit(ChLLRxDI(40));
  CNStageIntLLRInputS0xD(380)(0) <= LUT_4bit_to_3bit(ChLLRxDI(40));
  CNStageIntLLRInputS0xD(13)(0) <= LUT_4bit_to_3bit(ChLLRxDI(41));
  CNStageIntLLRInputS0xD(55)(0) <= LUT_4bit_to_3bit(ChLLRxDI(41));
  CNStageIntLLRInputS0xD(161)(0) <= LUT_4bit_to_3bit(ChLLRxDI(41));
  CNStageIntLLRInputS0xD(190)(0) <= LUT_4bit_to_3bit(ChLLRxDI(41));
  CNStageIntLLRInputS0xD(259)(0) <= LUT_4bit_to_3bit(ChLLRxDI(41));
  CNStageIntLLRInputS0xD(328)(0) <= LUT_4bit_to_3bit(ChLLRxDI(41));
  CNStageIntLLRInputS0xD(379)(0) <= LUT_4bit_to_3bit(ChLLRxDI(41));
  CNStageIntLLRInputS0xD(12)(0) <= LUT_4bit_to_3bit(ChLLRxDI(42));
  CNStageIntLLRInputS0xD(54)(0) <= LUT_4bit_to_3bit(ChLLRxDI(42));
  CNStageIntLLRInputS0xD(160)(0) <= LUT_4bit_to_3bit(ChLLRxDI(42));
  CNStageIntLLRInputS0xD(189)(0) <= LUT_4bit_to_3bit(ChLLRxDI(42));
  CNStageIntLLRInputS0xD(258)(0) <= LUT_4bit_to_3bit(ChLLRxDI(42));
  CNStageIntLLRInputS0xD(327)(0) <= LUT_4bit_to_3bit(ChLLRxDI(42));
  CNStageIntLLRInputS0xD(378)(0) <= LUT_4bit_to_3bit(ChLLRxDI(42));
  CNStageIntLLRInputS0xD(109)(0) <= LUT_4bit_to_3bit(ChLLRxDI(43));
  CNStageIntLLRInputS0xD(159)(0) <= LUT_4bit_to_3bit(ChLLRxDI(43));
  CNStageIntLLRInputS0xD(188)(0) <= LUT_4bit_to_3bit(ChLLRxDI(43));
  CNStageIntLLRInputS0xD(257)(0) <= LUT_4bit_to_3bit(ChLLRxDI(43));
  CNStageIntLLRInputS0xD(326)(0) <= LUT_4bit_to_3bit(ChLLRxDI(43));
  CNStageIntLLRInputS0xD(377)(0) <= LUT_4bit_to_3bit(ChLLRxDI(43));
  CNStageIntLLRInputS0xD(11)(0) <= LUT_4bit_to_3bit(ChLLRxDI(44));
  CNStageIntLLRInputS0xD(108)(0) <= LUT_4bit_to_3bit(ChLLRxDI(44));
  CNStageIntLLRInputS0xD(158)(0) <= LUT_4bit_to_3bit(ChLLRxDI(44));
  CNStageIntLLRInputS0xD(187)(0) <= LUT_4bit_to_3bit(ChLLRxDI(44));
  CNStageIntLLRInputS0xD(256)(0) <= LUT_4bit_to_3bit(ChLLRxDI(44));
  CNStageIntLLRInputS0xD(325)(0) <= LUT_4bit_to_3bit(ChLLRxDI(44));
  CNStageIntLLRInputS0xD(376)(0) <= LUT_4bit_to_3bit(ChLLRxDI(44));
  CNStageIntLLRInputS0xD(10)(0) <= LUT_4bit_to_3bit(ChLLRxDI(45));
  CNStageIntLLRInputS0xD(107)(0) <= LUT_4bit_to_3bit(ChLLRxDI(45));
  CNStageIntLLRInputS0xD(157)(0) <= LUT_4bit_to_3bit(ChLLRxDI(45));
  CNStageIntLLRInputS0xD(186)(0) <= LUT_4bit_to_3bit(ChLLRxDI(45));
  CNStageIntLLRInputS0xD(255)(0) <= LUT_4bit_to_3bit(ChLLRxDI(45));
  CNStageIntLLRInputS0xD(324)(0) <= LUT_4bit_to_3bit(ChLLRxDI(45));
  CNStageIntLLRInputS0xD(375)(0) <= LUT_4bit_to_3bit(ChLLRxDI(45));
  CNStageIntLLRInputS0xD(9)(0) <= LUT_4bit_to_3bit(ChLLRxDI(46));
  CNStageIntLLRInputS0xD(106)(0) <= LUT_4bit_to_3bit(ChLLRxDI(46));
  CNStageIntLLRInputS0xD(156)(0) <= LUT_4bit_to_3bit(ChLLRxDI(46));
  CNStageIntLLRInputS0xD(185)(0) <= LUT_4bit_to_3bit(ChLLRxDI(46));
  CNStageIntLLRInputS0xD(254)(0) <= LUT_4bit_to_3bit(ChLLRxDI(46));
  CNStageIntLLRInputS0xD(323)(0) <= LUT_4bit_to_3bit(ChLLRxDI(46));
  CNStageIntLLRInputS0xD(374)(0) <= LUT_4bit_to_3bit(ChLLRxDI(46));
  CNStageIntLLRInputS0xD(8)(0) <= LUT_4bit_to_3bit(ChLLRxDI(47));
  CNStageIntLLRInputS0xD(155)(0) <= LUT_4bit_to_3bit(ChLLRxDI(47));
  CNStageIntLLRInputS0xD(253)(0) <= LUT_4bit_to_3bit(ChLLRxDI(47));
  CNStageIntLLRInputS0xD(373)(0) <= LUT_4bit_to_3bit(ChLLRxDI(47));
  CNStageIntLLRInputS0xD(7)(0) <= LUT_4bit_to_3bit(ChLLRxDI(48));
  CNStageIntLLRInputS0xD(154)(0) <= LUT_4bit_to_3bit(ChLLRxDI(48));
  CNStageIntLLRInputS0xD(322)(0) <= LUT_4bit_to_3bit(ChLLRxDI(48));
  CNStageIntLLRInputS0xD(372)(0) <= LUT_4bit_to_3bit(ChLLRxDI(48));
  CNStageIntLLRInputS0xD(6)(0) <= LUT_4bit_to_3bit(ChLLRxDI(49));
  CNStageIntLLRInputS0xD(105)(0) <= LUT_4bit_to_3bit(ChLLRxDI(49));
  CNStageIntLLRInputS0xD(153)(0) <= LUT_4bit_to_3bit(ChLLRxDI(49));
  CNStageIntLLRInputS0xD(184)(0) <= LUT_4bit_to_3bit(ChLLRxDI(49));
  CNStageIntLLRInputS0xD(252)(0) <= LUT_4bit_to_3bit(ChLLRxDI(49));
  CNStageIntLLRInputS0xD(321)(0) <= LUT_4bit_to_3bit(ChLLRxDI(49));
  CNStageIntLLRInputS0xD(371)(0) <= LUT_4bit_to_3bit(ChLLRxDI(49));
  CNStageIntLLRInputS0xD(5)(0) <= LUT_4bit_to_3bit(ChLLRxDI(50));
  CNStageIntLLRInputS0xD(104)(0) <= LUT_4bit_to_3bit(ChLLRxDI(50));
  CNStageIntLLRInputS0xD(152)(0) <= LUT_4bit_to_3bit(ChLLRxDI(50));
  CNStageIntLLRInputS0xD(183)(0) <= LUT_4bit_to_3bit(ChLLRxDI(50));
  CNStageIntLLRInputS0xD(251)(0) <= LUT_4bit_to_3bit(ChLLRxDI(50));
  CNStageIntLLRInputS0xD(320)(0) <= LUT_4bit_to_3bit(ChLLRxDI(50));
  CNStageIntLLRInputS0xD(370)(0) <= LUT_4bit_to_3bit(ChLLRxDI(50));
  CNStageIntLLRInputS0xD(4)(0) <= LUT_4bit_to_3bit(ChLLRxDI(51));
  CNStageIntLLRInputS0xD(103)(0) <= LUT_4bit_to_3bit(ChLLRxDI(51));
  CNStageIntLLRInputS0xD(182)(0) <= LUT_4bit_to_3bit(ChLLRxDI(51));
  CNStageIntLLRInputS0xD(250)(0) <= LUT_4bit_to_3bit(ChLLRxDI(51));
  CNStageIntLLRInputS0xD(319)(0) <= LUT_4bit_to_3bit(ChLLRxDI(51));
  CNStageIntLLRInputS0xD(369)(0) <= LUT_4bit_to_3bit(ChLLRxDI(51));
  CNStageIntLLRInputS0xD(102)(0) <= LUT_4bit_to_3bit(ChLLRxDI(52));
  CNStageIntLLRInputS0xD(151)(0) <= LUT_4bit_to_3bit(ChLLRxDI(52));
  CNStageIntLLRInputS0xD(181)(0) <= LUT_4bit_to_3bit(ChLLRxDI(52));
  CNStageIntLLRInputS0xD(318)(0) <= LUT_4bit_to_3bit(ChLLRxDI(52));
  CNStageIntLLRInputS0xD(368)(0) <= LUT_4bit_to_3bit(ChLLRxDI(52));
  CNStageIntLLRInputS0xD(3)(0) <= LUT_4bit_to_3bit(ChLLRxDI(53));
  CNStageIntLLRInputS0xD(150)(0) <= LUT_4bit_to_3bit(ChLLRxDI(53));
  CNStageIntLLRInputS0xD(180)(0) <= LUT_4bit_to_3bit(ChLLRxDI(53));
  CNStageIntLLRInputS0xD(249)(0) <= LUT_4bit_to_3bit(ChLLRxDI(53));
  CNStageIntLLRInputS0xD(317)(0) <= LUT_4bit_to_3bit(ChLLRxDI(53));
  CNStageIntLLRInputS0xD(367)(0) <= LUT_4bit_to_3bit(ChLLRxDI(53));
  CNStageIntLLRInputS0xD(2)(0) <= LUT_4bit_to_3bit(ChLLRxDI(54));
  CNStageIntLLRInputS0xD(101)(0) <= LUT_4bit_to_3bit(ChLLRxDI(54));
  CNStageIntLLRInputS0xD(149)(0) <= LUT_4bit_to_3bit(ChLLRxDI(54));
  CNStageIntLLRInputS0xD(179)(0) <= LUT_4bit_to_3bit(ChLLRxDI(54));
  CNStageIntLLRInputS0xD(316)(0) <= LUT_4bit_to_3bit(ChLLRxDI(54));
  CNStageIntLLRInputS0xD(366)(0) <= LUT_4bit_to_3bit(ChLLRxDI(54));
  CNStageIntLLRInputS0xD(1)(0) <= LUT_4bit_to_3bit(ChLLRxDI(55));
  CNStageIntLLRInputS0xD(100)(0) <= LUT_4bit_to_3bit(ChLLRxDI(55));
  CNStageIntLLRInputS0xD(148)(0) <= LUT_4bit_to_3bit(ChLLRxDI(55));
  CNStageIntLLRInputS0xD(178)(0) <= LUT_4bit_to_3bit(ChLLRxDI(55));
  CNStageIntLLRInputS0xD(248)(0) <= LUT_4bit_to_3bit(ChLLRxDI(55));
  CNStageIntLLRInputS0xD(315)(0) <= LUT_4bit_to_3bit(ChLLRxDI(55));
  CNStageIntLLRInputS0xD(365)(0) <= LUT_4bit_to_3bit(ChLLRxDI(55));
  CNStageIntLLRInputS0xD(0)(0) <= LUT_4bit_to_3bit(ChLLRxDI(56));
  CNStageIntLLRInputS0xD(99)(0) <= LUT_4bit_to_3bit(ChLLRxDI(56));
  CNStageIntLLRInputS0xD(147)(0) <= LUT_4bit_to_3bit(ChLLRxDI(56));
  CNStageIntLLRInputS0xD(177)(0) <= LUT_4bit_to_3bit(ChLLRxDI(56));
  CNStageIntLLRInputS0xD(247)(0) <= LUT_4bit_to_3bit(ChLLRxDI(56));
  CNStageIntLLRInputS0xD(314)(0) <= LUT_4bit_to_3bit(ChLLRxDI(56));
  CNStageIntLLRInputS0xD(364)(0) <= LUT_4bit_to_3bit(ChLLRxDI(56));
  CNStageIntLLRInputS0xD(98)(0) <= LUT_4bit_to_3bit(ChLLRxDI(57));
  CNStageIntLLRInputS0xD(146)(0) <= LUT_4bit_to_3bit(ChLLRxDI(57));
  CNStageIntLLRInputS0xD(176)(0) <= LUT_4bit_to_3bit(ChLLRxDI(57));
  CNStageIntLLRInputS0xD(246)(0) <= LUT_4bit_to_3bit(ChLLRxDI(57));
  CNStageIntLLRInputS0xD(313)(0) <= LUT_4bit_to_3bit(ChLLRxDI(57));
  CNStageIntLLRInputS0xD(363)(0) <= LUT_4bit_to_3bit(ChLLRxDI(57));
  CNStageIntLLRInputS0xD(97)(0) <= LUT_4bit_to_3bit(ChLLRxDI(58));
  CNStageIntLLRInputS0xD(145)(0) <= LUT_4bit_to_3bit(ChLLRxDI(58));
  CNStageIntLLRInputS0xD(175)(0) <= LUT_4bit_to_3bit(ChLLRxDI(58));
  CNStageIntLLRInputS0xD(312)(0) <= LUT_4bit_to_3bit(ChLLRxDI(58));
  CNStageIntLLRInputS0xD(362)(0) <= LUT_4bit_to_3bit(ChLLRxDI(58));
  CNStageIntLLRInputS0xD(144)(0) <= LUT_4bit_to_3bit(ChLLRxDI(59));
  CNStageIntLLRInputS0xD(174)(0) <= LUT_4bit_to_3bit(ChLLRxDI(59));
  CNStageIntLLRInputS0xD(245)(0) <= LUT_4bit_to_3bit(ChLLRxDI(59));
  CNStageIntLLRInputS0xD(311)(0) <= LUT_4bit_to_3bit(ChLLRxDI(59));
  CNStageIntLLRInputS0xD(361)(0) <= LUT_4bit_to_3bit(ChLLRxDI(59));
  CNStageIntLLRInputS0xD(96)(0) <= LUT_4bit_to_3bit(ChLLRxDI(60));
  CNStageIntLLRInputS0xD(143)(0) <= LUT_4bit_to_3bit(ChLLRxDI(60));
  CNStageIntLLRInputS0xD(173)(0) <= LUT_4bit_to_3bit(ChLLRxDI(60));
  CNStageIntLLRInputS0xD(244)(0) <= LUT_4bit_to_3bit(ChLLRxDI(60));
  CNStageIntLLRInputS0xD(310)(0) <= LUT_4bit_to_3bit(ChLLRxDI(60));
  CNStageIntLLRInputS0xD(360)(0) <= LUT_4bit_to_3bit(ChLLRxDI(60));
  CNStageIntLLRInputS0xD(95)(0) <= LUT_4bit_to_3bit(ChLLRxDI(61));
  CNStageIntLLRInputS0xD(142)(0) <= LUT_4bit_to_3bit(ChLLRxDI(61));
  CNStageIntLLRInputS0xD(172)(0) <= LUT_4bit_to_3bit(ChLLRxDI(61));
  CNStageIntLLRInputS0xD(243)(0) <= LUT_4bit_to_3bit(ChLLRxDI(61));
  CNStageIntLLRInputS0xD(309)(0) <= LUT_4bit_to_3bit(ChLLRxDI(61));
  CNStageIntLLRInputS0xD(359)(0) <= LUT_4bit_to_3bit(ChLLRxDI(61));
  CNStageIntLLRInputS0xD(94)(0) <= LUT_4bit_to_3bit(ChLLRxDI(62));
  CNStageIntLLRInputS0xD(141)(0) <= LUT_4bit_to_3bit(ChLLRxDI(62));
  CNStageIntLLRInputS0xD(171)(0) <= LUT_4bit_to_3bit(ChLLRxDI(62));
  CNStageIntLLRInputS0xD(242)(0) <= LUT_4bit_to_3bit(ChLLRxDI(62));
  CNStageIntLLRInputS0xD(308)(0) <= LUT_4bit_to_3bit(ChLLRxDI(62));
  CNStageIntLLRInputS0xD(358)(0) <= LUT_4bit_to_3bit(ChLLRxDI(62));
  CNStageIntLLRInputS0xD(52)(0) <= LUT_4bit_to_3bit(ChLLRxDI(63));
  CNStageIntLLRInputS0xD(93)(0) <= LUT_4bit_to_3bit(ChLLRxDI(63));
  CNStageIntLLRInputS0xD(140)(0) <= LUT_4bit_to_3bit(ChLLRxDI(63));
  CNStageIntLLRInputS0xD(357)(0) <= LUT_4bit_to_3bit(ChLLRxDI(63));
  CNStageIntLLRInputS0xD(53)(1) <= LUT_4bit_to_3bit(ChLLRxDI(64));
  CNStageIntLLRInputS0xD(109)(1) <= LUT_4bit_to_3bit(ChLLRxDI(64));
  CNStageIntLLRInputS0xD(130)(1) <= LUT_4bit_to_3bit(ChLLRxDI(64));
  CNStageIntLLRInputS0xD(245)(1) <= LUT_4bit_to_3bit(ChLLRxDI(64));
  CNStageIntLLRInputS0xD(299)(1) <= LUT_4bit_to_3bit(ChLLRxDI(64));
  CNStageIntLLRInputS0xD(342)(1) <= LUT_4bit_to_3bit(ChLLRxDI(64));
  CNStageIntLLRInputS0xD(51)(1) <= LUT_4bit_to_3bit(ChLLRxDI(65));
  CNStageIntLLRInputS0xD(74)(1) <= LUT_4bit_to_3bit(ChLLRxDI(65));
  CNStageIntLLRInputS0xD(141)(1) <= LUT_4bit_to_3bit(ChLLRxDI(65));
  CNStageIntLLRInputS0xD(189)(1) <= LUT_4bit_to_3bit(ChLLRxDI(65));
  CNStageIntLLRInputS0xD(286)(1) <= LUT_4bit_to_3bit(ChLLRxDI(65));
  CNStageIntLLRInputS0xD(50)(1) <= LUT_4bit_to_3bit(ChLLRxDI(66));
  CNStageIntLLRInputS0xD(66)(1) <= LUT_4bit_to_3bit(ChLLRxDI(66));
  CNStageIntLLRInputS0xD(155)(1) <= LUT_4bit_to_3bit(ChLLRxDI(66));
  CNStageIntLLRInputS0xD(244)(1) <= LUT_4bit_to_3bit(ChLLRxDI(66));
  CNStageIntLLRInputS0xD(97)(1) <= LUT_4bit_to_3bit(ChLLRxDI(67));
  CNStageIntLLRInputS0xD(275)(1) <= LUT_4bit_to_3bit(ChLLRxDI(67));
  CNStageIntLLRInputS0xD(322)(1) <= LUT_4bit_to_3bit(ChLLRxDI(67));
  CNStageIntLLRInputS0xD(365)(1) <= LUT_4bit_to_3bit(ChLLRxDI(67));
  CNStageIntLLRInputS0xD(49)(1) <= LUT_4bit_to_3bit(ChLLRxDI(68));
  CNStageIntLLRInputS0xD(112)(1) <= LUT_4bit_to_3bit(ChLLRxDI(68));
  CNStageIntLLRInputS0xD(210)(1) <= LUT_4bit_to_3bit(ChLLRxDI(68));
  CNStageIntLLRInputS0xD(256)(1) <= LUT_4bit_to_3bit(ChLLRxDI(68));
  CNStageIntLLRInputS0xD(318)(1) <= LUT_4bit_to_3bit(ChLLRxDI(68));
  CNStageIntLLRInputS0xD(381)(1) <= LUT_4bit_to_3bit(ChLLRxDI(68));
  CNStageIntLLRInputS0xD(48)(1) <= LUT_4bit_to_3bit(ChLLRxDI(69));
  CNStageIntLLRInputS0xD(101)(1) <= LUT_4bit_to_3bit(ChLLRxDI(69));
  CNStageIntLLRInputS0xD(135)(1) <= LUT_4bit_to_3bit(ChLLRxDI(69));
  CNStageIntLLRInputS0xD(215)(1) <= LUT_4bit_to_3bit(ChLLRxDI(69));
  CNStageIntLLRInputS0xD(259)(1) <= LUT_4bit_to_3bit(ChLLRxDI(69));
  CNStageIntLLRInputS0xD(283)(1) <= LUT_4bit_to_3bit(ChLLRxDI(69));
  CNStageIntLLRInputS0xD(351)(1) <= LUT_4bit_to_3bit(ChLLRxDI(69));
  CNStageIntLLRInputS0xD(47)(1) <= LUT_4bit_to_3bit(ChLLRxDI(70));
  CNStageIntLLRInputS0xD(104)(1) <= LUT_4bit_to_3bit(ChLLRxDI(70));
  CNStageIntLLRInputS0xD(136)(1) <= LUT_4bit_to_3bit(ChLLRxDI(70));
  CNStageIntLLRInputS0xD(206)(1) <= LUT_4bit_to_3bit(ChLLRxDI(70));
  CNStageIntLLRInputS0xD(246)(1) <= LUT_4bit_to_3bit(ChLLRxDI(70));
  CNStageIntLLRInputS0xD(301)(1) <= LUT_4bit_to_3bit(ChLLRxDI(70));
  CNStageIntLLRInputS0xD(46)(1) <= LUT_4bit_to_3bit(ChLLRxDI(71));
  CNStageIntLLRInputS0xD(95)(1) <= LUT_4bit_to_3bit(ChLLRxDI(71));
  CNStageIntLLRInputS0xD(176)(1) <= LUT_4bit_to_3bit(ChLLRxDI(71));
  CNStageIntLLRInputS0xD(276)(1) <= LUT_4bit_to_3bit(ChLLRxDI(71));
  CNStageIntLLRInputS0xD(302)(1) <= LUT_4bit_to_3bit(ChLLRxDI(71));
  CNStageIntLLRInputS0xD(353)(1) <= LUT_4bit_to_3bit(ChLLRxDI(71));
  CNStageIntLLRInputS0xD(45)(1) <= LUT_4bit_to_3bit(ChLLRxDI(72));
  CNStageIntLLRInputS0xD(75)(1) <= LUT_4bit_to_3bit(ChLLRxDI(72));
  CNStageIntLLRInputS0xD(162)(1) <= LUT_4bit_to_3bit(ChLLRxDI(72));
  CNStageIntLLRInputS0xD(183)(1) <= LUT_4bit_to_3bit(ChLLRxDI(72));
  CNStageIntLLRInputS0xD(243)(1) <= LUT_4bit_to_3bit(ChLLRxDI(72));
  CNStageIntLLRInputS0xD(367)(1) <= LUT_4bit_to_3bit(ChLLRxDI(72));
  CNStageIntLLRInputS0xD(44)(1) <= LUT_4bit_to_3bit(ChLLRxDI(73));
  CNStageIntLLRInputS0xD(56)(1) <= LUT_4bit_to_3bit(ChLLRxDI(73));
  CNStageIntLLRInputS0xD(121)(1) <= LUT_4bit_to_3bit(ChLLRxDI(73));
  CNStageIntLLRInputS0xD(219)(1) <= LUT_4bit_to_3bit(ChLLRxDI(73));
  CNStageIntLLRInputS0xD(328)(1) <= LUT_4bit_to_3bit(ChLLRxDI(73));
  CNStageIntLLRInputS0xD(363)(1) <= LUT_4bit_to_3bit(ChLLRxDI(73));
  CNStageIntLLRInputS0xD(43)(1) <= LUT_4bit_to_3bit(ChLLRxDI(74));
  CNStageIntLLRInputS0xD(70)(1) <= LUT_4bit_to_3bit(ChLLRxDI(74));
  CNStageIntLLRInputS0xD(125)(1) <= LUT_4bit_to_3bit(ChLLRxDI(74));
  CNStageIntLLRInputS0xD(221)(1) <= LUT_4bit_to_3bit(ChLLRxDI(74));
  CNStageIntLLRInputS0xD(290)(1) <= LUT_4bit_to_3bit(ChLLRxDI(74));
  CNStageIntLLRInputS0xD(42)(1) <= LUT_4bit_to_3bit(ChLLRxDI(75));
  CNStageIntLLRInputS0xD(81)(1) <= LUT_4bit_to_3bit(ChLLRxDI(75));
  CNStageIntLLRInputS0xD(170)(1) <= LUT_4bit_to_3bit(ChLLRxDI(75));
  CNStageIntLLRInputS0xD(192)(1) <= LUT_4bit_to_3bit(ChLLRxDI(75));
  CNStageIntLLRInputS0xD(278)(1) <= LUT_4bit_to_3bit(ChLLRxDI(75));
  CNStageIntLLRInputS0xD(294)(1) <= LUT_4bit_to_3bit(ChLLRxDI(75));
  CNStageIntLLRInputS0xD(347)(1) <= LUT_4bit_to_3bit(ChLLRxDI(75));
  CNStageIntLLRInputS0xD(41)(1) <= LUT_4bit_to_3bit(ChLLRxDI(76));
  CNStageIntLLRInputS0xD(106)(1) <= LUT_4bit_to_3bit(ChLLRxDI(76));
  CNStageIntLLRInputS0xD(124)(1) <= LUT_4bit_to_3bit(ChLLRxDI(76));
  CNStageIntLLRInputS0xD(174)(1) <= LUT_4bit_to_3bit(ChLLRxDI(76));
  CNStageIntLLRInputS0xD(270)(1) <= LUT_4bit_to_3bit(ChLLRxDI(76));
  CNStageIntLLRInputS0xD(332)(1) <= LUT_4bit_to_3bit(ChLLRxDI(76));
  CNStageIntLLRInputS0xD(348)(1) <= LUT_4bit_to_3bit(ChLLRxDI(76));
  CNStageIntLLRInputS0xD(119)(1) <= LUT_4bit_to_3bit(ChLLRxDI(77));
  CNStageIntLLRInputS0xD(185)(1) <= LUT_4bit_to_3bit(ChLLRxDI(77));
  CNStageIntLLRInputS0xD(257)(1) <= LUT_4bit_to_3bit(ChLLRxDI(77));
  CNStageIntLLRInputS0xD(293)(1) <= LUT_4bit_to_3bit(ChLLRxDI(77));
  CNStageIntLLRInputS0xD(383)(1) <= LUT_4bit_to_3bit(ChLLRxDI(77));
  CNStageIntLLRInputS0xD(40)(1) <= LUT_4bit_to_3bit(ChLLRxDI(78));
  CNStageIntLLRInputS0xD(84)(1) <= LUT_4bit_to_3bit(ChLLRxDI(78));
  CNStageIntLLRInputS0xD(159)(1) <= LUT_4bit_to_3bit(ChLLRxDI(78));
  CNStageIntLLRInputS0xD(193)(1) <= LUT_4bit_to_3bit(ChLLRxDI(78));
  CNStageIntLLRInputS0xD(274)(1) <= LUT_4bit_to_3bit(ChLLRxDI(78));
  CNStageIntLLRInputS0xD(288)(1) <= LUT_4bit_to_3bit(ChLLRxDI(78));
  CNStageIntLLRInputS0xD(374)(1) <= LUT_4bit_to_3bit(ChLLRxDI(78));
  CNStageIntLLRInputS0xD(39)(1) <= LUT_4bit_to_3bit(ChLLRxDI(79));
  CNStageIntLLRInputS0xD(99)(1) <= LUT_4bit_to_3bit(ChLLRxDI(79));
  CNStageIntLLRInputS0xD(167)(1) <= LUT_4bit_to_3bit(ChLLRxDI(79));
  CNStageIntLLRInputS0xD(220)(1) <= LUT_4bit_to_3bit(ChLLRxDI(79));
  CNStageIntLLRInputS0xD(325)(1) <= LUT_4bit_to_3bit(ChLLRxDI(79));
  CNStageIntLLRInputS0xD(38)(1) <= LUT_4bit_to_3bit(ChLLRxDI(80));
  CNStageIntLLRInputS0xD(62)(1) <= LUT_4bit_to_3bit(ChLLRxDI(80));
  CNStageIntLLRInputS0xD(131)(1) <= LUT_4bit_to_3bit(ChLLRxDI(80));
  CNStageIntLLRInputS0xD(182)(1) <= LUT_4bit_to_3bit(ChLLRxDI(80));
  CNStageIntLLRInputS0xD(248)(1) <= LUT_4bit_to_3bit(ChLLRxDI(80));
  CNStageIntLLRInputS0xD(337)(1) <= LUT_4bit_to_3bit(ChLLRxDI(80));
  CNStageIntLLRInputS0xD(37)(1) <= LUT_4bit_to_3bit(ChLLRxDI(81));
  CNStageIntLLRInputS0xD(72)(1) <= LUT_4bit_to_3bit(ChLLRxDI(81));
  CNStageIntLLRInputS0xD(129)(1) <= LUT_4bit_to_3bit(ChLLRxDI(81));
  CNStageIntLLRInputS0xD(262)(1) <= LUT_4bit_to_3bit(ChLLRxDI(81));
  CNStageIntLLRInputS0xD(36)(1) <= LUT_4bit_to_3bit(ChLLRxDI(82));
  CNStageIntLLRInputS0xD(67)(1) <= LUT_4bit_to_3bit(ChLLRxDI(82));
  CNStageIntLLRInputS0xD(165)(1) <= LUT_4bit_to_3bit(ChLLRxDI(82));
  CNStageIntLLRInputS0xD(188)(1) <= LUT_4bit_to_3bit(ChLLRxDI(82));
  CNStageIntLLRInputS0xD(254)(1) <= LUT_4bit_to_3bit(ChLLRxDI(82));
  CNStageIntLLRInputS0xD(298)(1) <= LUT_4bit_to_3bit(ChLLRxDI(82));
  CNStageIntLLRInputS0xD(336)(1) <= LUT_4bit_to_3bit(ChLLRxDI(82));
  CNStageIntLLRInputS0xD(35)(1) <= LUT_4bit_to_3bit(ChLLRxDI(83));
  CNStageIntLLRInputS0xD(73)(1) <= LUT_4bit_to_3bit(ChLLRxDI(83));
  CNStageIntLLRInputS0xD(144)(1) <= LUT_4bit_to_3bit(ChLLRxDI(83));
  CNStageIntLLRInputS0xD(208)(1) <= LUT_4bit_to_3bit(ChLLRxDI(83));
  CNStageIntLLRInputS0xD(232)(1) <= LUT_4bit_to_3bit(ChLLRxDI(83));
  CNStageIntLLRInputS0xD(330)(1) <= LUT_4bit_to_3bit(ChLLRxDI(83));
  CNStageIntLLRInputS0xD(34)(1) <= LUT_4bit_to_3bit(ChLLRxDI(84));
  CNStageIntLLRInputS0xD(61)(1) <= LUT_4bit_to_3bit(ChLLRxDI(84));
  CNStageIntLLRInputS0xD(147)(1) <= LUT_4bit_to_3bit(ChLLRxDI(84));
  CNStageIntLLRInputS0xD(222)(1) <= LUT_4bit_to_3bit(ChLLRxDI(84));
  CNStageIntLLRInputS0xD(310)(1) <= LUT_4bit_to_3bit(ChLLRxDI(84));
  CNStageIntLLRInputS0xD(371)(1) <= LUT_4bit_to_3bit(ChLLRxDI(84));
  CNStageIntLLRInputS0xD(33)(1) <= LUT_4bit_to_3bit(ChLLRxDI(85));
  CNStageIntLLRInputS0xD(132)(1) <= LUT_4bit_to_3bit(ChLLRxDI(85));
  CNStageIntLLRInputS0xD(218)(1) <= LUT_4bit_to_3bit(ChLLRxDI(85));
  CNStageIntLLRInputS0xD(235)(1) <= LUT_4bit_to_3bit(ChLLRxDI(85));
  CNStageIntLLRInputS0xD(313)(1) <= LUT_4bit_to_3bit(ChLLRxDI(85));
  CNStageIntLLRInputS0xD(379)(1) <= LUT_4bit_to_3bit(ChLLRxDI(85));
  CNStageIntLLRInputS0xD(32)(1) <= LUT_4bit_to_3bit(ChLLRxDI(86));
  CNStageIntLLRInputS0xD(166)(1) <= LUT_4bit_to_3bit(ChLLRxDI(86));
  CNStageIntLLRInputS0xD(239)(1) <= LUT_4bit_to_3bit(ChLLRxDI(86));
  CNStageIntLLRInputS0xD(343)(1) <= LUT_4bit_to_3bit(ChLLRxDI(86));
  CNStageIntLLRInputS0xD(31)(1) <= LUT_4bit_to_3bit(ChLLRxDI(87));
  CNStageIntLLRInputS0xD(77)(1) <= LUT_4bit_to_3bit(ChLLRxDI(87));
  CNStageIntLLRInputS0xD(128)(1) <= LUT_4bit_to_3bit(ChLLRxDI(87));
  CNStageIntLLRInputS0xD(203)(1) <= LUT_4bit_to_3bit(ChLLRxDI(87));
  CNStageIntLLRInputS0xD(229)(1) <= LUT_4bit_to_3bit(ChLLRxDI(87));
  CNStageIntLLRInputS0xD(331)(1) <= LUT_4bit_to_3bit(ChLLRxDI(87));
  CNStageIntLLRInputS0xD(341)(1) <= LUT_4bit_to_3bit(ChLLRxDI(87));
  CNStageIntLLRInputS0xD(30)(1) <= LUT_4bit_to_3bit(ChLLRxDI(88));
  CNStageIntLLRInputS0xD(79)(1) <= LUT_4bit_to_3bit(ChLLRxDI(88));
  CNStageIntLLRInputS0xD(156)(1) <= LUT_4bit_to_3bit(ChLLRxDI(88));
  CNStageIntLLRInputS0xD(204)(1) <= LUT_4bit_to_3bit(ChLLRxDI(88));
  CNStageIntLLRInputS0xD(263)(1) <= LUT_4bit_to_3bit(ChLLRxDI(88));
  CNStageIntLLRInputS0xD(297)(1) <= LUT_4bit_to_3bit(ChLLRxDI(88));
  CNStageIntLLRInputS0xD(377)(1) <= LUT_4bit_to_3bit(ChLLRxDI(88));
  CNStageIntLLRInputS0xD(29)(1) <= LUT_4bit_to_3bit(ChLLRxDI(89));
  CNStageIntLLRInputS0xD(102)(1) <= LUT_4bit_to_3bit(ChLLRxDI(89));
  CNStageIntLLRInputS0xD(140)(1) <= LUT_4bit_to_3bit(ChLLRxDI(89));
  CNStageIntLLRInputS0xD(184)(1) <= LUT_4bit_to_3bit(ChLLRxDI(89));
  CNStageIntLLRInputS0xD(247)(1) <= LUT_4bit_to_3bit(ChLLRxDI(89));
  CNStageIntLLRInputS0xD(355)(1) <= LUT_4bit_to_3bit(ChLLRxDI(89));
  CNStageIntLLRInputS0xD(28)(1) <= LUT_4bit_to_3bit(ChLLRxDI(90));
  CNStageIntLLRInputS0xD(85)(1) <= LUT_4bit_to_3bit(ChLLRxDI(90));
  CNStageIntLLRInputS0xD(168)(1) <= LUT_4bit_to_3bit(ChLLRxDI(90));
  CNStageIntLLRInputS0xD(175)(1) <= LUT_4bit_to_3bit(ChLLRxDI(90));
  CNStageIntLLRInputS0xD(258)(1) <= LUT_4bit_to_3bit(ChLLRxDI(90));
  CNStageIntLLRInputS0xD(307)(1) <= LUT_4bit_to_3bit(ChLLRxDI(90));
  CNStageIntLLRInputS0xD(358)(1) <= LUT_4bit_to_3bit(ChLLRxDI(90));
  CNStageIntLLRInputS0xD(27)(1) <= LUT_4bit_to_3bit(ChLLRxDI(91));
  CNStageIntLLRInputS0xD(96)(1) <= LUT_4bit_to_3bit(ChLLRxDI(91));
  CNStageIntLLRInputS0xD(158)(1) <= LUT_4bit_to_3bit(ChLLRxDI(91));
  CNStageIntLLRInputS0xD(191)(1) <= LUT_4bit_to_3bit(ChLLRxDI(91));
  CNStageIntLLRInputS0xD(269)(1) <= LUT_4bit_to_3bit(ChLLRxDI(91));
  CNStageIntLLRInputS0xD(280)(1) <= LUT_4bit_to_3bit(ChLLRxDI(91));
  CNStageIntLLRInputS0xD(344)(1) <= LUT_4bit_to_3bit(ChLLRxDI(91));
  CNStageIntLLRInputS0xD(26)(1) <= LUT_4bit_to_3bit(ChLLRxDI(92));
  CNStageIntLLRInputS0xD(103)(1) <= LUT_4bit_to_3bit(ChLLRxDI(92));
  CNStageIntLLRInputS0xD(145)(1) <= LUT_4bit_to_3bit(ChLLRxDI(92));
  CNStageIntLLRInputS0xD(195)(1) <= LUT_4bit_to_3bit(ChLLRxDI(92));
  CNStageIntLLRInputS0xD(242)(1) <= LUT_4bit_to_3bit(ChLLRxDI(92));
  CNStageIntLLRInputS0xD(324)(1) <= LUT_4bit_to_3bit(ChLLRxDI(92));
  CNStageIntLLRInputS0xD(378)(1) <= LUT_4bit_to_3bit(ChLLRxDI(92));
  CNStageIntLLRInputS0xD(25)(1) <= LUT_4bit_to_3bit(ChLLRxDI(93));
  CNStageIntLLRInputS0xD(78)(1) <= LUT_4bit_to_3bit(ChLLRxDI(93));
  CNStageIntLLRInputS0xD(164)(1) <= LUT_4bit_to_3bit(ChLLRxDI(93));
  CNStageIntLLRInputS0xD(224)(1) <= LUT_4bit_to_3bit(ChLLRxDI(93));
  CNStageIntLLRInputS0xD(231)(1) <= LUT_4bit_to_3bit(ChLLRxDI(93));
  CNStageIntLLRInputS0xD(311)(1) <= LUT_4bit_to_3bit(ChLLRxDI(93));
  CNStageIntLLRInputS0xD(340)(1) <= LUT_4bit_to_3bit(ChLLRxDI(93));
  CNStageIntLLRInputS0xD(24)(1) <= LUT_4bit_to_3bit(ChLLRxDI(94));
  CNStageIntLLRInputS0xD(92)(1) <= LUT_4bit_to_3bit(ChLLRxDI(94));
  CNStageIntLLRInputS0xD(194)(1) <= LUT_4bit_to_3bit(ChLLRxDI(94));
  CNStageIntLLRInputS0xD(329)(1) <= LUT_4bit_to_3bit(ChLLRxDI(94));
  CNStageIntLLRInputS0xD(368)(1) <= LUT_4bit_to_3bit(ChLLRxDI(94));
  CNStageIntLLRInputS0xD(23)(1) <= LUT_4bit_to_3bit(ChLLRxDI(95));
  CNStageIntLLRInputS0xD(63)(1) <= LUT_4bit_to_3bit(ChLLRxDI(95));
  CNStageIntLLRInputS0xD(134)(1) <= LUT_4bit_to_3bit(ChLLRxDI(95));
  CNStageIntLLRInputS0xD(190)(1) <= LUT_4bit_to_3bit(ChLLRxDI(95));
  CNStageIntLLRInputS0xD(234)(1) <= LUT_4bit_to_3bit(ChLLRxDI(95));
  CNStageIntLLRInputS0xD(303)(1) <= LUT_4bit_to_3bit(ChLLRxDI(95));
  CNStageIntLLRInputS0xD(352)(1) <= LUT_4bit_to_3bit(ChLLRxDI(95));
  CNStageIntLLRInputS0xD(22)(1) <= LUT_4bit_to_3bit(ChLLRxDI(96));
  CNStageIntLLRInputS0xD(98)(1) <= LUT_4bit_to_3bit(ChLLRxDI(96));
  CNStageIntLLRInputS0xD(150)(1) <= LUT_4bit_to_3bit(ChLLRxDI(96));
  CNStageIntLLRInputS0xD(172)(1) <= LUT_4bit_to_3bit(ChLLRxDI(96));
  CNStageIntLLRInputS0xD(251)(1) <= LUT_4bit_to_3bit(ChLLRxDI(96));
  CNStageIntLLRInputS0xD(380)(1) <= LUT_4bit_to_3bit(ChLLRxDI(96));
  CNStageIntLLRInputS0xD(21)(1) <= LUT_4bit_to_3bit(ChLLRxDI(97));
  CNStageIntLLRInputS0xD(65)(1) <= LUT_4bit_to_3bit(ChLLRxDI(97));
  CNStageIntLLRInputS0xD(142)(1) <= LUT_4bit_to_3bit(ChLLRxDI(97));
  CNStageIntLLRInputS0xD(180)(1) <= LUT_4bit_to_3bit(ChLLRxDI(97));
  CNStageIntLLRInputS0xD(260)(1) <= LUT_4bit_to_3bit(ChLLRxDI(97));
  CNStageIntLLRInputS0xD(316)(1) <= LUT_4bit_to_3bit(ChLLRxDI(97));
  CNStageIntLLRInputS0xD(370)(1) <= LUT_4bit_to_3bit(ChLLRxDI(97));
  CNStageIntLLRInputS0xD(20)(1) <= LUT_4bit_to_3bit(ChLLRxDI(98));
  CNStageIntLLRInputS0xD(116)(1) <= LUT_4bit_to_3bit(ChLLRxDI(98));
  CNStageIntLLRInputS0xD(199)(1) <= LUT_4bit_to_3bit(ChLLRxDI(98));
  CNStageIntLLRInputS0xD(255)(1) <= LUT_4bit_to_3bit(ChLLRxDI(98));
  CNStageIntLLRInputS0xD(308)(1) <= LUT_4bit_to_3bit(ChLLRxDI(98));
  CNStageIntLLRInputS0xD(356)(1) <= LUT_4bit_to_3bit(ChLLRxDI(98));
  CNStageIntLLRInputS0xD(19)(1) <= LUT_4bit_to_3bit(ChLLRxDI(99));
  CNStageIntLLRInputS0xD(76)(1) <= LUT_4bit_to_3bit(ChLLRxDI(99));
  CNStageIntLLRInputS0xD(126)(1) <= LUT_4bit_to_3bit(ChLLRxDI(99));
  CNStageIntLLRInputS0xD(198)(1) <= LUT_4bit_to_3bit(ChLLRxDI(99));
  CNStageIntLLRInputS0xD(261)(1) <= LUT_4bit_to_3bit(ChLLRxDI(99));
  CNStageIntLLRInputS0xD(285)(1) <= LUT_4bit_to_3bit(ChLLRxDI(99));
  CNStageIntLLRInputS0xD(376)(1) <= LUT_4bit_to_3bit(ChLLRxDI(99));
  CNStageIntLLRInputS0xD(18)(1) <= LUT_4bit_to_3bit(ChLLRxDI(100));
  CNStageIntLLRInputS0xD(94)(1) <= LUT_4bit_to_3bit(ChLLRxDI(100));
  CNStageIntLLRInputS0xD(120)(1) <= LUT_4bit_to_3bit(ChLLRxDI(100));
  CNStageIntLLRInputS0xD(178)(1) <= LUT_4bit_to_3bit(ChLLRxDI(100));
  CNStageIntLLRInputS0xD(250)(1) <= LUT_4bit_to_3bit(ChLLRxDI(100));
  CNStageIntLLRInputS0xD(295)(1) <= LUT_4bit_to_3bit(ChLLRxDI(100));
  CNStageIntLLRInputS0xD(349)(1) <= LUT_4bit_to_3bit(ChLLRxDI(100));
  CNStageIntLLRInputS0xD(17)(1) <= LUT_4bit_to_3bit(ChLLRxDI(101));
  CNStageIntLLRInputS0xD(58)(1) <= LUT_4bit_to_3bit(ChLLRxDI(101));
  CNStageIntLLRInputS0xD(123)(1) <= LUT_4bit_to_3bit(ChLLRxDI(101));
  CNStageIntLLRInputS0xD(211)(1) <= LUT_4bit_to_3bit(ChLLRxDI(101));
  CNStageIntLLRInputS0xD(273)(1) <= LUT_4bit_to_3bit(ChLLRxDI(101));
  CNStageIntLLRInputS0xD(289)(1) <= LUT_4bit_to_3bit(ChLLRxDI(101));
  CNStageIntLLRInputS0xD(346)(1) <= LUT_4bit_to_3bit(ChLLRxDI(101));
  CNStageIntLLRInputS0xD(16)(1) <= LUT_4bit_to_3bit(ChLLRxDI(102));
  CNStageIntLLRInputS0xD(59)(1) <= LUT_4bit_to_3bit(ChLLRxDI(102));
  CNStageIntLLRInputS0xD(113)(1) <= LUT_4bit_to_3bit(ChLLRxDI(102));
  CNStageIntLLRInputS0xD(214)(1) <= LUT_4bit_to_3bit(ChLLRxDI(102));
  CNStageIntLLRInputS0xD(226)(1) <= LUT_4bit_to_3bit(ChLLRxDI(102));
  CNStageIntLLRInputS0xD(361)(1) <= LUT_4bit_to_3bit(ChLLRxDI(102));
  CNStageIntLLRInputS0xD(15)(1) <= LUT_4bit_to_3bit(ChLLRxDI(103));
  CNStageIntLLRInputS0xD(93)(1) <= LUT_4bit_to_3bit(ChLLRxDI(103));
  CNStageIntLLRInputS0xD(151)(1) <= LUT_4bit_to_3bit(ChLLRxDI(103));
  CNStageIntLLRInputS0xD(200)(1) <= LUT_4bit_to_3bit(ChLLRxDI(103));
  CNStageIntLLRInputS0xD(265)(1) <= LUT_4bit_to_3bit(ChLLRxDI(103));
  CNStageIntLLRInputS0xD(284)(1) <= LUT_4bit_to_3bit(ChLLRxDI(103));
  CNStageIntLLRInputS0xD(354)(1) <= LUT_4bit_to_3bit(ChLLRxDI(103));
  CNStageIntLLRInputS0xD(14)(1) <= LUT_4bit_to_3bit(ChLLRxDI(104));
  CNStageIntLLRInputS0xD(86)(1) <= LUT_4bit_to_3bit(ChLLRxDI(104));
  CNStageIntLLRInputS0xD(133)(1) <= LUT_4bit_to_3bit(ChLLRxDI(104));
  CNStageIntLLRInputS0xD(179)(1) <= LUT_4bit_to_3bit(ChLLRxDI(104));
  CNStageIntLLRInputS0xD(267)(1) <= LUT_4bit_to_3bit(ChLLRxDI(104));
  CNStageIntLLRInputS0xD(317)(1) <= LUT_4bit_to_3bit(ChLLRxDI(104));
  CNStageIntLLRInputS0xD(13)(1) <= LUT_4bit_to_3bit(ChLLRxDI(105));
  CNStageIntLLRInputS0xD(146)(1) <= LUT_4bit_to_3bit(ChLLRxDI(105));
  CNStageIntLLRInputS0xD(197)(1) <= LUT_4bit_to_3bit(ChLLRxDI(105));
  CNStageIntLLRInputS0xD(237)(1) <= LUT_4bit_to_3bit(ChLLRxDI(105));
  CNStageIntLLRInputS0xD(300)(1) <= LUT_4bit_to_3bit(ChLLRxDI(105));
  CNStageIntLLRInputS0xD(338)(1) <= LUT_4bit_to_3bit(ChLLRxDI(105));
  CNStageIntLLRInputS0xD(12)(1) <= LUT_4bit_to_3bit(ChLLRxDI(106));
  CNStageIntLLRInputS0xD(157)(1) <= LUT_4bit_to_3bit(ChLLRxDI(106));
  CNStageIntLLRInputS0xD(223)(1) <= LUT_4bit_to_3bit(ChLLRxDI(106));
  CNStageIntLLRInputS0xD(272)(1) <= LUT_4bit_to_3bit(ChLLRxDI(106));
  CNStageIntLLRInputS0xD(312)(1) <= LUT_4bit_to_3bit(ChLLRxDI(106));
  CNStageIntLLRInputS0xD(333)(1) <= LUT_4bit_to_3bit(ChLLRxDI(106));
  CNStageIntLLRInputS0xD(110)(1) <= LUT_4bit_to_3bit(ChLLRxDI(107));
  CNStageIntLLRInputS0xD(127)(1) <= LUT_4bit_to_3bit(ChLLRxDI(107));
  CNStageIntLLRInputS0xD(207)(1) <= LUT_4bit_to_3bit(ChLLRxDI(107));
  CNStageIntLLRInputS0xD(230)(1) <= LUT_4bit_to_3bit(ChLLRxDI(107));
  CNStageIntLLRInputS0xD(323)(1) <= LUT_4bit_to_3bit(ChLLRxDI(107));
  CNStageIntLLRInputS0xD(335)(1) <= LUT_4bit_to_3bit(ChLLRxDI(107));
  CNStageIntLLRInputS0xD(11)(1) <= LUT_4bit_to_3bit(ChLLRxDI(108));
  CNStageIntLLRInputS0xD(105)(1) <= LUT_4bit_to_3bit(ChLLRxDI(108));
  CNStageIntLLRInputS0xD(115)(1) <= LUT_4bit_to_3bit(ChLLRxDI(108));
  CNStageIntLLRInputS0xD(181)(1) <= LUT_4bit_to_3bit(ChLLRxDI(108));
  CNStageIntLLRInputS0xD(238)(1) <= LUT_4bit_to_3bit(ChLLRxDI(108));
  CNStageIntLLRInputS0xD(296)(1) <= LUT_4bit_to_3bit(ChLLRxDI(108));
  CNStageIntLLRInputS0xD(10)(1) <= LUT_4bit_to_3bit(ChLLRxDI(109));
  CNStageIntLLRInputS0xD(100)(1) <= LUT_4bit_to_3bit(ChLLRxDI(109));
  CNStageIntLLRInputS0xD(160)(1) <= LUT_4bit_to_3bit(ChLLRxDI(109));
  CNStageIntLLRInputS0xD(171)(1) <= LUT_4bit_to_3bit(ChLLRxDI(109));
  CNStageIntLLRInputS0xD(266)(1) <= LUT_4bit_to_3bit(ChLLRxDI(109));
  CNStageIntLLRInputS0xD(362)(1) <= LUT_4bit_to_3bit(ChLLRxDI(109));
  CNStageIntLLRInputS0xD(9)(1) <= LUT_4bit_to_3bit(ChLLRxDI(110));
  CNStageIntLLRInputS0xD(83)(1) <= LUT_4bit_to_3bit(ChLLRxDI(110));
  CNStageIntLLRInputS0xD(118)(1) <= LUT_4bit_to_3bit(ChLLRxDI(110));
  CNStageIntLLRInputS0xD(212)(1) <= LUT_4bit_to_3bit(ChLLRxDI(110));
  CNStageIntLLRInputS0xD(225)(1) <= LUT_4bit_to_3bit(ChLLRxDI(110));
  CNStageIntLLRInputS0xD(326)(1) <= LUT_4bit_to_3bit(ChLLRxDI(110));
  CNStageIntLLRInputS0xD(345)(1) <= LUT_4bit_to_3bit(ChLLRxDI(110));
  CNStageIntLLRInputS0xD(8)(1) <= LUT_4bit_to_3bit(ChLLRxDI(111));
  CNStageIntLLRInputS0xD(90)(1) <= LUT_4bit_to_3bit(ChLLRxDI(111));
  CNStageIntLLRInputS0xD(138)(1) <= LUT_4bit_to_3bit(ChLLRxDI(111));
  CNStageIntLLRInputS0xD(177)(1) <= LUT_4bit_to_3bit(ChLLRxDI(111));
  CNStageIntLLRInputS0xD(252)(1) <= LUT_4bit_to_3bit(ChLLRxDI(111));
  CNStageIntLLRInputS0xD(287)(1) <= LUT_4bit_to_3bit(ChLLRxDI(111));
  CNStageIntLLRInputS0xD(357)(1) <= LUT_4bit_to_3bit(ChLLRxDI(111));
  CNStageIntLLRInputS0xD(7)(1) <= LUT_4bit_to_3bit(ChLLRxDI(112));
  CNStageIntLLRInputS0xD(54)(1) <= LUT_4bit_to_3bit(ChLLRxDI(112));
  CNStageIntLLRInputS0xD(148)(1) <= LUT_4bit_to_3bit(ChLLRxDI(112));
  CNStageIntLLRInputS0xD(205)(1) <= LUT_4bit_to_3bit(ChLLRxDI(112));
  CNStageIntLLRInputS0xD(233)(1) <= LUT_4bit_to_3bit(ChLLRxDI(112));
  CNStageIntLLRInputS0xD(305)(1) <= LUT_4bit_to_3bit(ChLLRxDI(112));
  CNStageIntLLRInputS0xD(369)(1) <= LUT_4bit_to_3bit(ChLLRxDI(112));
  CNStageIntLLRInputS0xD(6)(1) <= LUT_4bit_to_3bit(ChLLRxDI(113));
  CNStageIntLLRInputS0xD(108)(1) <= LUT_4bit_to_3bit(ChLLRxDI(113));
  CNStageIntLLRInputS0xD(143)(1) <= LUT_4bit_to_3bit(ChLLRxDI(113));
  CNStageIntLLRInputS0xD(202)(1) <= LUT_4bit_to_3bit(ChLLRxDI(113));
  CNStageIntLLRInputS0xD(253)(1) <= LUT_4bit_to_3bit(ChLLRxDI(113));
  CNStageIntLLRInputS0xD(314)(1) <= LUT_4bit_to_3bit(ChLLRxDI(113));
  CNStageIntLLRInputS0xD(339)(1) <= LUT_4bit_to_3bit(ChLLRxDI(113));
  CNStageIntLLRInputS0xD(5)(1) <= LUT_4bit_to_3bit(ChLLRxDI(114));
  CNStageIntLLRInputS0xD(88)(1) <= LUT_4bit_to_3bit(ChLLRxDI(114));
  CNStageIntLLRInputS0xD(149)(1) <= LUT_4bit_to_3bit(ChLLRxDI(114));
  CNStageIntLLRInputS0xD(216)(1) <= LUT_4bit_to_3bit(ChLLRxDI(114));
  CNStageIntLLRInputS0xD(268)(1) <= LUT_4bit_to_3bit(ChLLRxDI(114));
  CNStageIntLLRInputS0xD(309)(1) <= LUT_4bit_to_3bit(ChLLRxDI(114));
  CNStageIntLLRInputS0xD(4)(1) <= LUT_4bit_to_3bit(ChLLRxDI(115));
  CNStageIntLLRInputS0xD(68)(1) <= LUT_4bit_to_3bit(ChLLRxDI(115));
  CNStageIntLLRInputS0xD(137)(1) <= LUT_4bit_to_3bit(ChLLRxDI(115));
  CNStageIntLLRInputS0xD(209)(1) <= LUT_4bit_to_3bit(ChLLRxDI(115));
  CNStageIntLLRInputS0xD(264)(1) <= LUT_4bit_to_3bit(ChLLRxDI(115));
  CNStageIntLLRInputS0xD(315)(1) <= LUT_4bit_to_3bit(ChLLRxDI(115));
  CNStageIntLLRInputS0xD(372)(1) <= LUT_4bit_to_3bit(ChLLRxDI(115));
  CNStageIntLLRInputS0xD(71)(1) <= LUT_4bit_to_3bit(ChLLRxDI(116));
  CNStageIntLLRInputS0xD(163)(1) <= LUT_4bit_to_3bit(ChLLRxDI(116));
  CNStageIntLLRInputS0xD(187)(1) <= LUT_4bit_to_3bit(ChLLRxDI(116));
  CNStageIntLLRInputS0xD(228)(1) <= LUT_4bit_to_3bit(ChLLRxDI(116));
  CNStageIntLLRInputS0xD(304)(1) <= LUT_4bit_to_3bit(ChLLRxDI(116));
  CNStageIntLLRInputS0xD(3)(1) <= LUT_4bit_to_3bit(ChLLRxDI(117));
  CNStageIntLLRInputS0xD(55)(1) <= LUT_4bit_to_3bit(ChLLRxDI(117));
  CNStageIntLLRInputS0xD(111)(1) <= LUT_4bit_to_3bit(ChLLRxDI(117));
  CNStageIntLLRInputS0xD(196)(1) <= LUT_4bit_to_3bit(ChLLRxDI(117));
  CNStageIntLLRInputS0xD(2)(1) <= LUT_4bit_to_3bit(ChLLRxDI(118));
  CNStageIntLLRInputS0xD(89)(1) <= LUT_4bit_to_3bit(ChLLRxDI(118));
  CNStageIntLLRInputS0xD(152)(1) <= LUT_4bit_to_3bit(ChLLRxDI(118));
  CNStageIntLLRInputS0xD(249)(1) <= LUT_4bit_to_3bit(ChLLRxDI(118));
  CNStageIntLLRInputS0xD(282)(1) <= LUT_4bit_to_3bit(ChLLRxDI(118));
  CNStageIntLLRInputS0xD(359)(1) <= LUT_4bit_to_3bit(ChLLRxDI(118));
  CNStageIntLLRInputS0xD(1)(1) <= LUT_4bit_to_3bit(ChLLRxDI(119));
  CNStageIntLLRInputS0xD(107)(1) <= LUT_4bit_to_3bit(ChLLRxDI(119));
  CNStageIntLLRInputS0xD(154)(1) <= LUT_4bit_to_3bit(ChLLRxDI(119));
  CNStageIntLLRInputS0xD(227)(1) <= LUT_4bit_to_3bit(ChLLRxDI(119));
  CNStageIntLLRInputS0xD(319)(1) <= LUT_4bit_to_3bit(ChLLRxDI(119));
  CNStageIntLLRInputS0xD(0)(1) <= LUT_4bit_to_3bit(ChLLRxDI(120));
  CNStageIntLLRInputS0xD(80)(1) <= LUT_4bit_to_3bit(ChLLRxDI(120));
  CNStageIntLLRInputS0xD(321)(1) <= LUT_4bit_to_3bit(ChLLRxDI(120));
  CNStageIntLLRInputS0xD(360)(1) <= LUT_4bit_to_3bit(ChLLRxDI(120));
  CNStageIntLLRInputS0xD(64)(1) <= LUT_4bit_to_3bit(ChLLRxDI(121));
  CNStageIntLLRInputS0xD(161)(1) <= LUT_4bit_to_3bit(ChLLRxDI(121));
  CNStageIntLLRInputS0xD(217)(1) <= LUT_4bit_to_3bit(ChLLRxDI(121));
  CNStageIntLLRInputS0xD(236)(1) <= LUT_4bit_to_3bit(ChLLRxDI(121));
  CNStageIntLLRInputS0xD(291)(1) <= LUT_4bit_to_3bit(ChLLRxDI(121));
  CNStageIntLLRInputS0xD(350)(1) <= LUT_4bit_to_3bit(ChLLRxDI(121));
  CNStageIntLLRInputS0xD(91)(1) <= LUT_4bit_to_3bit(ChLLRxDI(122));
  CNStageIntLLRInputS0xD(114)(1) <= LUT_4bit_to_3bit(ChLLRxDI(122));
  CNStageIntLLRInputS0xD(201)(1) <= LUT_4bit_to_3bit(ChLLRxDI(122));
  CNStageIntLLRInputS0xD(241)(1) <= LUT_4bit_to_3bit(ChLLRxDI(122));
  CNStageIntLLRInputS0xD(327)(1) <= LUT_4bit_to_3bit(ChLLRxDI(122));
  CNStageIntLLRInputS0xD(375)(1) <= LUT_4bit_to_3bit(ChLLRxDI(122));
  CNStageIntLLRInputS0xD(82)(1) <= LUT_4bit_to_3bit(ChLLRxDI(123));
  CNStageIntLLRInputS0xD(122)(1) <= LUT_4bit_to_3bit(ChLLRxDI(123));
  CNStageIntLLRInputS0xD(213)(1) <= LUT_4bit_to_3bit(ChLLRxDI(123));
  CNStageIntLLRInputS0xD(279)(1) <= LUT_4bit_to_3bit(ChLLRxDI(123));
  CNStageIntLLRInputS0xD(382)(1) <= LUT_4bit_to_3bit(ChLLRxDI(123));
  CNStageIntLLRInputS0xD(69)(1) <= LUT_4bit_to_3bit(ChLLRxDI(124));
  CNStageIntLLRInputS0xD(153)(1) <= LUT_4bit_to_3bit(ChLLRxDI(124));
  CNStageIntLLRInputS0xD(240)(1) <= LUT_4bit_to_3bit(ChLLRxDI(124));
  CNStageIntLLRInputS0xD(292)(1) <= LUT_4bit_to_3bit(ChLLRxDI(124));
  CNStageIntLLRInputS0xD(364)(1) <= LUT_4bit_to_3bit(ChLLRxDI(124));
  CNStageIntLLRInputS0xD(87)(1) <= LUT_4bit_to_3bit(ChLLRxDI(125));
  CNStageIntLLRInputS0xD(169)(1) <= LUT_4bit_to_3bit(ChLLRxDI(125));
  CNStageIntLLRInputS0xD(320)(1) <= LUT_4bit_to_3bit(ChLLRxDI(125));
  CNStageIntLLRInputS0xD(366)(1) <= LUT_4bit_to_3bit(ChLLRxDI(125));
  CNStageIntLLRInputS0xD(60)(1) <= LUT_4bit_to_3bit(ChLLRxDI(126));
  CNStageIntLLRInputS0xD(139)(1) <= LUT_4bit_to_3bit(ChLLRxDI(126));
  CNStageIntLLRInputS0xD(186)(1) <= LUT_4bit_to_3bit(ChLLRxDI(126));
  CNStageIntLLRInputS0xD(271)(1) <= LUT_4bit_to_3bit(ChLLRxDI(126));
  CNStageIntLLRInputS0xD(281)(1) <= LUT_4bit_to_3bit(ChLLRxDI(126));
  CNStageIntLLRInputS0xD(334)(1) <= LUT_4bit_to_3bit(ChLLRxDI(126));
  CNStageIntLLRInputS0xD(52)(1) <= LUT_4bit_to_3bit(ChLLRxDI(127));
  CNStageIntLLRInputS0xD(57)(1) <= LUT_4bit_to_3bit(ChLLRxDI(127));
  CNStageIntLLRInputS0xD(117)(1) <= LUT_4bit_to_3bit(ChLLRxDI(127));
  CNStageIntLLRInputS0xD(173)(1) <= LUT_4bit_to_3bit(ChLLRxDI(127));
  CNStageIntLLRInputS0xD(277)(1) <= LUT_4bit_to_3bit(ChLLRxDI(127));
  CNStageIntLLRInputS0xD(306)(1) <= LUT_4bit_to_3bit(ChLLRxDI(127));
  CNStageIntLLRInputS0xD(373)(1) <= LUT_4bit_to_3bit(ChLLRxDI(127));
  CNStageIntLLRInputS0xD(53)(2) <= LUT_4bit_to_3bit(ChLLRxDI(128));
  CNStageIntLLRInputS0xD(108)(2) <= LUT_4bit_to_3bit(ChLLRxDI(128));
  CNStageIntLLRInputS0xD(129)(2) <= LUT_4bit_to_3bit(ChLLRxDI(128));
  CNStageIntLLRInputS0xD(198)(2) <= LUT_4bit_to_3bit(ChLLRxDI(128));
  CNStageIntLLRInputS0xD(244)(2) <= LUT_4bit_to_3bit(ChLLRxDI(128));
  CNStageIntLLRInputS0xD(298)(2) <= LUT_4bit_to_3bit(ChLLRxDI(128));
  CNStageIntLLRInputS0xD(341)(2) <= LUT_4bit_to_3bit(ChLLRxDI(128));
  CNStageIntLLRInputS0xD(51)(2) <= LUT_4bit_to_3bit(ChLLRxDI(129));
  CNStageIntLLRInputS0xD(56)(2) <= LUT_4bit_to_3bit(ChLLRxDI(129));
  CNStageIntLLRInputS0xD(116)(2) <= LUT_4bit_to_3bit(ChLLRxDI(129));
  CNStageIntLLRInputS0xD(172)(2) <= LUT_4bit_to_3bit(ChLLRxDI(129));
  CNStageIntLLRInputS0xD(276)(2) <= LUT_4bit_to_3bit(ChLLRxDI(129));
  CNStageIntLLRInputS0xD(305)(2) <= LUT_4bit_to_3bit(ChLLRxDI(129));
  CNStageIntLLRInputS0xD(372)(2) <= LUT_4bit_to_3bit(ChLLRxDI(129));
  CNStageIntLLRInputS0xD(50)(2) <= LUT_4bit_to_3bit(ChLLRxDI(130));
  CNStageIntLLRInputS0xD(73)(2) <= LUT_4bit_to_3bit(ChLLRxDI(130));
  CNStageIntLLRInputS0xD(140)(2) <= LUT_4bit_to_3bit(ChLLRxDI(130));
  CNStageIntLLRInputS0xD(188)(2) <= LUT_4bit_to_3bit(ChLLRxDI(130));
  CNStageIntLLRInputS0xD(245)(2) <= LUT_4bit_to_3bit(ChLLRxDI(130));
  CNStageIntLLRInputS0xD(285)(2) <= LUT_4bit_to_3bit(ChLLRxDI(130));
  CNStageIntLLRInputS0xD(65)(2) <= LUT_4bit_to_3bit(ChLLRxDI(131));
  CNStageIntLLRInputS0xD(154)(2) <= LUT_4bit_to_3bit(ChLLRxDI(131));
  CNStageIntLLRInputS0xD(206)(2) <= LUT_4bit_to_3bit(ChLLRxDI(131));
  CNStageIntLLRInputS0xD(243)(2) <= LUT_4bit_to_3bit(ChLLRxDI(131));
  CNStageIntLLRInputS0xD(307)(2) <= LUT_4bit_to_3bit(ChLLRxDI(131));
  CNStageIntLLRInputS0xD(334)(2) <= LUT_4bit_to_3bit(ChLLRxDI(131));
  CNStageIntLLRInputS0xD(49)(2) <= LUT_4bit_to_3bit(ChLLRxDI(132));
  CNStageIntLLRInputS0xD(151)(2) <= LUT_4bit_to_3bit(ChLLRxDI(132));
  CNStageIntLLRInputS0xD(214)(2) <= LUT_4bit_to_3bit(ChLLRxDI(132));
  CNStageIntLLRInputS0xD(274)(2) <= LUT_4bit_to_3bit(ChLLRxDI(132));
  CNStageIntLLRInputS0xD(321)(2) <= LUT_4bit_to_3bit(ChLLRxDI(132));
  CNStageIntLLRInputS0xD(364)(2) <= LUT_4bit_to_3bit(ChLLRxDI(132));
  CNStageIntLLRInputS0xD(48)(2) <= LUT_4bit_to_3bit(ChLLRxDI(133));
  CNStageIntLLRInputS0xD(209)(2) <= LUT_4bit_to_3bit(ChLLRxDI(133));
  CNStageIntLLRInputS0xD(255)(2) <= LUT_4bit_to_3bit(ChLLRxDI(133));
  CNStageIntLLRInputS0xD(317)(2) <= LUT_4bit_to_3bit(ChLLRxDI(133));
  CNStageIntLLRInputS0xD(380)(2) <= LUT_4bit_to_3bit(ChLLRxDI(133));
  CNStageIntLLRInputS0xD(47)(2) <= LUT_4bit_to_3bit(ChLLRxDI(134));
  CNStageIntLLRInputS0xD(100)(2) <= LUT_4bit_to_3bit(ChLLRxDI(134));
  CNStageIntLLRInputS0xD(134)(2) <= LUT_4bit_to_3bit(ChLLRxDI(134));
  CNStageIntLLRInputS0xD(258)(2) <= LUT_4bit_to_3bit(ChLLRxDI(134));
  CNStageIntLLRInputS0xD(46)(2) <= LUT_4bit_to_3bit(ChLLRxDI(135));
  CNStageIntLLRInputS0xD(103)(2) <= LUT_4bit_to_3bit(ChLLRxDI(135));
  CNStageIntLLRInputS0xD(135)(2) <= LUT_4bit_to_3bit(ChLLRxDI(135));
  CNStageIntLLRInputS0xD(205)(2) <= LUT_4bit_to_3bit(ChLLRxDI(135));
  CNStageIntLLRInputS0xD(45)(2) <= LUT_4bit_to_3bit(ChLLRxDI(136));
  CNStageIntLLRInputS0xD(94)(2) <= LUT_4bit_to_3bit(ChLLRxDI(136));
  CNStageIntLLRInputS0xD(111)(2) <= LUT_4bit_to_3bit(ChLLRxDI(136));
  CNStageIntLLRInputS0xD(175)(2) <= LUT_4bit_to_3bit(ChLLRxDI(136));
  CNStageIntLLRInputS0xD(275)(2) <= LUT_4bit_to_3bit(ChLLRxDI(136));
  CNStageIntLLRInputS0xD(301)(2) <= LUT_4bit_to_3bit(ChLLRxDI(136));
  CNStageIntLLRInputS0xD(352)(2) <= LUT_4bit_to_3bit(ChLLRxDI(136));
  CNStageIntLLRInputS0xD(44)(2) <= LUT_4bit_to_3bit(ChLLRxDI(137));
  CNStageIntLLRInputS0xD(74)(2) <= LUT_4bit_to_3bit(ChLLRxDI(137));
  CNStageIntLLRInputS0xD(161)(2) <= LUT_4bit_to_3bit(ChLLRxDI(137));
  CNStageIntLLRInputS0xD(182)(2) <= LUT_4bit_to_3bit(ChLLRxDI(137));
  CNStageIntLLRInputS0xD(242)(2) <= LUT_4bit_to_3bit(ChLLRxDI(137));
  CNStageIntLLRInputS0xD(282)(2) <= LUT_4bit_to_3bit(ChLLRxDI(137));
  CNStageIntLLRInputS0xD(366)(2) <= LUT_4bit_to_3bit(ChLLRxDI(137));
  CNStageIntLLRInputS0xD(43)(2) <= LUT_4bit_to_3bit(ChLLRxDI(138));
  CNStageIntLLRInputS0xD(55)(2) <= LUT_4bit_to_3bit(ChLLRxDI(138));
  CNStageIntLLRInputS0xD(120)(2) <= LUT_4bit_to_3bit(ChLLRxDI(138));
  CNStageIntLLRInputS0xD(218)(2) <= LUT_4bit_to_3bit(ChLLRxDI(138));
  CNStageIntLLRInputS0xD(268)(2) <= LUT_4bit_to_3bit(ChLLRxDI(138));
  CNStageIntLLRInputS0xD(327)(2) <= LUT_4bit_to_3bit(ChLLRxDI(138));
  CNStageIntLLRInputS0xD(362)(2) <= LUT_4bit_to_3bit(ChLLRxDI(138));
  CNStageIntLLRInputS0xD(42)(2) <= LUT_4bit_to_3bit(ChLLRxDI(139));
  CNStageIntLLRInputS0xD(69)(2) <= LUT_4bit_to_3bit(ChLLRxDI(139));
  CNStageIntLLRInputS0xD(124)(2) <= LUT_4bit_to_3bit(ChLLRxDI(139));
  CNStageIntLLRInputS0xD(220)(2) <= LUT_4bit_to_3bit(ChLLRxDI(139));
  CNStageIntLLRInputS0xD(252)(2) <= LUT_4bit_to_3bit(ChLLRxDI(139));
  CNStageIntLLRInputS0xD(289)(2) <= LUT_4bit_to_3bit(ChLLRxDI(139));
  CNStageIntLLRInputS0xD(383)(2) <= LUT_4bit_to_3bit(ChLLRxDI(139));
  CNStageIntLLRInputS0xD(41)(2) <= LUT_4bit_to_3bit(ChLLRxDI(140));
  CNStageIntLLRInputS0xD(80)(2) <= LUT_4bit_to_3bit(ChLLRxDI(140));
  CNStageIntLLRInputS0xD(170)(2) <= LUT_4bit_to_3bit(ChLLRxDI(140));
  CNStageIntLLRInputS0xD(191)(2) <= LUT_4bit_to_3bit(ChLLRxDI(140));
  CNStageIntLLRInputS0xD(277)(2) <= LUT_4bit_to_3bit(ChLLRxDI(140));
  CNStageIntLLRInputS0xD(293)(2) <= LUT_4bit_to_3bit(ChLLRxDI(140));
  CNStageIntLLRInputS0xD(346)(2) <= LUT_4bit_to_3bit(ChLLRxDI(140));
  CNStageIntLLRInputS0xD(123)(2) <= LUT_4bit_to_3bit(ChLLRxDI(141));
  CNStageIntLLRInputS0xD(173)(2) <= LUT_4bit_to_3bit(ChLLRxDI(141));
  CNStageIntLLRInputS0xD(269)(2) <= LUT_4bit_to_3bit(ChLLRxDI(141));
  CNStageIntLLRInputS0xD(332)(2) <= LUT_4bit_to_3bit(ChLLRxDI(141));
  CNStageIntLLRInputS0xD(347)(2) <= LUT_4bit_to_3bit(ChLLRxDI(141));
  CNStageIntLLRInputS0xD(40)(2) <= LUT_4bit_to_3bit(ChLLRxDI(142));
  CNStageIntLLRInputS0xD(96)(2) <= LUT_4bit_to_3bit(ChLLRxDI(142));
  CNStageIntLLRInputS0xD(118)(2) <= LUT_4bit_to_3bit(ChLLRxDI(142));
  CNStageIntLLRInputS0xD(256)(2) <= LUT_4bit_to_3bit(ChLLRxDI(142));
  CNStageIntLLRInputS0xD(382)(2) <= LUT_4bit_to_3bit(ChLLRxDI(142));
  CNStageIntLLRInputS0xD(39)(2) <= LUT_4bit_to_3bit(ChLLRxDI(143));
  CNStageIntLLRInputS0xD(83)(2) <= LUT_4bit_to_3bit(ChLLRxDI(143));
  CNStageIntLLRInputS0xD(158)(2) <= LUT_4bit_to_3bit(ChLLRxDI(143));
  CNStageIntLLRInputS0xD(192)(2) <= LUT_4bit_to_3bit(ChLLRxDI(143));
  CNStageIntLLRInputS0xD(273)(2) <= LUT_4bit_to_3bit(ChLLRxDI(143));
  CNStageIntLLRInputS0xD(287)(2) <= LUT_4bit_to_3bit(ChLLRxDI(143));
  CNStageIntLLRInputS0xD(373)(2) <= LUT_4bit_to_3bit(ChLLRxDI(143));
  CNStageIntLLRInputS0xD(38)(2) <= LUT_4bit_to_3bit(ChLLRxDI(144));
  CNStageIntLLRInputS0xD(98)(2) <= LUT_4bit_to_3bit(ChLLRxDI(144));
  CNStageIntLLRInputS0xD(166)(2) <= LUT_4bit_to_3bit(ChLLRxDI(144));
  CNStageIntLLRInputS0xD(219)(2) <= LUT_4bit_to_3bit(ChLLRxDI(144));
  CNStageIntLLRInputS0xD(249)(2) <= LUT_4bit_to_3bit(ChLLRxDI(144));
  CNStageIntLLRInputS0xD(324)(2) <= LUT_4bit_to_3bit(ChLLRxDI(144));
  CNStageIntLLRInputS0xD(333)(2) <= LUT_4bit_to_3bit(ChLLRxDI(144));
  CNStageIntLLRInputS0xD(37)(2) <= LUT_4bit_to_3bit(ChLLRxDI(145));
  CNStageIntLLRInputS0xD(61)(2) <= LUT_4bit_to_3bit(ChLLRxDI(145));
  CNStageIntLLRInputS0xD(130)(2) <= LUT_4bit_to_3bit(ChLLRxDI(145));
  CNStageIntLLRInputS0xD(181)(2) <= LUT_4bit_to_3bit(ChLLRxDI(145));
  CNStageIntLLRInputS0xD(247)(2) <= LUT_4bit_to_3bit(ChLLRxDI(145));
  CNStageIntLLRInputS0xD(331)(2) <= LUT_4bit_to_3bit(ChLLRxDI(145));
  CNStageIntLLRInputS0xD(336)(2) <= LUT_4bit_to_3bit(ChLLRxDI(145));
  CNStageIntLLRInputS0xD(36)(2) <= LUT_4bit_to_3bit(ChLLRxDI(146));
  CNStageIntLLRInputS0xD(71)(2) <= LUT_4bit_to_3bit(ChLLRxDI(146));
  CNStageIntLLRInputS0xD(128)(2) <= LUT_4bit_to_3bit(ChLLRxDI(146));
  CNStageIntLLRInputS0xD(261)(2) <= LUT_4bit_to_3bit(ChLLRxDI(146));
  CNStageIntLLRInputS0xD(299)(2) <= LUT_4bit_to_3bit(ChLLRxDI(146));
  CNStageIntLLRInputS0xD(35)(2) <= LUT_4bit_to_3bit(ChLLRxDI(147));
  CNStageIntLLRInputS0xD(66)(2) <= LUT_4bit_to_3bit(ChLLRxDI(147));
  CNStageIntLLRInputS0xD(164)(2) <= LUT_4bit_to_3bit(ChLLRxDI(147));
  CNStageIntLLRInputS0xD(187)(2) <= LUT_4bit_to_3bit(ChLLRxDI(147));
  CNStageIntLLRInputS0xD(253)(2) <= LUT_4bit_to_3bit(ChLLRxDI(147));
  CNStageIntLLRInputS0xD(297)(2) <= LUT_4bit_to_3bit(ChLLRxDI(147));
  CNStageIntLLRInputS0xD(335)(2) <= LUT_4bit_to_3bit(ChLLRxDI(147));
  CNStageIntLLRInputS0xD(34)(2) <= LUT_4bit_to_3bit(ChLLRxDI(148));
  CNStageIntLLRInputS0xD(72)(2) <= LUT_4bit_to_3bit(ChLLRxDI(148));
  CNStageIntLLRInputS0xD(143)(2) <= LUT_4bit_to_3bit(ChLLRxDI(148));
  CNStageIntLLRInputS0xD(207)(2) <= LUT_4bit_to_3bit(ChLLRxDI(148));
  CNStageIntLLRInputS0xD(231)(2) <= LUT_4bit_to_3bit(ChLLRxDI(148));
  CNStageIntLLRInputS0xD(329)(2) <= LUT_4bit_to_3bit(ChLLRxDI(148));
  CNStageIntLLRInputS0xD(33)(2) <= LUT_4bit_to_3bit(ChLLRxDI(149));
  CNStageIntLLRInputS0xD(60)(2) <= LUT_4bit_to_3bit(ChLLRxDI(149));
  CNStageIntLLRInputS0xD(146)(2) <= LUT_4bit_to_3bit(ChLLRxDI(149));
  CNStageIntLLRInputS0xD(221)(2) <= LUT_4bit_to_3bit(ChLLRxDI(149));
  CNStageIntLLRInputS0xD(241)(2) <= LUT_4bit_to_3bit(ChLLRxDI(149));
  CNStageIntLLRInputS0xD(309)(2) <= LUT_4bit_to_3bit(ChLLRxDI(149));
  CNStageIntLLRInputS0xD(370)(2) <= LUT_4bit_to_3bit(ChLLRxDI(149));
  CNStageIntLLRInputS0xD(32)(2) <= LUT_4bit_to_3bit(ChLLRxDI(150));
  CNStageIntLLRInputS0xD(86)(2) <= LUT_4bit_to_3bit(ChLLRxDI(150));
  CNStageIntLLRInputS0xD(131)(2) <= LUT_4bit_to_3bit(ChLLRxDI(150));
  CNStageIntLLRInputS0xD(217)(2) <= LUT_4bit_to_3bit(ChLLRxDI(150));
  CNStageIntLLRInputS0xD(312)(2) <= LUT_4bit_to_3bit(ChLLRxDI(150));
  CNStageIntLLRInputS0xD(378)(2) <= LUT_4bit_to_3bit(ChLLRxDI(150));
  CNStageIntLLRInputS0xD(31)(2) <= LUT_4bit_to_3bit(ChLLRxDI(151));
  CNStageIntLLRInputS0xD(92)(2) <= LUT_4bit_to_3bit(ChLLRxDI(151));
  CNStageIntLLRInputS0xD(165)(2) <= LUT_4bit_to_3bit(ChLLRxDI(151));
  CNStageIntLLRInputS0xD(184)(2) <= LUT_4bit_to_3bit(ChLLRxDI(151));
  CNStageIntLLRInputS0xD(238)(2) <= LUT_4bit_to_3bit(ChLLRxDI(151));
  CNStageIntLLRInputS0xD(342)(2) <= LUT_4bit_to_3bit(ChLLRxDI(151));
  CNStageIntLLRInputS0xD(30)(2) <= LUT_4bit_to_3bit(ChLLRxDI(152));
  CNStageIntLLRInputS0xD(76)(2) <= LUT_4bit_to_3bit(ChLLRxDI(152));
  CNStageIntLLRInputS0xD(127)(2) <= LUT_4bit_to_3bit(ChLLRxDI(152));
  CNStageIntLLRInputS0xD(202)(2) <= LUT_4bit_to_3bit(ChLLRxDI(152));
  CNStageIntLLRInputS0xD(228)(2) <= LUT_4bit_to_3bit(ChLLRxDI(152));
  CNStageIntLLRInputS0xD(330)(2) <= LUT_4bit_to_3bit(ChLLRxDI(152));
  CNStageIntLLRInputS0xD(340)(2) <= LUT_4bit_to_3bit(ChLLRxDI(152));
  CNStageIntLLRInputS0xD(29)(2) <= LUT_4bit_to_3bit(ChLLRxDI(153));
  CNStageIntLLRInputS0xD(78)(2) <= LUT_4bit_to_3bit(ChLLRxDI(153));
  CNStageIntLLRInputS0xD(155)(2) <= LUT_4bit_to_3bit(ChLLRxDI(153));
  CNStageIntLLRInputS0xD(203)(2) <= LUT_4bit_to_3bit(ChLLRxDI(153));
  CNStageIntLLRInputS0xD(262)(2) <= LUT_4bit_to_3bit(ChLLRxDI(153));
  CNStageIntLLRInputS0xD(296)(2) <= LUT_4bit_to_3bit(ChLLRxDI(153));
  CNStageIntLLRInputS0xD(376)(2) <= LUT_4bit_to_3bit(ChLLRxDI(153));
  CNStageIntLLRInputS0xD(28)(2) <= LUT_4bit_to_3bit(ChLLRxDI(154));
  CNStageIntLLRInputS0xD(139)(2) <= LUT_4bit_to_3bit(ChLLRxDI(154));
  CNStageIntLLRInputS0xD(183)(2) <= LUT_4bit_to_3bit(ChLLRxDI(154));
  CNStageIntLLRInputS0xD(246)(2) <= LUT_4bit_to_3bit(ChLLRxDI(154));
  CNStageIntLLRInputS0xD(322)(2) <= LUT_4bit_to_3bit(ChLLRxDI(154));
  CNStageIntLLRInputS0xD(27)(2) <= LUT_4bit_to_3bit(ChLLRxDI(155));
  CNStageIntLLRInputS0xD(84)(2) <= LUT_4bit_to_3bit(ChLLRxDI(155));
  CNStageIntLLRInputS0xD(167)(2) <= LUT_4bit_to_3bit(ChLLRxDI(155));
  CNStageIntLLRInputS0xD(174)(2) <= LUT_4bit_to_3bit(ChLLRxDI(155));
  CNStageIntLLRInputS0xD(257)(2) <= LUT_4bit_to_3bit(ChLLRxDI(155));
  CNStageIntLLRInputS0xD(306)(2) <= LUT_4bit_to_3bit(ChLLRxDI(155));
  CNStageIntLLRInputS0xD(357)(2) <= LUT_4bit_to_3bit(ChLLRxDI(155));
  CNStageIntLLRInputS0xD(26)(2) <= LUT_4bit_to_3bit(ChLLRxDI(156));
  CNStageIntLLRInputS0xD(95)(2) <= LUT_4bit_to_3bit(ChLLRxDI(156));
  CNStageIntLLRInputS0xD(157)(2) <= LUT_4bit_to_3bit(ChLLRxDI(156));
  CNStageIntLLRInputS0xD(343)(2) <= LUT_4bit_to_3bit(ChLLRxDI(156));
  CNStageIntLLRInputS0xD(25)(2) <= LUT_4bit_to_3bit(ChLLRxDI(157));
  CNStageIntLLRInputS0xD(102)(2) <= LUT_4bit_to_3bit(ChLLRxDI(157));
  CNStageIntLLRInputS0xD(144)(2) <= LUT_4bit_to_3bit(ChLLRxDI(157));
  CNStageIntLLRInputS0xD(194)(2) <= LUT_4bit_to_3bit(ChLLRxDI(157));
  CNStageIntLLRInputS0xD(323)(2) <= LUT_4bit_to_3bit(ChLLRxDI(157));
  CNStageIntLLRInputS0xD(377)(2) <= LUT_4bit_to_3bit(ChLLRxDI(157));
  CNStageIntLLRInputS0xD(24)(2) <= LUT_4bit_to_3bit(ChLLRxDI(158));
  CNStageIntLLRInputS0xD(77)(2) <= LUT_4bit_to_3bit(ChLLRxDI(158));
  CNStageIntLLRInputS0xD(163)(2) <= LUT_4bit_to_3bit(ChLLRxDI(158));
  CNStageIntLLRInputS0xD(224)(2) <= LUT_4bit_to_3bit(ChLLRxDI(158));
  CNStageIntLLRInputS0xD(230)(2) <= LUT_4bit_to_3bit(ChLLRxDI(158));
  CNStageIntLLRInputS0xD(310)(2) <= LUT_4bit_to_3bit(ChLLRxDI(158));
  CNStageIntLLRInputS0xD(339)(2) <= LUT_4bit_to_3bit(ChLLRxDI(158));
  CNStageIntLLRInputS0xD(23)(2) <= LUT_4bit_to_3bit(ChLLRxDI(159));
  CNStageIntLLRInputS0xD(91)(2) <= LUT_4bit_to_3bit(ChLLRxDI(159));
  CNStageIntLLRInputS0xD(136)(2) <= LUT_4bit_to_3bit(ChLLRxDI(159));
  CNStageIntLLRInputS0xD(271)(2) <= LUT_4bit_to_3bit(ChLLRxDI(159));
  CNStageIntLLRInputS0xD(367)(2) <= LUT_4bit_to_3bit(ChLLRxDI(159));
  CNStageIntLLRInputS0xD(22)(2) <= LUT_4bit_to_3bit(ChLLRxDI(160));
  CNStageIntLLRInputS0xD(62)(2) <= LUT_4bit_to_3bit(ChLLRxDI(160));
  CNStageIntLLRInputS0xD(133)(2) <= LUT_4bit_to_3bit(ChLLRxDI(160));
  CNStageIntLLRInputS0xD(189)(2) <= LUT_4bit_to_3bit(ChLLRxDI(160));
  CNStageIntLLRInputS0xD(233)(2) <= LUT_4bit_to_3bit(ChLLRxDI(160));
  CNStageIntLLRInputS0xD(302)(2) <= LUT_4bit_to_3bit(ChLLRxDI(160));
  CNStageIntLLRInputS0xD(351)(2) <= LUT_4bit_to_3bit(ChLLRxDI(160));
  CNStageIntLLRInputS0xD(21)(2) <= LUT_4bit_to_3bit(ChLLRxDI(161));
  CNStageIntLLRInputS0xD(97)(2) <= LUT_4bit_to_3bit(ChLLRxDI(161));
  CNStageIntLLRInputS0xD(149)(2) <= LUT_4bit_to_3bit(ChLLRxDI(161));
  CNStageIntLLRInputS0xD(171)(2) <= LUT_4bit_to_3bit(ChLLRxDI(161));
  CNStageIntLLRInputS0xD(250)(2) <= LUT_4bit_to_3bit(ChLLRxDI(161));
  CNStageIntLLRInputS0xD(300)(2) <= LUT_4bit_to_3bit(ChLLRxDI(161));
  CNStageIntLLRInputS0xD(379)(2) <= LUT_4bit_to_3bit(ChLLRxDI(161));
  CNStageIntLLRInputS0xD(20)(2) <= LUT_4bit_to_3bit(ChLLRxDI(162));
  CNStageIntLLRInputS0xD(64)(2) <= LUT_4bit_to_3bit(ChLLRxDI(162));
  CNStageIntLLRInputS0xD(141)(2) <= LUT_4bit_to_3bit(ChLLRxDI(162));
  CNStageIntLLRInputS0xD(179)(2) <= LUT_4bit_to_3bit(ChLLRxDI(162));
  CNStageIntLLRInputS0xD(259)(2) <= LUT_4bit_to_3bit(ChLLRxDI(162));
  CNStageIntLLRInputS0xD(315)(2) <= LUT_4bit_to_3bit(ChLLRxDI(162));
  CNStageIntLLRInputS0xD(369)(2) <= LUT_4bit_to_3bit(ChLLRxDI(162));
  CNStageIntLLRInputS0xD(19)(2) <= LUT_4bit_to_3bit(ChLLRxDI(163));
  CNStageIntLLRInputS0xD(79)(2) <= LUT_4bit_to_3bit(ChLLRxDI(163));
  CNStageIntLLRInputS0xD(115)(2) <= LUT_4bit_to_3bit(ChLLRxDI(163));
  CNStageIntLLRInputS0xD(254)(2) <= LUT_4bit_to_3bit(ChLLRxDI(163));
  CNStageIntLLRInputS0xD(355)(2) <= LUT_4bit_to_3bit(ChLLRxDI(163));
  CNStageIntLLRInputS0xD(18)(2) <= LUT_4bit_to_3bit(ChLLRxDI(164));
  CNStageIntLLRInputS0xD(75)(2) <= LUT_4bit_to_3bit(ChLLRxDI(164));
  CNStageIntLLRInputS0xD(125)(2) <= LUT_4bit_to_3bit(ChLLRxDI(164));
  CNStageIntLLRInputS0xD(197)(2) <= LUT_4bit_to_3bit(ChLLRxDI(164));
  CNStageIntLLRInputS0xD(260)(2) <= LUT_4bit_to_3bit(ChLLRxDI(164));
  CNStageIntLLRInputS0xD(375)(2) <= LUT_4bit_to_3bit(ChLLRxDI(164));
  CNStageIntLLRInputS0xD(17)(2) <= LUT_4bit_to_3bit(ChLLRxDI(165));
  CNStageIntLLRInputS0xD(93)(2) <= LUT_4bit_to_3bit(ChLLRxDI(165));
  CNStageIntLLRInputS0xD(119)(2) <= LUT_4bit_to_3bit(ChLLRxDI(165));
  CNStageIntLLRInputS0xD(177)(2) <= LUT_4bit_to_3bit(ChLLRxDI(165));
  CNStageIntLLRInputS0xD(294)(2) <= LUT_4bit_to_3bit(ChLLRxDI(165));
  CNStageIntLLRInputS0xD(348)(2) <= LUT_4bit_to_3bit(ChLLRxDI(165));
  CNStageIntLLRInputS0xD(16)(2) <= LUT_4bit_to_3bit(ChLLRxDI(166));
  CNStageIntLLRInputS0xD(57)(2) <= LUT_4bit_to_3bit(ChLLRxDI(166));
  CNStageIntLLRInputS0xD(122)(2) <= LUT_4bit_to_3bit(ChLLRxDI(166));
  CNStageIntLLRInputS0xD(210)(2) <= LUT_4bit_to_3bit(ChLLRxDI(166));
  CNStageIntLLRInputS0xD(288)(2) <= LUT_4bit_to_3bit(ChLLRxDI(166));
  CNStageIntLLRInputS0xD(345)(2) <= LUT_4bit_to_3bit(ChLLRxDI(166));
  CNStageIntLLRInputS0xD(15)(2) <= LUT_4bit_to_3bit(ChLLRxDI(167));
  CNStageIntLLRInputS0xD(58)(2) <= LUT_4bit_to_3bit(ChLLRxDI(167));
  CNStageIntLLRInputS0xD(112)(2) <= LUT_4bit_to_3bit(ChLLRxDI(167));
  CNStageIntLLRInputS0xD(213)(2) <= LUT_4bit_to_3bit(ChLLRxDI(167));
  CNStageIntLLRInputS0xD(225)(2) <= LUT_4bit_to_3bit(ChLLRxDI(167));
  CNStageIntLLRInputS0xD(292)(2) <= LUT_4bit_to_3bit(ChLLRxDI(167));
  CNStageIntLLRInputS0xD(360)(2) <= LUT_4bit_to_3bit(ChLLRxDI(167));
  CNStageIntLLRInputS0xD(14)(2) <= LUT_4bit_to_3bit(ChLLRxDI(168));
  CNStageIntLLRInputS0xD(150)(2) <= LUT_4bit_to_3bit(ChLLRxDI(168));
  CNStageIntLLRInputS0xD(199)(2) <= LUT_4bit_to_3bit(ChLLRxDI(168));
  CNStageIntLLRInputS0xD(264)(2) <= LUT_4bit_to_3bit(ChLLRxDI(168));
  CNStageIntLLRInputS0xD(283)(2) <= LUT_4bit_to_3bit(ChLLRxDI(168));
  CNStageIntLLRInputS0xD(353)(2) <= LUT_4bit_to_3bit(ChLLRxDI(168));
  CNStageIntLLRInputS0xD(13)(2) <= LUT_4bit_to_3bit(ChLLRxDI(169));
  CNStageIntLLRInputS0xD(85)(2) <= LUT_4bit_to_3bit(ChLLRxDI(169));
  CNStageIntLLRInputS0xD(132)(2) <= LUT_4bit_to_3bit(ChLLRxDI(169));
  CNStageIntLLRInputS0xD(178)(2) <= LUT_4bit_to_3bit(ChLLRxDI(169));
  CNStageIntLLRInputS0xD(266)(2) <= LUT_4bit_to_3bit(ChLLRxDI(169));
  CNStageIntLLRInputS0xD(316)(2) <= LUT_4bit_to_3bit(ChLLRxDI(169));
  CNStageIntLLRInputS0xD(12)(2) <= LUT_4bit_to_3bit(ChLLRxDI(170));
  CNStageIntLLRInputS0xD(101)(2) <= LUT_4bit_to_3bit(ChLLRxDI(170));
  CNStageIntLLRInputS0xD(145)(2) <= LUT_4bit_to_3bit(ChLLRxDI(170));
  CNStageIntLLRInputS0xD(236)(2) <= LUT_4bit_to_3bit(ChLLRxDI(170));
  CNStageIntLLRInputS0xD(337)(2) <= LUT_4bit_to_3bit(ChLLRxDI(170));
  CNStageIntLLRInputS0xD(105)(2) <= LUT_4bit_to_3bit(ChLLRxDI(171));
  CNStageIntLLRInputS0xD(156)(2) <= LUT_4bit_to_3bit(ChLLRxDI(171));
  CNStageIntLLRInputS0xD(222)(2) <= LUT_4bit_to_3bit(ChLLRxDI(171));
  CNStageIntLLRInputS0xD(311)(2) <= LUT_4bit_to_3bit(ChLLRxDI(171));
  CNStageIntLLRInputS0xD(11)(2) <= LUT_4bit_to_3bit(ChLLRxDI(172));
  CNStageIntLLRInputS0xD(110)(2) <= LUT_4bit_to_3bit(ChLLRxDI(172));
  CNStageIntLLRInputS0xD(126)(2) <= LUT_4bit_to_3bit(ChLLRxDI(172));
  CNStageIntLLRInputS0xD(229)(2) <= LUT_4bit_to_3bit(ChLLRxDI(172));
  CNStageIntLLRInputS0xD(10)(2) <= LUT_4bit_to_3bit(ChLLRxDI(173));
  CNStageIntLLRInputS0xD(104)(2) <= LUT_4bit_to_3bit(ChLLRxDI(173));
  CNStageIntLLRInputS0xD(114)(2) <= LUT_4bit_to_3bit(ChLLRxDI(173));
  CNStageIntLLRInputS0xD(180)(2) <= LUT_4bit_to_3bit(ChLLRxDI(173));
  CNStageIntLLRInputS0xD(237)(2) <= LUT_4bit_to_3bit(ChLLRxDI(173));
  CNStageIntLLRInputS0xD(295)(2) <= LUT_4bit_to_3bit(ChLLRxDI(173));
  CNStageIntLLRInputS0xD(9)(2) <= LUT_4bit_to_3bit(ChLLRxDI(174));
  CNStageIntLLRInputS0xD(99)(2) <= LUT_4bit_to_3bit(ChLLRxDI(174));
  CNStageIntLLRInputS0xD(159)(2) <= LUT_4bit_to_3bit(ChLLRxDI(174));
  CNStageIntLLRInputS0xD(265)(2) <= LUT_4bit_to_3bit(ChLLRxDI(174));
  CNStageIntLLRInputS0xD(361)(2) <= LUT_4bit_to_3bit(ChLLRxDI(174));
  CNStageIntLLRInputS0xD(8)(2) <= LUT_4bit_to_3bit(ChLLRxDI(175));
  CNStageIntLLRInputS0xD(82)(2) <= LUT_4bit_to_3bit(ChLLRxDI(175));
  CNStageIntLLRInputS0xD(117)(2) <= LUT_4bit_to_3bit(ChLLRxDI(175));
  CNStageIntLLRInputS0xD(211)(2) <= LUT_4bit_to_3bit(ChLLRxDI(175));
  CNStageIntLLRInputS0xD(278)(2) <= LUT_4bit_to_3bit(ChLLRxDI(175));
  CNStageIntLLRInputS0xD(325)(2) <= LUT_4bit_to_3bit(ChLLRxDI(175));
  CNStageIntLLRInputS0xD(344)(2) <= LUT_4bit_to_3bit(ChLLRxDI(175));
  CNStageIntLLRInputS0xD(7)(2) <= LUT_4bit_to_3bit(ChLLRxDI(176));
  CNStageIntLLRInputS0xD(89)(2) <= LUT_4bit_to_3bit(ChLLRxDI(176));
  CNStageIntLLRInputS0xD(137)(2) <= LUT_4bit_to_3bit(ChLLRxDI(176));
  CNStageIntLLRInputS0xD(176)(2) <= LUT_4bit_to_3bit(ChLLRxDI(176));
  CNStageIntLLRInputS0xD(251)(2) <= LUT_4bit_to_3bit(ChLLRxDI(176));
  CNStageIntLLRInputS0xD(286)(2) <= LUT_4bit_to_3bit(ChLLRxDI(176));
  CNStageIntLLRInputS0xD(356)(2) <= LUT_4bit_to_3bit(ChLLRxDI(176));
  CNStageIntLLRInputS0xD(6)(2) <= LUT_4bit_to_3bit(ChLLRxDI(177));
  CNStageIntLLRInputS0xD(109)(2) <= LUT_4bit_to_3bit(ChLLRxDI(177));
  CNStageIntLLRInputS0xD(147)(2) <= LUT_4bit_to_3bit(ChLLRxDI(177));
  CNStageIntLLRInputS0xD(204)(2) <= LUT_4bit_to_3bit(ChLLRxDI(177));
  CNStageIntLLRInputS0xD(232)(2) <= LUT_4bit_to_3bit(ChLLRxDI(177));
  CNStageIntLLRInputS0xD(304)(2) <= LUT_4bit_to_3bit(ChLLRxDI(177));
  CNStageIntLLRInputS0xD(368)(2) <= LUT_4bit_to_3bit(ChLLRxDI(177));
  CNStageIntLLRInputS0xD(5)(2) <= LUT_4bit_to_3bit(ChLLRxDI(178));
  CNStageIntLLRInputS0xD(107)(2) <= LUT_4bit_to_3bit(ChLLRxDI(178));
  CNStageIntLLRInputS0xD(142)(2) <= LUT_4bit_to_3bit(ChLLRxDI(178));
  CNStageIntLLRInputS0xD(201)(2) <= LUT_4bit_to_3bit(ChLLRxDI(178));
  CNStageIntLLRInputS0xD(313)(2) <= LUT_4bit_to_3bit(ChLLRxDI(178));
  CNStageIntLLRInputS0xD(338)(2) <= LUT_4bit_to_3bit(ChLLRxDI(178));
  CNStageIntLLRInputS0xD(4)(2) <= LUT_4bit_to_3bit(ChLLRxDI(179));
  CNStageIntLLRInputS0xD(87)(2) <= LUT_4bit_to_3bit(ChLLRxDI(179));
  CNStageIntLLRInputS0xD(148)(2) <= LUT_4bit_to_3bit(ChLLRxDI(179));
  CNStageIntLLRInputS0xD(215)(2) <= LUT_4bit_to_3bit(ChLLRxDI(179));
  CNStageIntLLRInputS0xD(267)(2) <= LUT_4bit_to_3bit(ChLLRxDI(179));
  CNStageIntLLRInputS0xD(308)(2) <= LUT_4bit_to_3bit(ChLLRxDI(179));
  CNStageIntLLRInputS0xD(67)(2) <= LUT_4bit_to_3bit(ChLLRxDI(180));
  CNStageIntLLRInputS0xD(208)(2) <= LUT_4bit_to_3bit(ChLLRxDI(180));
  CNStageIntLLRInputS0xD(263)(2) <= LUT_4bit_to_3bit(ChLLRxDI(180));
  CNStageIntLLRInputS0xD(314)(2) <= LUT_4bit_to_3bit(ChLLRxDI(180));
  CNStageIntLLRInputS0xD(371)(2) <= LUT_4bit_to_3bit(ChLLRxDI(180));
  CNStageIntLLRInputS0xD(3)(2) <= LUT_4bit_to_3bit(ChLLRxDI(181));
  CNStageIntLLRInputS0xD(70)(2) <= LUT_4bit_to_3bit(ChLLRxDI(181));
  CNStageIntLLRInputS0xD(162)(2) <= LUT_4bit_to_3bit(ChLLRxDI(181));
  CNStageIntLLRInputS0xD(186)(2) <= LUT_4bit_to_3bit(ChLLRxDI(181));
  CNStageIntLLRInputS0xD(227)(2) <= LUT_4bit_to_3bit(ChLLRxDI(181));
  CNStageIntLLRInputS0xD(303)(2) <= LUT_4bit_to_3bit(ChLLRxDI(181));
  CNStageIntLLRInputS0xD(2)(2) <= LUT_4bit_to_3bit(ChLLRxDI(182));
  CNStageIntLLRInputS0xD(54)(2) <= LUT_4bit_to_3bit(ChLLRxDI(182));
  CNStageIntLLRInputS0xD(169)(2) <= LUT_4bit_to_3bit(ChLLRxDI(182));
  CNStageIntLLRInputS0xD(195)(2) <= LUT_4bit_to_3bit(ChLLRxDI(182));
  CNStageIntLLRInputS0xD(248)(2) <= LUT_4bit_to_3bit(ChLLRxDI(182));
  CNStageIntLLRInputS0xD(328)(2) <= LUT_4bit_to_3bit(ChLLRxDI(182));
  CNStageIntLLRInputS0xD(350)(2) <= LUT_4bit_to_3bit(ChLLRxDI(182));
  CNStageIntLLRInputS0xD(1)(2) <= LUT_4bit_to_3bit(ChLLRxDI(183));
  CNStageIntLLRInputS0xD(88)(2) <= LUT_4bit_to_3bit(ChLLRxDI(183));
  CNStageIntLLRInputS0xD(190)(2) <= LUT_4bit_to_3bit(ChLLRxDI(183));
  CNStageIntLLRInputS0xD(281)(2) <= LUT_4bit_to_3bit(ChLLRxDI(183));
  CNStageIntLLRInputS0xD(358)(2) <= LUT_4bit_to_3bit(ChLLRxDI(183));
  CNStageIntLLRInputS0xD(0)(2) <= LUT_4bit_to_3bit(ChLLRxDI(184));
  CNStageIntLLRInputS0xD(106)(2) <= LUT_4bit_to_3bit(ChLLRxDI(184));
  CNStageIntLLRInputS0xD(153)(2) <= LUT_4bit_to_3bit(ChLLRxDI(184));
  CNStageIntLLRInputS0xD(193)(2) <= LUT_4bit_to_3bit(ChLLRxDI(184));
  CNStageIntLLRInputS0xD(226)(2) <= LUT_4bit_to_3bit(ChLLRxDI(184));
  CNStageIntLLRInputS0xD(318)(2) <= LUT_4bit_to_3bit(ChLLRxDI(184));
  CNStageIntLLRInputS0xD(354)(2) <= LUT_4bit_to_3bit(ChLLRxDI(184));
  CNStageIntLLRInputS0xD(121)(2) <= LUT_4bit_to_3bit(ChLLRxDI(185));
  CNStageIntLLRInputS0xD(272)(2) <= LUT_4bit_to_3bit(ChLLRxDI(185));
  CNStageIntLLRInputS0xD(320)(2) <= LUT_4bit_to_3bit(ChLLRxDI(185));
  CNStageIntLLRInputS0xD(359)(2) <= LUT_4bit_to_3bit(ChLLRxDI(185));
  CNStageIntLLRInputS0xD(63)(2) <= LUT_4bit_to_3bit(ChLLRxDI(186));
  CNStageIntLLRInputS0xD(160)(2) <= LUT_4bit_to_3bit(ChLLRxDI(186));
  CNStageIntLLRInputS0xD(216)(2) <= LUT_4bit_to_3bit(ChLLRxDI(186));
  CNStageIntLLRInputS0xD(235)(2) <= LUT_4bit_to_3bit(ChLLRxDI(186));
  CNStageIntLLRInputS0xD(290)(2) <= LUT_4bit_to_3bit(ChLLRxDI(186));
  CNStageIntLLRInputS0xD(349)(2) <= LUT_4bit_to_3bit(ChLLRxDI(186));
  CNStageIntLLRInputS0xD(90)(2) <= LUT_4bit_to_3bit(ChLLRxDI(187));
  CNStageIntLLRInputS0xD(113)(2) <= LUT_4bit_to_3bit(ChLLRxDI(187));
  CNStageIntLLRInputS0xD(200)(2) <= LUT_4bit_to_3bit(ChLLRxDI(187));
  CNStageIntLLRInputS0xD(240)(2) <= LUT_4bit_to_3bit(ChLLRxDI(187));
  CNStageIntLLRInputS0xD(326)(2) <= LUT_4bit_to_3bit(ChLLRxDI(187));
  CNStageIntLLRInputS0xD(374)(2) <= LUT_4bit_to_3bit(ChLLRxDI(187));
  CNStageIntLLRInputS0xD(81)(2) <= LUT_4bit_to_3bit(ChLLRxDI(188));
  CNStageIntLLRInputS0xD(212)(2) <= LUT_4bit_to_3bit(ChLLRxDI(188));
  CNStageIntLLRInputS0xD(279)(2) <= LUT_4bit_to_3bit(ChLLRxDI(188));
  CNStageIntLLRInputS0xD(284)(2) <= LUT_4bit_to_3bit(ChLLRxDI(188));
  CNStageIntLLRInputS0xD(381)(2) <= LUT_4bit_to_3bit(ChLLRxDI(188));
  CNStageIntLLRInputS0xD(68)(2) <= LUT_4bit_to_3bit(ChLLRxDI(189));
  CNStageIntLLRInputS0xD(152)(2) <= LUT_4bit_to_3bit(ChLLRxDI(189));
  CNStageIntLLRInputS0xD(223)(2) <= LUT_4bit_to_3bit(ChLLRxDI(189));
  CNStageIntLLRInputS0xD(239)(2) <= LUT_4bit_to_3bit(ChLLRxDI(189));
  CNStageIntLLRInputS0xD(291)(2) <= LUT_4bit_to_3bit(ChLLRxDI(189));
  CNStageIntLLRInputS0xD(363)(2) <= LUT_4bit_to_3bit(ChLLRxDI(189));
  CNStageIntLLRInputS0xD(168)(2) <= LUT_4bit_to_3bit(ChLLRxDI(190));
  CNStageIntLLRInputS0xD(196)(2) <= LUT_4bit_to_3bit(ChLLRxDI(190));
  CNStageIntLLRInputS0xD(234)(2) <= LUT_4bit_to_3bit(ChLLRxDI(190));
  CNStageIntLLRInputS0xD(319)(2) <= LUT_4bit_to_3bit(ChLLRxDI(190));
  CNStageIntLLRInputS0xD(365)(2) <= LUT_4bit_to_3bit(ChLLRxDI(190));
  CNStageIntLLRInputS0xD(52)(2) <= LUT_4bit_to_3bit(ChLLRxDI(191));
  CNStageIntLLRInputS0xD(59)(2) <= LUT_4bit_to_3bit(ChLLRxDI(191));
  CNStageIntLLRInputS0xD(138)(2) <= LUT_4bit_to_3bit(ChLLRxDI(191));
  CNStageIntLLRInputS0xD(185)(2) <= LUT_4bit_to_3bit(ChLLRxDI(191));
  CNStageIntLLRInputS0xD(270)(2) <= LUT_4bit_to_3bit(ChLLRxDI(191));
  CNStageIntLLRInputS0xD(280)(2) <= LUT_4bit_to_3bit(ChLLRxDI(191));
  CNStageIntLLRInputS0xD(53)(3) <= LUT_4bit_to_3bit(ChLLRxDI(192));
  CNStageIntLLRInputS0xD(107)(3) <= LUT_4bit_to_3bit(ChLLRxDI(192));
  CNStageIntLLRInputS0xD(128)(3) <= LUT_4bit_to_3bit(ChLLRxDI(192));
  CNStageIntLLRInputS0xD(197)(3) <= LUT_4bit_to_3bit(ChLLRxDI(192));
  CNStageIntLLRInputS0xD(243)(3) <= LUT_4bit_to_3bit(ChLLRxDI(192));
  CNStageIntLLRInputS0xD(297)(3) <= LUT_4bit_to_3bit(ChLLRxDI(192));
  CNStageIntLLRInputS0xD(340)(3) <= LUT_4bit_to_3bit(ChLLRxDI(192));
  CNStageIntLLRInputS0xD(51)(3) <= LUT_4bit_to_3bit(ChLLRxDI(193));
  CNStageIntLLRInputS0xD(58)(3) <= LUT_4bit_to_3bit(ChLLRxDI(193));
  CNStageIntLLRInputS0xD(137)(3) <= LUT_4bit_to_3bit(ChLLRxDI(193));
  CNStageIntLLRInputS0xD(269)(3) <= LUT_4bit_to_3bit(ChLLRxDI(193));
  CNStageIntLLRInputS0xD(333)(3) <= LUT_4bit_to_3bit(ChLLRxDI(193));
  CNStageIntLLRInputS0xD(50)(3) <= LUT_4bit_to_3bit(ChLLRxDI(194));
  CNStageIntLLRInputS0xD(55)(3) <= LUT_4bit_to_3bit(ChLLRxDI(194));
  CNStageIntLLRInputS0xD(115)(3) <= LUT_4bit_to_3bit(ChLLRxDI(194));
  CNStageIntLLRInputS0xD(171)(3) <= LUT_4bit_to_3bit(ChLLRxDI(194));
  CNStageIntLLRInputS0xD(275)(3) <= LUT_4bit_to_3bit(ChLLRxDI(194));
  CNStageIntLLRInputS0xD(304)(3) <= LUT_4bit_to_3bit(ChLLRxDI(194));
  CNStageIntLLRInputS0xD(371)(3) <= LUT_4bit_to_3bit(ChLLRxDI(194));
  CNStageIntLLRInputS0xD(72)(3) <= LUT_4bit_to_3bit(ChLLRxDI(195));
  CNStageIntLLRInputS0xD(139)(3) <= LUT_4bit_to_3bit(ChLLRxDI(195));
  CNStageIntLLRInputS0xD(187)(3) <= LUT_4bit_to_3bit(ChLLRxDI(195));
  CNStageIntLLRInputS0xD(244)(3) <= LUT_4bit_to_3bit(ChLLRxDI(195));
  CNStageIntLLRInputS0xD(49)(3) <= LUT_4bit_to_3bit(ChLLRxDI(196));
  CNStageIntLLRInputS0xD(64)(3) <= LUT_4bit_to_3bit(ChLLRxDI(196));
  CNStageIntLLRInputS0xD(153)(3) <= LUT_4bit_to_3bit(ChLLRxDI(196));
  CNStageIntLLRInputS0xD(205)(3) <= LUT_4bit_to_3bit(ChLLRxDI(196));
  CNStageIntLLRInputS0xD(242)(3) <= LUT_4bit_to_3bit(ChLLRxDI(196));
  CNStageIntLLRInputS0xD(306)(3) <= LUT_4bit_to_3bit(ChLLRxDI(196));
  CNStageIntLLRInputS0xD(48)(3) <= LUT_4bit_to_3bit(ChLLRxDI(197));
  CNStageIntLLRInputS0xD(96)(3) <= LUT_4bit_to_3bit(ChLLRxDI(197));
  CNStageIntLLRInputS0xD(150)(3) <= LUT_4bit_to_3bit(ChLLRxDI(197));
  CNStageIntLLRInputS0xD(213)(3) <= LUT_4bit_to_3bit(ChLLRxDI(197));
  CNStageIntLLRInputS0xD(273)(3) <= LUT_4bit_to_3bit(ChLLRxDI(197));
  CNStageIntLLRInputS0xD(320)(3) <= LUT_4bit_to_3bit(ChLLRxDI(197));
  CNStageIntLLRInputS0xD(363)(3) <= LUT_4bit_to_3bit(ChLLRxDI(197));
  CNStageIntLLRInputS0xD(47)(3) <= LUT_4bit_to_3bit(ChLLRxDI(198));
  CNStageIntLLRInputS0xD(105)(3) <= LUT_4bit_to_3bit(ChLLRxDI(198));
  CNStageIntLLRInputS0xD(111)(3) <= LUT_4bit_to_3bit(ChLLRxDI(198));
  CNStageIntLLRInputS0xD(208)(3) <= LUT_4bit_to_3bit(ChLLRxDI(198));
  CNStageIntLLRInputS0xD(254)(3) <= LUT_4bit_to_3bit(ChLLRxDI(198));
  CNStageIntLLRInputS0xD(316)(3) <= LUT_4bit_to_3bit(ChLLRxDI(198));
  CNStageIntLLRInputS0xD(379)(3) <= LUT_4bit_to_3bit(ChLLRxDI(198));
  CNStageIntLLRInputS0xD(46)(3) <= LUT_4bit_to_3bit(ChLLRxDI(199));
  CNStageIntLLRInputS0xD(99)(3) <= LUT_4bit_to_3bit(ChLLRxDI(199));
  CNStageIntLLRInputS0xD(133)(3) <= LUT_4bit_to_3bit(ChLLRxDI(199));
  CNStageIntLLRInputS0xD(214)(3) <= LUT_4bit_to_3bit(ChLLRxDI(199));
  CNStageIntLLRInputS0xD(257)(3) <= LUT_4bit_to_3bit(ChLLRxDI(199));
  CNStageIntLLRInputS0xD(282)(3) <= LUT_4bit_to_3bit(ChLLRxDI(199));
  CNStageIntLLRInputS0xD(350)(3) <= LUT_4bit_to_3bit(ChLLRxDI(199));
  CNStageIntLLRInputS0xD(45)(3) <= LUT_4bit_to_3bit(ChLLRxDI(200));
  CNStageIntLLRInputS0xD(102)(3) <= LUT_4bit_to_3bit(ChLLRxDI(200));
  CNStageIntLLRInputS0xD(134)(3) <= LUT_4bit_to_3bit(ChLLRxDI(200));
  CNStageIntLLRInputS0xD(204)(3) <= LUT_4bit_to_3bit(ChLLRxDI(200));
  CNStageIntLLRInputS0xD(245)(3) <= LUT_4bit_to_3bit(ChLLRxDI(200));
  CNStageIntLLRInputS0xD(300)(3) <= LUT_4bit_to_3bit(ChLLRxDI(200));
  CNStageIntLLRInputS0xD(44)(3) <= LUT_4bit_to_3bit(ChLLRxDI(201));
  CNStageIntLLRInputS0xD(93)(3) <= LUT_4bit_to_3bit(ChLLRxDI(201));
  CNStageIntLLRInputS0xD(169)(3) <= LUT_4bit_to_3bit(ChLLRxDI(201));
  CNStageIntLLRInputS0xD(174)(3) <= LUT_4bit_to_3bit(ChLLRxDI(201));
  CNStageIntLLRInputS0xD(274)(3) <= LUT_4bit_to_3bit(ChLLRxDI(201));
  CNStageIntLLRInputS0xD(351)(3) <= LUT_4bit_to_3bit(ChLLRxDI(201));
  CNStageIntLLRInputS0xD(43)(3) <= LUT_4bit_to_3bit(ChLLRxDI(202));
  CNStageIntLLRInputS0xD(73)(3) <= LUT_4bit_to_3bit(ChLLRxDI(202));
  CNStageIntLLRInputS0xD(160)(3) <= LUT_4bit_to_3bit(ChLLRxDI(202));
  CNStageIntLLRInputS0xD(181)(3) <= LUT_4bit_to_3bit(ChLLRxDI(202));
  CNStageIntLLRInputS0xD(281)(3) <= LUT_4bit_to_3bit(ChLLRxDI(202));
  CNStageIntLLRInputS0xD(365)(3) <= LUT_4bit_to_3bit(ChLLRxDI(202));
  CNStageIntLLRInputS0xD(42)(3) <= LUT_4bit_to_3bit(ChLLRxDI(203));
  CNStageIntLLRInputS0xD(54)(3) <= LUT_4bit_to_3bit(ChLLRxDI(203));
  CNStageIntLLRInputS0xD(119)(3) <= LUT_4bit_to_3bit(ChLLRxDI(203));
  CNStageIntLLRInputS0xD(217)(3) <= LUT_4bit_to_3bit(ChLLRxDI(203));
  CNStageIntLLRInputS0xD(267)(3) <= LUT_4bit_to_3bit(ChLLRxDI(203));
  CNStageIntLLRInputS0xD(326)(3) <= LUT_4bit_to_3bit(ChLLRxDI(203));
  CNStageIntLLRInputS0xD(361)(3) <= LUT_4bit_to_3bit(ChLLRxDI(203));
  CNStageIntLLRInputS0xD(41)(3) <= LUT_4bit_to_3bit(ChLLRxDI(204));
  CNStageIntLLRInputS0xD(68)(3) <= LUT_4bit_to_3bit(ChLLRxDI(204));
  CNStageIntLLRInputS0xD(123)(3) <= LUT_4bit_to_3bit(ChLLRxDI(204));
  CNStageIntLLRInputS0xD(219)(3) <= LUT_4bit_to_3bit(ChLLRxDI(204));
  CNStageIntLLRInputS0xD(251)(3) <= LUT_4bit_to_3bit(ChLLRxDI(204));
  CNStageIntLLRInputS0xD(288)(3) <= LUT_4bit_to_3bit(ChLLRxDI(204));
  CNStageIntLLRInputS0xD(382)(3) <= LUT_4bit_to_3bit(ChLLRxDI(204));
  CNStageIntLLRInputS0xD(170)(3) <= LUT_4bit_to_3bit(ChLLRxDI(205));
  CNStageIntLLRInputS0xD(276)(3) <= LUT_4bit_to_3bit(ChLLRxDI(205));
  CNStageIntLLRInputS0xD(345)(3) <= LUT_4bit_to_3bit(ChLLRxDI(205));
  CNStageIntLLRInputS0xD(40)(3) <= LUT_4bit_to_3bit(ChLLRxDI(206));
  CNStageIntLLRInputS0xD(122)(3) <= LUT_4bit_to_3bit(ChLLRxDI(206));
  CNStageIntLLRInputS0xD(172)(3) <= LUT_4bit_to_3bit(ChLLRxDI(206));
  CNStageIntLLRInputS0xD(332)(3) <= LUT_4bit_to_3bit(ChLLRxDI(206));
  CNStageIntLLRInputS0xD(346)(3) <= LUT_4bit_to_3bit(ChLLRxDI(206));
  CNStageIntLLRInputS0xD(39)(3) <= LUT_4bit_to_3bit(ChLLRxDI(207));
  CNStageIntLLRInputS0xD(95)(3) <= LUT_4bit_to_3bit(ChLLRxDI(207));
  CNStageIntLLRInputS0xD(117)(3) <= LUT_4bit_to_3bit(ChLLRxDI(207));
  CNStageIntLLRInputS0xD(255)(3) <= LUT_4bit_to_3bit(ChLLRxDI(207));
  CNStageIntLLRInputS0xD(292)(3) <= LUT_4bit_to_3bit(ChLLRxDI(207));
  CNStageIntLLRInputS0xD(381)(3) <= LUT_4bit_to_3bit(ChLLRxDI(207));
  CNStageIntLLRInputS0xD(38)(3) <= LUT_4bit_to_3bit(ChLLRxDI(208));
  CNStageIntLLRInputS0xD(82)(3) <= LUT_4bit_to_3bit(ChLLRxDI(208));
  CNStageIntLLRInputS0xD(157)(3) <= LUT_4bit_to_3bit(ChLLRxDI(208));
  CNStageIntLLRInputS0xD(191)(3) <= LUT_4bit_to_3bit(ChLLRxDI(208));
  CNStageIntLLRInputS0xD(286)(3) <= LUT_4bit_to_3bit(ChLLRxDI(208));
  CNStageIntLLRInputS0xD(372)(3) <= LUT_4bit_to_3bit(ChLLRxDI(208));
  CNStageIntLLRInputS0xD(37)(3) <= LUT_4bit_to_3bit(ChLLRxDI(209));
  CNStageIntLLRInputS0xD(97)(3) <= LUT_4bit_to_3bit(ChLLRxDI(209));
  CNStageIntLLRInputS0xD(165)(3) <= LUT_4bit_to_3bit(ChLLRxDI(209));
  CNStageIntLLRInputS0xD(218)(3) <= LUT_4bit_to_3bit(ChLLRxDI(209));
  CNStageIntLLRInputS0xD(323)(3) <= LUT_4bit_to_3bit(ChLLRxDI(209));
  CNStageIntLLRInputS0xD(36)(3) <= LUT_4bit_to_3bit(ChLLRxDI(210));
  CNStageIntLLRInputS0xD(60)(3) <= LUT_4bit_to_3bit(ChLLRxDI(210));
  CNStageIntLLRInputS0xD(129)(3) <= LUT_4bit_to_3bit(ChLLRxDI(210));
  CNStageIntLLRInputS0xD(180)(3) <= LUT_4bit_to_3bit(ChLLRxDI(210));
  CNStageIntLLRInputS0xD(246)(3) <= LUT_4bit_to_3bit(ChLLRxDI(210));
  CNStageIntLLRInputS0xD(330)(3) <= LUT_4bit_to_3bit(ChLLRxDI(210));
  CNStageIntLLRInputS0xD(335)(3) <= LUT_4bit_to_3bit(ChLLRxDI(210));
  CNStageIntLLRInputS0xD(35)(3) <= LUT_4bit_to_3bit(ChLLRxDI(211));
  CNStageIntLLRInputS0xD(70)(3) <= LUT_4bit_to_3bit(ChLLRxDI(211));
  CNStageIntLLRInputS0xD(127)(3) <= LUT_4bit_to_3bit(ChLLRxDI(211));
  CNStageIntLLRInputS0xD(206)(3) <= LUT_4bit_to_3bit(ChLLRxDI(211));
  CNStageIntLLRInputS0xD(260)(3) <= LUT_4bit_to_3bit(ChLLRxDI(211));
  CNStageIntLLRInputS0xD(298)(3) <= LUT_4bit_to_3bit(ChLLRxDI(211));
  CNStageIntLLRInputS0xD(34)(3) <= LUT_4bit_to_3bit(ChLLRxDI(212));
  CNStageIntLLRInputS0xD(65)(3) <= LUT_4bit_to_3bit(ChLLRxDI(212));
  CNStageIntLLRInputS0xD(163)(3) <= LUT_4bit_to_3bit(ChLLRxDI(212));
  CNStageIntLLRInputS0xD(186)(3) <= LUT_4bit_to_3bit(ChLLRxDI(212));
  CNStageIntLLRInputS0xD(296)(3) <= LUT_4bit_to_3bit(ChLLRxDI(212));
  CNStageIntLLRInputS0xD(33)(3) <= LUT_4bit_to_3bit(ChLLRxDI(213));
  CNStageIntLLRInputS0xD(71)(3) <= LUT_4bit_to_3bit(ChLLRxDI(213));
  CNStageIntLLRInputS0xD(142)(3) <= LUT_4bit_to_3bit(ChLLRxDI(213));
  CNStageIntLLRInputS0xD(230)(3) <= LUT_4bit_to_3bit(ChLLRxDI(213));
  CNStageIntLLRInputS0xD(32)(3) <= LUT_4bit_to_3bit(ChLLRxDI(214));
  CNStageIntLLRInputS0xD(59)(3) <= LUT_4bit_to_3bit(ChLLRxDI(214));
  CNStageIntLLRInputS0xD(145)(3) <= LUT_4bit_to_3bit(ChLLRxDI(214));
  CNStageIntLLRInputS0xD(220)(3) <= LUT_4bit_to_3bit(ChLLRxDI(214));
  CNStageIntLLRInputS0xD(240)(3) <= LUT_4bit_to_3bit(ChLLRxDI(214));
  CNStageIntLLRInputS0xD(308)(3) <= LUT_4bit_to_3bit(ChLLRxDI(214));
  CNStageIntLLRInputS0xD(369)(3) <= LUT_4bit_to_3bit(ChLLRxDI(214));
  CNStageIntLLRInputS0xD(31)(3) <= LUT_4bit_to_3bit(ChLLRxDI(215));
  CNStageIntLLRInputS0xD(85)(3) <= LUT_4bit_to_3bit(ChLLRxDI(215));
  CNStageIntLLRInputS0xD(130)(3) <= LUT_4bit_to_3bit(ChLLRxDI(215));
  CNStageIntLLRInputS0xD(216)(3) <= LUT_4bit_to_3bit(ChLLRxDI(215));
  CNStageIntLLRInputS0xD(234)(3) <= LUT_4bit_to_3bit(ChLLRxDI(215));
  CNStageIntLLRInputS0xD(311)(3) <= LUT_4bit_to_3bit(ChLLRxDI(215));
  CNStageIntLLRInputS0xD(377)(3) <= LUT_4bit_to_3bit(ChLLRxDI(215));
  CNStageIntLLRInputS0xD(30)(3) <= LUT_4bit_to_3bit(ChLLRxDI(216));
  CNStageIntLLRInputS0xD(91)(3) <= LUT_4bit_to_3bit(ChLLRxDI(216));
  CNStageIntLLRInputS0xD(164)(3) <= LUT_4bit_to_3bit(ChLLRxDI(216));
  CNStageIntLLRInputS0xD(183)(3) <= LUT_4bit_to_3bit(ChLLRxDI(216));
  CNStageIntLLRInputS0xD(237)(3) <= LUT_4bit_to_3bit(ChLLRxDI(216));
  CNStageIntLLRInputS0xD(299)(3) <= LUT_4bit_to_3bit(ChLLRxDI(216));
  CNStageIntLLRInputS0xD(341)(3) <= LUT_4bit_to_3bit(ChLLRxDI(216));
  CNStageIntLLRInputS0xD(29)(3) <= LUT_4bit_to_3bit(ChLLRxDI(217));
  CNStageIntLLRInputS0xD(75)(3) <= LUT_4bit_to_3bit(ChLLRxDI(217));
  CNStageIntLLRInputS0xD(126)(3) <= LUT_4bit_to_3bit(ChLLRxDI(217));
  CNStageIntLLRInputS0xD(201)(3) <= LUT_4bit_to_3bit(ChLLRxDI(217));
  CNStageIntLLRInputS0xD(227)(3) <= LUT_4bit_to_3bit(ChLLRxDI(217));
  CNStageIntLLRInputS0xD(329)(3) <= LUT_4bit_to_3bit(ChLLRxDI(217));
  CNStageIntLLRInputS0xD(339)(3) <= LUT_4bit_to_3bit(ChLLRxDI(217));
  CNStageIntLLRInputS0xD(28)(3) <= LUT_4bit_to_3bit(ChLLRxDI(218));
  CNStageIntLLRInputS0xD(77)(3) <= LUT_4bit_to_3bit(ChLLRxDI(218));
  CNStageIntLLRInputS0xD(154)(3) <= LUT_4bit_to_3bit(ChLLRxDI(218));
  CNStageIntLLRInputS0xD(202)(3) <= LUT_4bit_to_3bit(ChLLRxDI(218));
  CNStageIntLLRInputS0xD(261)(3) <= LUT_4bit_to_3bit(ChLLRxDI(218));
  CNStageIntLLRInputS0xD(295)(3) <= LUT_4bit_to_3bit(ChLLRxDI(218));
  CNStageIntLLRInputS0xD(375)(3) <= LUT_4bit_to_3bit(ChLLRxDI(218));
  CNStageIntLLRInputS0xD(27)(3) <= LUT_4bit_to_3bit(ChLLRxDI(219));
  CNStageIntLLRInputS0xD(101)(3) <= LUT_4bit_to_3bit(ChLLRxDI(219));
  CNStageIntLLRInputS0xD(138)(3) <= LUT_4bit_to_3bit(ChLLRxDI(219));
  CNStageIntLLRInputS0xD(182)(3) <= LUT_4bit_to_3bit(ChLLRxDI(219));
  CNStageIntLLRInputS0xD(321)(3) <= LUT_4bit_to_3bit(ChLLRxDI(219));
  CNStageIntLLRInputS0xD(354)(3) <= LUT_4bit_to_3bit(ChLLRxDI(219));
  CNStageIntLLRInputS0xD(26)(3) <= LUT_4bit_to_3bit(ChLLRxDI(220));
  CNStageIntLLRInputS0xD(83)(3) <= LUT_4bit_to_3bit(ChLLRxDI(220));
  CNStageIntLLRInputS0xD(166)(3) <= LUT_4bit_to_3bit(ChLLRxDI(220));
  CNStageIntLLRInputS0xD(173)(3) <= LUT_4bit_to_3bit(ChLLRxDI(220));
  CNStageIntLLRInputS0xD(256)(3) <= LUT_4bit_to_3bit(ChLLRxDI(220));
  CNStageIntLLRInputS0xD(305)(3) <= LUT_4bit_to_3bit(ChLLRxDI(220));
  CNStageIntLLRInputS0xD(356)(3) <= LUT_4bit_to_3bit(ChLLRxDI(220));
  CNStageIntLLRInputS0xD(25)(3) <= LUT_4bit_to_3bit(ChLLRxDI(221));
  CNStageIntLLRInputS0xD(94)(3) <= LUT_4bit_to_3bit(ChLLRxDI(221));
  CNStageIntLLRInputS0xD(156)(3) <= LUT_4bit_to_3bit(ChLLRxDI(221));
  CNStageIntLLRInputS0xD(190)(3) <= LUT_4bit_to_3bit(ChLLRxDI(221));
  CNStageIntLLRInputS0xD(268)(3) <= LUT_4bit_to_3bit(ChLLRxDI(221));
  CNStageIntLLRInputS0xD(331)(3) <= LUT_4bit_to_3bit(ChLLRxDI(221));
  CNStageIntLLRInputS0xD(342)(3) <= LUT_4bit_to_3bit(ChLLRxDI(221));
  CNStageIntLLRInputS0xD(24)(3) <= LUT_4bit_to_3bit(ChLLRxDI(222));
  CNStageIntLLRInputS0xD(143)(3) <= LUT_4bit_to_3bit(ChLLRxDI(222));
  CNStageIntLLRInputS0xD(241)(3) <= LUT_4bit_to_3bit(ChLLRxDI(222));
  CNStageIntLLRInputS0xD(376)(3) <= LUT_4bit_to_3bit(ChLLRxDI(222));
  CNStageIntLLRInputS0xD(23)(3) <= LUT_4bit_to_3bit(ChLLRxDI(223));
  CNStageIntLLRInputS0xD(76)(3) <= LUT_4bit_to_3bit(ChLLRxDI(223));
  CNStageIntLLRInputS0xD(162)(3) <= LUT_4bit_to_3bit(ChLLRxDI(223));
  CNStageIntLLRInputS0xD(224)(3) <= LUT_4bit_to_3bit(ChLLRxDI(223));
  CNStageIntLLRInputS0xD(229)(3) <= LUT_4bit_to_3bit(ChLLRxDI(223));
  CNStageIntLLRInputS0xD(309)(3) <= LUT_4bit_to_3bit(ChLLRxDI(223));
  CNStageIntLLRInputS0xD(338)(3) <= LUT_4bit_to_3bit(ChLLRxDI(223));
  CNStageIntLLRInputS0xD(22)(3) <= LUT_4bit_to_3bit(ChLLRxDI(224));
  CNStageIntLLRInputS0xD(90)(3) <= LUT_4bit_to_3bit(ChLLRxDI(224));
  CNStageIntLLRInputS0xD(135)(3) <= LUT_4bit_to_3bit(ChLLRxDI(224));
  CNStageIntLLRInputS0xD(193)(3) <= LUT_4bit_to_3bit(ChLLRxDI(224));
  CNStageIntLLRInputS0xD(270)(3) <= LUT_4bit_to_3bit(ChLLRxDI(224));
  CNStageIntLLRInputS0xD(328)(3) <= LUT_4bit_to_3bit(ChLLRxDI(224));
  CNStageIntLLRInputS0xD(366)(3) <= LUT_4bit_to_3bit(ChLLRxDI(224));
  CNStageIntLLRInputS0xD(21)(3) <= LUT_4bit_to_3bit(ChLLRxDI(225));
  CNStageIntLLRInputS0xD(61)(3) <= LUT_4bit_to_3bit(ChLLRxDI(225));
  CNStageIntLLRInputS0xD(132)(3) <= LUT_4bit_to_3bit(ChLLRxDI(225));
  CNStageIntLLRInputS0xD(188)(3) <= LUT_4bit_to_3bit(ChLLRxDI(225));
  CNStageIntLLRInputS0xD(232)(3) <= LUT_4bit_to_3bit(ChLLRxDI(225));
  CNStageIntLLRInputS0xD(301)(3) <= LUT_4bit_to_3bit(ChLLRxDI(225));
  CNStageIntLLRInputS0xD(20)(3) <= LUT_4bit_to_3bit(ChLLRxDI(226));
  CNStageIntLLRInputS0xD(148)(3) <= LUT_4bit_to_3bit(ChLLRxDI(226));
  CNStageIntLLRInputS0xD(378)(3) <= LUT_4bit_to_3bit(ChLLRxDI(226));
  CNStageIntLLRInputS0xD(19)(3) <= LUT_4bit_to_3bit(ChLLRxDI(227));
  CNStageIntLLRInputS0xD(63)(3) <= LUT_4bit_to_3bit(ChLLRxDI(227));
  CNStageIntLLRInputS0xD(140)(3) <= LUT_4bit_to_3bit(ChLLRxDI(227));
  CNStageIntLLRInputS0xD(178)(3) <= LUT_4bit_to_3bit(ChLLRxDI(227));
  CNStageIntLLRInputS0xD(258)(3) <= LUT_4bit_to_3bit(ChLLRxDI(227));
  CNStageIntLLRInputS0xD(314)(3) <= LUT_4bit_to_3bit(ChLLRxDI(227));
  CNStageIntLLRInputS0xD(368)(3) <= LUT_4bit_to_3bit(ChLLRxDI(227));
  CNStageIntLLRInputS0xD(18)(3) <= LUT_4bit_to_3bit(ChLLRxDI(228));
  CNStageIntLLRInputS0xD(78)(3) <= LUT_4bit_to_3bit(ChLLRxDI(228));
  CNStageIntLLRInputS0xD(114)(3) <= LUT_4bit_to_3bit(ChLLRxDI(228));
  CNStageIntLLRInputS0xD(198)(3) <= LUT_4bit_to_3bit(ChLLRxDI(228));
  CNStageIntLLRInputS0xD(253)(3) <= LUT_4bit_to_3bit(ChLLRxDI(228));
  CNStageIntLLRInputS0xD(307)(3) <= LUT_4bit_to_3bit(ChLLRxDI(228));
  CNStageIntLLRInputS0xD(17)(3) <= LUT_4bit_to_3bit(ChLLRxDI(229));
  CNStageIntLLRInputS0xD(74)(3) <= LUT_4bit_to_3bit(ChLLRxDI(229));
  CNStageIntLLRInputS0xD(124)(3) <= LUT_4bit_to_3bit(ChLLRxDI(229));
  CNStageIntLLRInputS0xD(259)(3) <= LUT_4bit_to_3bit(ChLLRxDI(229));
  CNStageIntLLRInputS0xD(374)(3) <= LUT_4bit_to_3bit(ChLLRxDI(229));
  CNStageIntLLRInputS0xD(16)(3) <= LUT_4bit_to_3bit(ChLLRxDI(230));
  CNStageIntLLRInputS0xD(118)(3) <= LUT_4bit_to_3bit(ChLLRxDI(230));
  CNStageIntLLRInputS0xD(176)(3) <= LUT_4bit_to_3bit(ChLLRxDI(230));
  CNStageIntLLRInputS0xD(249)(3) <= LUT_4bit_to_3bit(ChLLRxDI(230));
  CNStageIntLLRInputS0xD(293)(3) <= LUT_4bit_to_3bit(ChLLRxDI(230));
  CNStageIntLLRInputS0xD(347)(3) <= LUT_4bit_to_3bit(ChLLRxDI(230));
  CNStageIntLLRInputS0xD(15)(3) <= LUT_4bit_to_3bit(ChLLRxDI(231));
  CNStageIntLLRInputS0xD(56)(3) <= LUT_4bit_to_3bit(ChLLRxDI(231));
  CNStageIntLLRInputS0xD(209)(3) <= LUT_4bit_to_3bit(ChLLRxDI(231));
  CNStageIntLLRInputS0xD(272)(3) <= LUT_4bit_to_3bit(ChLLRxDI(231));
  CNStageIntLLRInputS0xD(287)(3) <= LUT_4bit_to_3bit(ChLLRxDI(231));
  CNStageIntLLRInputS0xD(344)(3) <= LUT_4bit_to_3bit(ChLLRxDI(231));
  CNStageIntLLRInputS0xD(14)(3) <= LUT_4bit_to_3bit(ChLLRxDI(232));
  CNStageIntLLRInputS0xD(57)(3) <= LUT_4bit_to_3bit(ChLLRxDI(232));
  CNStageIntLLRInputS0xD(212)(3) <= LUT_4bit_to_3bit(ChLLRxDI(232));
  CNStageIntLLRInputS0xD(278)(3) <= LUT_4bit_to_3bit(ChLLRxDI(232));
  CNStageIntLLRInputS0xD(291)(3) <= LUT_4bit_to_3bit(ChLLRxDI(232));
  CNStageIntLLRInputS0xD(359)(3) <= LUT_4bit_to_3bit(ChLLRxDI(232));
  CNStageIntLLRInputS0xD(13)(3) <= LUT_4bit_to_3bit(ChLLRxDI(233));
  CNStageIntLLRInputS0xD(92)(3) <= LUT_4bit_to_3bit(ChLLRxDI(233));
  CNStageIntLLRInputS0xD(149)(3) <= LUT_4bit_to_3bit(ChLLRxDI(233));
  CNStageIntLLRInputS0xD(263)(3) <= LUT_4bit_to_3bit(ChLLRxDI(233));
  CNStageIntLLRInputS0xD(352)(3) <= LUT_4bit_to_3bit(ChLLRxDI(233));
  CNStageIntLLRInputS0xD(12)(3) <= LUT_4bit_to_3bit(ChLLRxDI(234));
  CNStageIntLLRInputS0xD(84)(3) <= LUT_4bit_to_3bit(ChLLRxDI(234));
  CNStageIntLLRInputS0xD(131)(3) <= LUT_4bit_to_3bit(ChLLRxDI(234));
  CNStageIntLLRInputS0xD(177)(3) <= LUT_4bit_to_3bit(ChLLRxDI(234));
  CNStageIntLLRInputS0xD(265)(3) <= LUT_4bit_to_3bit(ChLLRxDI(234));
  CNStageIntLLRInputS0xD(315)(3) <= LUT_4bit_to_3bit(ChLLRxDI(234));
  CNStageIntLLRInputS0xD(100)(3) <= LUT_4bit_to_3bit(ChLLRxDI(235));
  CNStageIntLLRInputS0xD(144)(3) <= LUT_4bit_to_3bit(ChLLRxDI(235));
  CNStageIntLLRInputS0xD(196)(3) <= LUT_4bit_to_3bit(ChLLRxDI(235));
  CNStageIntLLRInputS0xD(235)(3) <= LUT_4bit_to_3bit(ChLLRxDI(235));
  CNStageIntLLRInputS0xD(336)(3) <= LUT_4bit_to_3bit(ChLLRxDI(235));
  CNStageIntLLRInputS0xD(11)(3) <= LUT_4bit_to_3bit(ChLLRxDI(236));
  CNStageIntLLRInputS0xD(104)(3) <= LUT_4bit_to_3bit(ChLLRxDI(236));
  CNStageIntLLRInputS0xD(155)(3) <= LUT_4bit_to_3bit(ChLLRxDI(236));
  CNStageIntLLRInputS0xD(221)(3) <= LUT_4bit_to_3bit(ChLLRxDI(236));
  CNStageIntLLRInputS0xD(271)(3) <= LUT_4bit_to_3bit(ChLLRxDI(236));
  CNStageIntLLRInputS0xD(310)(3) <= LUT_4bit_to_3bit(ChLLRxDI(236));
  CNStageIntLLRInputS0xD(10)(3) <= LUT_4bit_to_3bit(ChLLRxDI(237));
  CNStageIntLLRInputS0xD(110)(3) <= LUT_4bit_to_3bit(ChLLRxDI(237));
  CNStageIntLLRInputS0xD(125)(3) <= LUT_4bit_to_3bit(ChLLRxDI(237));
  CNStageIntLLRInputS0xD(228)(3) <= LUT_4bit_to_3bit(ChLLRxDI(237));
  CNStageIntLLRInputS0xD(322)(3) <= LUT_4bit_to_3bit(ChLLRxDI(237));
  CNStageIntLLRInputS0xD(334)(3) <= LUT_4bit_to_3bit(ChLLRxDI(237));
  CNStageIntLLRInputS0xD(9)(3) <= LUT_4bit_to_3bit(ChLLRxDI(238));
  CNStageIntLLRInputS0xD(103)(3) <= LUT_4bit_to_3bit(ChLLRxDI(238));
  CNStageIntLLRInputS0xD(113)(3) <= LUT_4bit_to_3bit(ChLLRxDI(238));
  CNStageIntLLRInputS0xD(179)(3) <= LUT_4bit_to_3bit(ChLLRxDI(238));
  CNStageIntLLRInputS0xD(236)(3) <= LUT_4bit_to_3bit(ChLLRxDI(238));
  CNStageIntLLRInputS0xD(294)(3) <= LUT_4bit_to_3bit(ChLLRxDI(238));
  CNStageIntLLRInputS0xD(383)(3) <= LUT_4bit_to_3bit(ChLLRxDI(238));
  CNStageIntLLRInputS0xD(8)(3) <= LUT_4bit_to_3bit(ChLLRxDI(239));
  CNStageIntLLRInputS0xD(98)(3) <= LUT_4bit_to_3bit(ChLLRxDI(239));
  CNStageIntLLRInputS0xD(158)(3) <= LUT_4bit_to_3bit(ChLLRxDI(239));
  CNStageIntLLRInputS0xD(223)(3) <= LUT_4bit_to_3bit(ChLLRxDI(239));
  CNStageIntLLRInputS0xD(264)(3) <= LUT_4bit_to_3bit(ChLLRxDI(239));
  CNStageIntLLRInputS0xD(284)(3) <= LUT_4bit_to_3bit(ChLLRxDI(239));
  CNStageIntLLRInputS0xD(360)(3) <= LUT_4bit_to_3bit(ChLLRxDI(239));
  CNStageIntLLRInputS0xD(7)(3) <= LUT_4bit_to_3bit(ChLLRxDI(240));
  CNStageIntLLRInputS0xD(81)(3) <= LUT_4bit_to_3bit(ChLLRxDI(240));
  CNStageIntLLRInputS0xD(116)(3) <= LUT_4bit_to_3bit(ChLLRxDI(240));
  CNStageIntLLRInputS0xD(210)(3) <= LUT_4bit_to_3bit(ChLLRxDI(240));
  CNStageIntLLRInputS0xD(277)(3) <= LUT_4bit_to_3bit(ChLLRxDI(240));
  CNStageIntLLRInputS0xD(324)(3) <= LUT_4bit_to_3bit(ChLLRxDI(240));
  CNStageIntLLRInputS0xD(343)(3) <= LUT_4bit_to_3bit(ChLLRxDI(240));
  CNStageIntLLRInputS0xD(6)(3) <= LUT_4bit_to_3bit(ChLLRxDI(241));
  CNStageIntLLRInputS0xD(88)(3) <= LUT_4bit_to_3bit(ChLLRxDI(241));
  CNStageIntLLRInputS0xD(175)(3) <= LUT_4bit_to_3bit(ChLLRxDI(241));
  CNStageIntLLRInputS0xD(250)(3) <= LUT_4bit_to_3bit(ChLLRxDI(241));
  CNStageIntLLRInputS0xD(285)(3) <= LUT_4bit_to_3bit(ChLLRxDI(241));
  CNStageIntLLRInputS0xD(355)(3) <= LUT_4bit_to_3bit(ChLLRxDI(241));
  CNStageIntLLRInputS0xD(5)(3) <= LUT_4bit_to_3bit(ChLLRxDI(242));
  CNStageIntLLRInputS0xD(108)(3) <= LUT_4bit_to_3bit(ChLLRxDI(242));
  CNStageIntLLRInputS0xD(146)(3) <= LUT_4bit_to_3bit(ChLLRxDI(242));
  CNStageIntLLRInputS0xD(203)(3) <= LUT_4bit_to_3bit(ChLLRxDI(242));
  CNStageIntLLRInputS0xD(231)(3) <= LUT_4bit_to_3bit(ChLLRxDI(242));
  CNStageIntLLRInputS0xD(303)(3) <= LUT_4bit_to_3bit(ChLLRxDI(242));
  CNStageIntLLRInputS0xD(367)(3) <= LUT_4bit_to_3bit(ChLLRxDI(242));
  CNStageIntLLRInputS0xD(4)(3) <= LUT_4bit_to_3bit(ChLLRxDI(243));
  CNStageIntLLRInputS0xD(106)(3) <= LUT_4bit_to_3bit(ChLLRxDI(243));
  CNStageIntLLRInputS0xD(141)(3) <= LUT_4bit_to_3bit(ChLLRxDI(243));
  CNStageIntLLRInputS0xD(200)(3) <= LUT_4bit_to_3bit(ChLLRxDI(243));
  CNStageIntLLRInputS0xD(252)(3) <= LUT_4bit_to_3bit(ChLLRxDI(243));
  CNStageIntLLRInputS0xD(312)(3) <= LUT_4bit_to_3bit(ChLLRxDI(243));
  CNStageIntLLRInputS0xD(337)(3) <= LUT_4bit_to_3bit(ChLLRxDI(243));
  CNStageIntLLRInputS0xD(147)(3) <= LUT_4bit_to_3bit(ChLLRxDI(244));
  CNStageIntLLRInputS0xD(266)(3) <= LUT_4bit_to_3bit(ChLLRxDI(244));
  CNStageIntLLRInputS0xD(3)(3) <= LUT_4bit_to_3bit(ChLLRxDI(245));
  CNStageIntLLRInputS0xD(66)(3) <= LUT_4bit_to_3bit(ChLLRxDI(245));
  CNStageIntLLRInputS0xD(136)(3) <= LUT_4bit_to_3bit(ChLLRxDI(245));
  CNStageIntLLRInputS0xD(207)(3) <= LUT_4bit_to_3bit(ChLLRxDI(245));
  CNStageIntLLRInputS0xD(262)(3) <= LUT_4bit_to_3bit(ChLLRxDI(245));
  CNStageIntLLRInputS0xD(313)(3) <= LUT_4bit_to_3bit(ChLLRxDI(245));
  CNStageIntLLRInputS0xD(370)(3) <= LUT_4bit_to_3bit(ChLLRxDI(245));
  CNStageIntLLRInputS0xD(2)(3) <= LUT_4bit_to_3bit(ChLLRxDI(246));
  CNStageIntLLRInputS0xD(69)(3) <= LUT_4bit_to_3bit(ChLLRxDI(246));
  CNStageIntLLRInputS0xD(161)(3) <= LUT_4bit_to_3bit(ChLLRxDI(246));
  CNStageIntLLRInputS0xD(185)(3) <= LUT_4bit_to_3bit(ChLLRxDI(246));
  CNStageIntLLRInputS0xD(226)(3) <= LUT_4bit_to_3bit(ChLLRxDI(246));
  CNStageIntLLRInputS0xD(302)(3) <= LUT_4bit_to_3bit(ChLLRxDI(246));
  CNStageIntLLRInputS0xD(1)(3) <= LUT_4bit_to_3bit(ChLLRxDI(247));
  CNStageIntLLRInputS0xD(109)(3) <= LUT_4bit_to_3bit(ChLLRxDI(247));
  CNStageIntLLRInputS0xD(168)(3) <= LUT_4bit_to_3bit(ChLLRxDI(247));
  CNStageIntLLRInputS0xD(194)(3) <= LUT_4bit_to_3bit(ChLLRxDI(247));
  CNStageIntLLRInputS0xD(247)(3) <= LUT_4bit_to_3bit(ChLLRxDI(247));
  CNStageIntLLRInputS0xD(327)(3) <= LUT_4bit_to_3bit(ChLLRxDI(247));
  CNStageIntLLRInputS0xD(349)(3) <= LUT_4bit_to_3bit(ChLLRxDI(247));
  CNStageIntLLRInputS0xD(0)(3) <= LUT_4bit_to_3bit(ChLLRxDI(248));
  CNStageIntLLRInputS0xD(87)(3) <= LUT_4bit_to_3bit(ChLLRxDI(248));
  CNStageIntLLRInputS0xD(151)(3) <= LUT_4bit_to_3bit(ChLLRxDI(248));
  CNStageIntLLRInputS0xD(189)(3) <= LUT_4bit_to_3bit(ChLLRxDI(248));
  CNStageIntLLRInputS0xD(248)(3) <= LUT_4bit_to_3bit(ChLLRxDI(248));
  CNStageIntLLRInputS0xD(280)(3) <= LUT_4bit_to_3bit(ChLLRxDI(248));
  CNStageIntLLRInputS0xD(357)(3) <= LUT_4bit_to_3bit(ChLLRxDI(248));
  CNStageIntLLRInputS0xD(152)(3) <= LUT_4bit_to_3bit(ChLLRxDI(249));
  CNStageIntLLRInputS0xD(192)(3) <= LUT_4bit_to_3bit(ChLLRxDI(249));
  CNStageIntLLRInputS0xD(225)(3) <= LUT_4bit_to_3bit(ChLLRxDI(249));
  CNStageIntLLRInputS0xD(317)(3) <= LUT_4bit_to_3bit(ChLLRxDI(249));
  CNStageIntLLRInputS0xD(353)(3) <= LUT_4bit_to_3bit(ChLLRxDI(249));
  CNStageIntLLRInputS0xD(79)(3) <= LUT_4bit_to_3bit(ChLLRxDI(250));
  CNStageIntLLRInputS0xD(120)(3) <= LUT_4bit_to_3bit(ChLLRxDI(250));
  CNStageIntLLRInputS0xD(184)(3) <= LUT_4bit_to_3bit(ChLLRxDI(250));
  CNStageIntLLRInputS0xD(319)(3) <= LUT_4bit_to_3bit(ChLLRxDI(250));
  CNStageIntLLRInputS0xD(358)(3) <= LUT_4bit_to_3bit(ChLLRxDI(250));
  CNStageIntLLRInputS0xD(62)(3) <= LUT_4bit_to_3bit(ChLLRxDI(251));
  CNStageIntLLRInputS0xD(159)(3) <= LUT_4bit_to_3bit(ChLLRxDI(251));
  CNStageIntLLRInputS0xD(215)(3) <= LUT_4bit_to_3bit(ChLLRxDI(251));
  CNStageIntLLRInputS0xD(289)(3) <= LUT_4bit_to_3bit(ChLLRxDI(251));
  CNStageIntLLRInputS0xD(348)(3) <= LUT_4bit_to_3bit(ChLLRxDI(251));
  CNStageIntLLRInputS0xD(89)(3) <= LUT_4bit_to_3bit(ChLLRxDI(252));
  CNStageIntLLRInputS0xD(112)(3) <= LUT_4bit_to_3bit(ChLLRxDI(252));
  CNStageIntLLRInputS0xD(199)(3) <= LUT_4bit_to_3bit(ChLLRxDI(252));
  CNStageIntLLRInputS0xD(239)(3) <= LUT_4bit_to_3bit(ChLLRxDI(252));
  CNStageIntLLRInputS0xD(325)(3) <= LUT_4bit_to_3bit(ChLLRxDI(252));
  CNStageIntLLRInputS0xD(373)(3) <= LUT_4bit_to_3bit(ChLLRxDI(252));
  CNStageIntLLRInputS0xD(80)(3) <= LUT_4bit_to_3bit(ChLLRxDI(253));
  CNStageIntLLRInputS0xD(121)(3) <= LUT_4bit_to_3bit(ChLLRxDI(253));
  CNStageIntLLRInputS0xD(211)(3) <= LUT_4bit_to_3bit(ChLLRxDI(253));
  CNStageIntLLRInputS0xD(279)(3) <= LUT_4bit_to_3bit(ChLLRxDI(253));
  CNStageIntLLRInputS0xD(283)(3) <= LUT_4bit_to_3bit(ChLLRxDI(253));
  CNStageIntLLRInputS0xD(380)(3) <= LUT_4bit_to_3bit(ChLLRxDI(253));
  CNStageIntLLRInputS0xD(67)(3) <= LUT_4bit_to_3bit(ChLLRxDI(254));
  CNStageIntLLRInputS0xD(222)(3) <= LUT_4bit_to_3bit(ChLLRxDI(254));
  CNStageIntLLRInputS0xD(238)(3) <= LUT_4bit_to_3bit(ChLLRxDI(254));
  CNStageIntLLRInputS0xD(290)(3) <= LUT_4bit_to_3bit(ChLLRxDI(254));
  CNStageIntLLRInputS0xD(362)(3) <= LUT_4bit_to_3bit(ChLLRxDI(254));
  CNStageIntLLRInputS0xD(52)(3) <= LUT_4bit_to_3bit(ChLLRxDI(255));
  CNStageIntLLRInputS0xD(86)(3) <= LUT_4bit_to_3bit(ChLLRxDI(255));
  CNStageIntLLRInputS0xD(167)(3) <= LUT_4bit_to_3bit(ChLLRxDI(255));
  CNStageIntLLRInputS0xD(195)(3) <= LUT_4bit_to_3bit(ChLLRxDI(255));
  CNStageIntLLRInputS0xD(233)(3) <= LUT_4bit_to_3bit(ChLLRxDI(255));
  CNStageIntLLRInputS0xD(318)(3) <= LUT_4bit_to_3bit(ChLLRxDI(255));
  CNStageIntLLRInputS0xD(364)(3) <= LUT_4bit_to_3bit(ChLLRxDI(255));
  CNStageIntLLRInputS0xD(53)(4) <= LUT_4bit_to_3bit(ChLLRxDI(256));
  CNStageIntLLRInputS0xD(106)(4) <= LUT_4bit_to_3bit(ChLLRxDI(256));
  CNStageIntLLRInputS0xD(127)(4) <= LUT_4bit_to_3bit(ChLLRxDI(256));
  CNStageIntLLRInputS0xD(242)(4) <= LUT_4bit_to_3bit(ChLLRxDI(256));
  CNStageIntLLRInputS0xD(296)(4) <= LUT_4bit_to_3bit(ChLLRxDI(256));
  CNStageIntLLRInputS0xD(339)(4) <= LUT_4bit_to_3bit(ChLLRxDI(256));
  CNStageIntLLRInputS0xD(51)(4) <= LUT_4bit_to_3bit(ChLLRxDI(257));
  CNStageIntLLRInputS0xD(85)(4) <= LUT_4bit_to_3bit(ChLLRxDI(257));
  CNStageIntLLRInputS0xD(166)(4) <= LUT_4bit_to_3bit(ChLLRxDI(257));
  CNStageIntLLRInputS0xD(194)(4) <= LUT_4bit_to_3bit(ChLLRxDI(257));
  CNStageIntLLRInputS0xD(232)(4) <= LUT_4bit_to_3bit(ChLLRxDI(257));
  CNStageIntLLRInputS0xD(317)(4) <= LUT_4bit_to_3bit(ChLLRxDI(257));
  CNStageIntLLRInputS0xD(363)(4) <= LUT_4bit_to_3bit(ChLLRxDI(257));
  CNStageIntLLRInputS0xD(50)(4) <= LUT_4bit_to_3bit(ChLLRxDI(258));
  CNStageIntLLRInputS0xD(57)(4) <= LUT_4bit_to_3bit(ChLLRxDI(258));
  CNStageIntLLRInputS0xD(331)(4) <= LUT_4bit_to_3bit(ChLLRxDI(258));
  CNStageIntLLRInputS0xD(54)(4) <= LUT_4bit_to_3bit(ChLLRxDI(259));
  CNStageIntLLRInputS0xD(114)(4) <= LUT_4bit_to_3bit(ChLLRxDI(259));
  CNStageIntLLRInputS0xD(274)(4) <= LUT_4bit_to_3bit(ChLLRxDI(259));
  CNStageIntLLRInputS0xD(303)(4) <= LUT_4bit_to_3bit(ChLLRxDI(259));
  CNStageIntLLRInputS0xD(370)(4) <= LUT_4bit_to_3bit(ChLLRxDI(259));
  CNStageIntLLRInputS0xD(49)(4) <= LUT_4bit_to_3bit(ChLLRxDI(260));
  CNStageIntLLRInputS0xD(71)(4) <= LUT_4bit_to_3bit(ChLLRxDI(260));
  CNStageIntLLRInputS0xD(138)(4) <= LUT_4bit_to_3bit(ChLLRxDI(260));
  CNStageIntLLRInputS0xD(186)(4) <= LUT_4bit_to_3bit(ChLLRxDI(260));
  CNStageIntLLRInputS0xD(243)(4) <= LUT_4bit_to_3bit(ChLLRxDI(260));
  CNStageIntLLRInputS0xD(383)(4) <= LUT_4bit_to_3bit(ChLLRxDI(260));
  CNStageIntLLRInputS0xD(48)(4) <= LUT_4bit_to_3bit(ChLLRxDI(261));
  CNStageIntLLRInputS0xD(63)(4) <= LUT_4bit_to_3bit(ChLLRxDI(261));
  CNStageIntLLRInputS0xD(152)(4) <= LUT_4bit_to_3bit(ChLLRxDI(261));
  CNStageIntLLRInputS0xD(204)(4) <= LUT_4bit_to_3bit(ChLLRxDI(261));
  CNStageIntLLRInputS0xD(305)(4) <= LUT_4bit_to_3bit(ChLLRxDI(261));
  CNStageIntLLRInputS0xD(333)(4) <= LUT_4bit_to_3bit(ChLLRxDI(261));
  CNStageIntLLRInputS0xD(47)(4) <= LUT_4bit_to_3bit(ChLLRxDI(262));
  CNStageIntLLRInputS0xD(95)(4) <= LUT_4bit_to_3bit(ChLLRxDI(262));
  CNStageIntLLRInputS0xD(149)(4) <= LUT_4bit_to_3bit(ChLLRxDI(262));
  CNStageIntLLRInputS0xD(212)(4) <= LUT_4bit_to_3bit(ChLLRxDI(262));
  CNStageIntLLRInputS0xD(319)(4) <= LUT_4bit_to_3bit(ChLLRxDI(262));
  CNStageIntLLRInputS0xD(362)(4) <= LUT_4bit_to_3bit(ChLLRxDI(262));
  CNStageIntLLRInputS0xD(46)(4) <= LUT_4bit_to_3bit(ChLLRxDI(263));
  CNStageIntLLRInputS0xD(104)(4) <= LUT_4bit_to_3bit(ChLLRxDI(263));
  CNStageIntLLRInputS0xD(169)(4) <= LUT_4bit_to_3bit(ChLLRxDI(263));
  CNStageIntLLRInputS0xD(207)(4) <= LUT_4bit_to_3bit(ChLLRxDI(263));
  CNStageIntLLRInputS0xD(253)(4) <= LUT_4bit_to_3bit(ChLLRxDI(263));
  CNStageIntLLRInputS0xD(315)(4) <= LUT_4bit_to_3bit(ChLLRxDI(263));
  CNStageIntLLRInputS0xD(378)(4) <= LUT_4bit_to_3bit(ChLLRxDI(263));
  CNStageIntLLRInputS0xD(45)(4) <= LUT_4bit_to_3bit(ChLLRxDI(264));
  CNStageIntLLRInputS0xD(98)(4) <= LUT_4bit_to_3bit(ChLLRxDI(264));
  CNStageIntLLRInputS0xD(132)(4) <= LUT_4bit_to_3bit(ChLLRxDI(264));
  CNStageIntLLRInputS0xD(213)(4) <= LUT_4bit_to_3bit(ChLLRxDI(264));
  CNStageIntLLRInputS0xD(256)(4) <= LUT_4bit_to_3bit(ChLLRxDI(264));
  CNStageIntLLRInputS0xD(281)(4) <= LUT_4bit_to_3bit(ChLLRxDI(264));
  CNStageIntLLRInputS0xD(349)(4) <= LUT_4bit_to_3bit(ChLLRxDI(264));
  CNStageIntLLRInputS0xD(44)(4) <= LUT_4bit_to_3bit(ChLLRxDI(265));
  CNStageIntLLRInputS0xD(133)(4) <= LUT_4bit_to_3bit(ChLLRxDI(265));
  CNStageIntLLRInputS0xD(203)(4) <= LUT_4bit_to_3bit(ChLLRxDI(265));
  CNStageIntLLRInputS0xD(244)(4) <= LUT_4bit_to_3bit(ChLLRxDI(265));
  CNStageIntLLRInputS0xD(43)(4) <= LUT_4bit_to_3bit(ChLLRxDI(266));
  CNStageIntLLRInputS0xD(168)(4) <= LUT_4bit_to_3bit(ChLLRxDI(266));
  CNStageIntLLRInputS0xD(173)(4) <= LUT_4bit_to_3bit(ChLLRxDI(266));
  CNStageIntLLRInputS0xD(273)(4) <= LUT_4bit_to_3bit(ChLLRxDI(266));
  CNStageIntLLRInputS0xD(300)(4) <= LUT_4bit_to_3bit(ChLLRxDI(266));
  CNStageIntLLRInputS0xD(42)(4) <= LUT_4bit_to_3bit(ChLLRxDI(267));
  CNStageIntLLRInputS0xD(72)(4) <= LUT_4bit_to_3bit(ChLLRxDI(267));
  CNStageIntLLRInputS0xD(159)(4) <= LUT_4bit_to_3bit(ChLLRxDI(267));
  CNStageIntLLRInputS0xD(180)(4) <= LUT_4bit_to_3bit(ChLLRxDI(267));
  CNStageIntLLRInputS0xD(241)(4) <= LUT_4bit_to_3bit(ChLLRxDI(267));
  CNStageIntLLRInputS0xD(280)(4) <= LUT_4bit_to_3bit(ChLLRxDI(267));
  CNStageIntLLRInputS0xD(364)(4) <= LUT_4bit_to_3bit(ChLLRxDI(267));
  CNStageIntLLRInputS0xD(41)(4) <= LUT_4bit_to_3bit(ChLLRxDI(268));
  CNStageIntLLRInputS0xD(109)(4) <= LUT_4bit_to_3bit(ChLLRxDI(268));
  CNStageIntLLRInputS0xD(118)(4) <= LUT_4bit_to_3bit(ChLLRxDI(268));
  CNStageIntLLRInputS0xD(216)(4) <= LUT_4bit_to_3bit(ChLLRxDI(268));
  CNStageIntLLRInputS0xD(266)(4) <= LUT_4bit_to_3bit(ChLLRxDI(268));
  CNStageIntLLRInputS0xD(325)(4) <= LUT_4bit_to_3bit(ChLLRxDI(268));
  CNStageIntLLRInputS0xD(360)(4) <= LUT_4bit_to_3bit(ChLLRxDI(268));
  CNStageIntLLRInputS0xD(67)(4) <= LUT_4bit_to_3bit(ChLLRxDI(269));
  CNStageIntLLRInputS0xD(122)(4) <= LUT_4bit_to_3bit(ChLLRxDI(269));
  CNStageIntLLRInputS0xD(218)(4) <= LUT_4bit_to_3bit(ChLLRxDI(269));
  CNStageIntLLRInputS0xD(250)(4) <= LUT_4bit_to_3bit(ChLLRxDI(269));
  CNStageIntLLRInputS0xD(287)(4) <= LUT_4bit_to_3bit(ChLLRxDI(269));
  CNStageIntLLRInputS0xD(381)(4) <= LUT_4bit_to_3bit(ChLLRxDI(269));
  CNStageIntLLRInputS0xD(40)(4) <= LUT_4bit_to_3bit(ChLLRxDI(270));
  CNStageIntLLRInputS0xD(79)(4) <= LUT_4bit_to_3bit(ChLLRxDI(270));
  CNStageIntLLRInputS0xD(170)(4) <= LUT_4bit_to_3bit(ChLLRxDI(270));
  CNStageIntLLRInputS0xD(190)(4) <= LUT_4bit_to_3bit(ChLLRxDI(270));
  CNStageIntLLRInputS0xD(275)(4) <= LUT_4bit_to_3bit(ChLLRxDI(270));
  CNStageIntLLRInputS0xD(292)(4) <= LUT_4bit_to_3bit(ChLLRxDI(270));
  CNStageIntLLRInputS0xD(344)(4) <= LUT_4bit_to_3bit(ChLLRxDI(270));
  CNStageIntLLRInputS0xD(39)(4) <= LUT_4bit_to_3bit(ChLLRxDI(271));
  CNStageIntLLRInputS0xD(105)(4) <= LUT_4bit_to_3bit(ChLLRxDI(271));
  CNStageIntLLRInputS0xD(171)(4) <= LUT_4bit_to_3bit(ChLLRxDI(271));
  CNStageIntLLRInputS0xD(268)(4) <= LUT_4bit_to_3bit(ChLLRxDI(271));
  CNStageIntLLRInputS0xD(332)(4) <= LUT_4bit_to_3bit(ChLLRxDI(271));
  CNStageIntLLRInputS0xD(345)(4) <= LUT_4bit_to_3bit(ChLLRxDI(271));
  CNStageIntLLRInputS0xD(38)(4) <= LUT_4bit_to_3bit(ChLLRxDI(272));
  CNStageIntLLRInputS0xD(94)(4) <= LUT_4bit_to_3bit(ChLLRxDI(272));
  CNStageIntLLRInputS0xD(116)(4) <= LUT_4bit_to_3bit(ChLLRxDI(272));
  CNStageIntLLRInputS0xD(184)(4) <= LUT_4bit_to_3bit(ChLLRxDI(272));
  CNStageIntLLRInputS0xD(254)(4) <= LUT_4bit_to_3bit(ChLLRxDI(272));
  CNStageIntLLRInputS0xD(291)(4) <= LUT_4bit_to_3bit(ChLLRxDI(272));
  CNStageIntLLRInputS0xD(380)(4) <= LUT_4bit_to_3bit(ChLLRxDI(272));
  CNStageIntLLRInputS0xD(37)(4) <= LUT_4bit_to_3bit(ChLLRxDI(273));
  CNStageIntLLRInputS0xD(81)(4) <= LUT_4bit_to_3bit(ChLLRxDI(273));
  CNStageIntLLRInputS0xD(156)(4) <= LUT_4bit_to_3bit(ChLLRxDI(273));
  CNStageIntLLRInputS0xD(272)(4) <= LUT_4bit_to_3bit(ChLLRxDI(273));
  CNStageIntLLRInputS0xD(285)(4) <= LUT_4bit_to_3bit(ChLLRxDI(273));
  CNStageIntLLRInputS0xD(371)(4) <= LUT_4bit_to_3bit(ChLLRxDI(273));
  CNStageIntLLRInputS0xD(36)(4) <= LUT_4bit_to_3bit(ChLLRxDI(274));
  CNStageIntLLRInputS0xD(164)(4) <= LUT_4bit_to_3bit(ChLLRxDI(274));
  CNStageIntLLRInputS0xD(217)(4) <= LUT_4bit_to_3bit(ChLLRxDI(274));
  CNStageIntLLRInputS0xD(248)(4) <= LUT_4bit_to_3bit(ChLLRxDI(274));
  CNStageIntLLRInputS0xD(35)(4) <= LUT_4bit_to_3bit(ChLLRxDI(275));
  CNStageIntLLRInputS0xD(59)(4) <= LUT_4bit_to_3bit(ChLLRxDI(275));
  CNStageIntLLRInputS0xD(128)(4) <= LUT_4bit_to_3bit(ChLLRxDI(275));
  CNStageIntLLRInputS0xD(179)(4) <= LUT_4bit_to_3bit(ChLLRxDI(275));
  CNStageIntLLRInputS0xD(329)(4) <= LUT_4bit_to_3bit(ChLLRxDI(275));
  CNStageIntLLRInputS0xD(34)(4) <= LUT_4bit_to_3bit(ChLLRxDI(276));
  CNStageIntLLRInputS0xD(69)(4) <= LUT_4bit_to_3bit(ChLLRxDI(276));
  CNStageIntLLRInputS0xD(126)(4) <= LUT_4bit_to_3bit(ChLLRxDI(276));
  CNStageIntLLRInputS0xD(205)(4) <= LUT_4bit_to_3bit(ChLLRxDI(276));
  CNStageIntLLRInputS0xD(259)(4) <= LUT_4bit_to_3bit(ChLLRxDI(276));
  CNStageIntLLRInputS0xD(297)(4) <= LUT_4bit_to_3bit(ChLLRxDI(276));
  CNStageIntLLRInputS0xD(33)(4) <= LUT_4bit_to_3bit(ChLLRxDI(277));
  CNStageIntLLRInputS0xD(64)(4) <= LUT_4bit_to_3bit(ChLLRxDI(277));
  CNStageIntLLRInputS0xD(162)(4) <= LUT_4bit_to_3bit(ChLLRxDI(277));
  CNStageIntLLRInputS0xD(185)(4) <= LUT_4bit_to_3bit(ChLLRxDI(277));
  CNStageIntLLRInputS0xD(252)(4) <= LUT_4bit_to_3bit(ChLLRxDI(277));
  CNStageIntLLRInputS0xD(295)(4) <= LUT_4bit_to_3bit(ChLLRxDI(277));
  CNStageIntLLRInputS0xD(334)(4) <= LUT_4bit_to_3bit(ChLLRxDI(277));
  CNStageIntLLRInputS0xD(32)(4) <= LUT_4bit_to_3bit(ChLLRxDI(278));
  CNStageIntLLRInputS0xD(70)(4) <= LUT_4bit_to_3bit(ChLLRxDI(278));
  CNStageIntLLRInputS0xD(141)(4) <= LUT_4bit_to_3bit(ChLLRxDI(278));
  CNStageIntLLRInputS0xD(229)(4) <= LUT_4bit_to_3bit(ChLLRxDI(278));
  CNStageIntLLRInputS0xD(328)(4) <= LUT_4bit_to_3bit(ChLLRxDI(278));
  CNStageIntLLRInputS0xD(31)(4) <= LUT_4bit_to_3bit(ChLLRxDI(279));
  CNStageIntLLRInputS0xD(58)(4) <= LUT_4bit_to_3bit(ChLLRxDI(279));
  CNStageIntLLRInputS0xD(144)(4) <= LUT_4bit_to_3bit(ChLLRxDI(279));
  CNStageIntLLRInputS0xD(219)(4) <= LUT_4bit_to_3bit(ChLLRxDI(279));
  CNStageIntLLRInputS0xD(239)(4) <= LUT_4bit_to_3bit(ChLLRxDI(279));
  CNStageIntLLRInputS0xD(368)(4) <= LUT_4bit_to_3bit(ChLLRxDI(279));
  CNStageIntLLRInputS0xD(30)(4) <= LUT_4bit_to_3bit(ChLLRxDI(280));
  CNStageIntLLRInputS0xD(84)(4) <= LUT_4bit_to_3bit(ChLLRxDI(280));
  CNStageIntLLRInputS0xD(129)(4) <= LUT_4bit_to_3bit(ChLLRxDI(280));
  CNStageIntLLRInputS0xD(215)(4) <= LUT_4bit_to_3bit(ChLLRxDI(280));
  CNStageIntLLRInputS0xD(233)(4) <= LUT_4bit_to_3bit(ChLLRxDI(280));
  CNStageIntLLRInputS0xD(310)(4) <= LUT_4bit_to_3bit(ChLLRxDI(280));
  CNStageIntLLRInputS0xD(376)(4) <= LUT_4bit_to_3bit(ChLLRxDI(280));
  CNStageIntLLRInputS0xD(29)(4) <= LUT_4bit_to_3bit(ChLLRxDI(281));
  CNStageIntLLRInputS0xD(90)(4) <= LUT_4bit_to_3bit(ChLLRxDI(281));
  CNStageIntLLRInputS0xD(163)(4) <= LUT_4bit_to_3bit(ChLLRxDI(281));
  CNStageIntLLRInputS0xD(182)(4) <= LUT_4bit_to_3bit(ChLLRxDI(281));
  CNStageIntLLRInputS0xD(236)(4) <= LUT_4bit_to_3bit(ChLLRxDI(281));
  CNStageIntLLRInputS0xD(298)(4) <= LUT_4bit_to_3bit(ChLLRxDI(281));
  CNStageIntLLRInputS0xD(340)(4) <= LUT_4bit_to_3bit(ChLLRxDI(281));
  CNStageIntLLRInputS0xD(28)(4) <= LUT_4bit_to_3bit(ChLLRxDI(282));
  CNStageIntLLRInputS0xD(74)(4) <= LUT_4bit_to_3bit(ChLLRxDI(282));
  CNStageIntLLRInputS0xD(125)(4) <= LUT_4bit_to_3bit(ChLLRxDI(282));
  CNStageIntLLRInputS0xD(200)(4) <= LUT_4bit_to_3bit(ChLLRxDI(282));
  CNStageIntLLRInputS0xD(226)(4) <= LUT_4bit_to_3bit(ChLLRxDI(282));
  CNStageIntLLRInputS0xD(338)(4) <= LUT_4bit_to_3bit(ChLLRxDI(282));
  CNStageIntLLRInputS0xD(27)(4) <= LUT_4bit_to_3bit(ChLLRxDI(283));
  CNStageIntLLRInputS0xD(76)(4) <= LUT_4bit_to_3bit(ChLLRxDI(283));
  CNStageIntLLRInputS0xD(153)(4) <= LUT_4bit_to_3bit(ChLLRxDI(283));
  CNStageIntLLRInputS0xD(201)(4) <= LUT_4bit_to_3bit(ChLLRxDI(283));
  CNStageIntLLRInputS0xD(260)(4) <= LUT_4bit_to_3bit(ChLLRxDI(283));
  CNStageIntLLRInputS0xD(294)(4) <= LUT_4bit_to_3bit(ChLLRxDI(283));
  CNStageIntLLRInputS0xD(374)(4) <= LUT_4bit_to_3bit(ChLLRxDI(283));
  CNStageIntLLRInputS0xD(26)(4) <= LUT_4bit_to_3bit(ChLLRxDI(284));
  CNStageIntLLRInputS0xD(100)(4) <= LUT_4bit_to_3bit(ChLLRxDI(284));
  CNStageIntLLRInputS0xD(137)(4) <= LUT_4bit_to_3bit(ChLLRxDI(284));
  CNStageIntLLRInputS0xD(181)(4) <= LUT_4bit_to_3bit(ChLLRxDI(284));
  CNStageIntLLRInputS0xD(245)(4) <= LUT_4bit_to_3bit(ChLLRxDI(284));
  CNStageIntLLRInputS0xD(320)(4) <= LUT_4bit_to_3bit(ChLLRxDI(284));
  CNStageIntLLRInputS0xD(353)(4) <= LUT_4bit_to_3bit(ChLLRxDI(284));
  CNStageIntLLRInputS0xD(25)(4) <= LUT_4bit_to_3bit(ChLLRxDI(285));
  CNStageIntLLRInputS0xD(82)(4) <= LUT_4bit_to_3bit(ChLLRxDI(285));
  CNStageIntLLRInputS0xD(165)(4) <= LUT_4bit_to_3bit(ChLLRxDI(285));
  CNStageIntLLRInputS0xD(172)(4) <= LUT_4bit_to_3bit(ChLLRxDI(285));
  CNStageIntLLRInputS0xD(255)(4) <= LUT_4bit_to_3bit(ChLLRxDI(285));
  CNStageIntLLRInputS0xD(304)(4) <= LUT_4bit_to_3bit(ChLLRxDI(285));
  CNStageIntLLRInputS0xD(355)(4) <= LUT_4bit_to_3bit(ChLLRxDI(285));
  CNStageIntLLRInputS0xD(24)(4) <= LUT_4bit_to_3bit(ChLLRxDI(286));
  CNStageIntLLRInputS0xD(93)(4) <= LUT_4bit_to_3bit(ChLLRxDI(286));
  CNStageIntLLRInputS0xD(155)(4) <= LUT_4bit_to_3bit(ChLLRxDI(286));
  CNStageIntLLRInputS0xD(189)(4) <= LUT_4bit_to_3bit(ChLLRxDI(286));
  CNStageIntLLRInputS0xD(267)(4) <= LUT_4bit_to_3bit(ChLLRxDI(286));
  CNStageIntLLRInputS0xD(330)(4) <= LUT_4bit_to_3bit(ChLLRxDI(286));
  CNStageIntLLRInputS0xD(341)(4) <= LUT_4bit_to_3bit(ChLLRxDI(286));
  CNStageIntLLRInputS0xD(23)(4) <= LUT_4bit_to_3bit(ChLLRxDI(287));
  CNStageIntLLRInputS0xD(101)(4) <= LUT_4bit_to_3bit(ChLLRxDI(287));
  CNStageIntLLRInputS0xD(142)(4) <= LUT_4bit_to_3bit(ChLLRxDI(287));
  CNStageIntLLRInputS0xD(193)(4) <= LUT_4bit_to_3bit(ChLLRxDI(287));
  CNStageIntLLRInputS0xD(240)(4) <= LUT_4bit_to_3bit(ChLLRxDI(287));
  CNStageIntLLRInputS0xD(322)(4) <= LUT_4bit_to_3bit(ChLLRxDI(287));
  CNStageIntLLRInputS0xD(375)(4) <= LUT_4bit_to_3bit(ChLLRxDI(287));
  CNStageIntLLRInputS0xD(22)(4) <= LUT_4bit_to_3bit(ChLLRxDI(288));
  CNStageIntLLRInputS0xD(75)(4) <= LUT_4bit_to_3bit(ChLLRxDI(288));
  CNStageIntLLRInputS0xD(161)(4) <= LUT_4bit_to_3bit(ChLLRxDI(288));
  CNStageIntLLRInputS0xD(224)(4) <= LUT_4bit_to_3bit(ChLLRxDI(288));
  CNStageIntLLRInputS0xD(228)(4) <= LUT_4bit_to_3bit(ChLLRxDI(288));
  CNStageIntLLRInputS0xD(308)(4) <= LUT_4bit_to_3bit(ChLLRxDI(288));
  CNStageIntLLRInputS0xD(337)(4) <= LUT_4bit_to_3bit(ChLLRxDI(288));
  CNStageIntLLRInputS0xD(21)(4) <= LUT_4bit_to_3bit(ChLLRxDI(289));
  CNStageIntLLRInputS0xD(89)(4) <= LUT_4bit_to_3bit(ChLLRxDI(289));
  CNStageIntLLRInputS0xD(134)(4) <= LUT_4bit_to_3bit(ChLLRxDI(289));
  CNStageIntLLRInputS0xD(192)(4) <= LUT_4bit_to_3bit(ChLLRxDI(289));
  CNStageIntLLRInputS0xD(269)(4) <= LUT_4bit_to_3bit(ChLLRxDI(289));
  CNStageIntLLRInputS0xD(327)(4) <= LUT_4bit_to_3bit(ChLLRxDI(289));
  CNStageIntLLRInputS0xD(365)(4) <= LUT_4bit_to_3bit(ChLLRxDI(289));
  CNStageIntLLRInputS0xD(20)(4) <= LUT_4bit_to_3bit(ChLLRxDI(290));
  CNStageIntLLRInputS0xD(60)(4) <= LUT_4bit_to_3bit(ChLLRxDI(290));
  CNStageIntLLRInputS0xD(131)(4) <= LUT_4bit_to_3bit(ChLLRxDI(290));
  CNStageIntLLRInputS0xD(187)(4) <= LUT_4bit_to_3bit(ChLLRxDI(290));
  CNStageIntLLRInputS0xD(231)(4) <= LUT_4bit_to_3bit(ChLLRxDI(290));
  CNStageIntLLRInputS0xD(350)(4) <= LUT_4bit_to_3bit(ChLLRxDI(290));
  CNStageIntLLRInputS0xD(19)(4) <= LUT_4bit_to_3bit(ChLLRxDI(291));
  CNStageIntLLRInputS0xD(96)(4) <= LUT_4bit_to_3bit(ChLLRxDI(291));
  CNStageIntLLRInputS0xD(147)(4) <= LUT_4bit_to_3bit(ChLLRxDI(291));
  CNStageIntLLRInputS0xD(223)(4) <= LUT_4bit_to_3bit(ChLLRxDI(291));
  CNStageIntLLRInputS0xD(249)(4) <= LUT_4bit_to_3bit(ChLLRxDI(291));
  CNStageIntLLRInputS0xD(377)(4) <= LUT_4bit_to_3bit(ChLLRxDI(291));
  CNStageIntLLRInputS0xD(18)(4) <= LUT_4bit_to_3bit(ChLLRxDI(292));
  CNStageIntLLRInputS0xD(62)(4) <= LUT_4bit_to_3bit(ChLLRxDI(292));
  CNStageIntLLRInputS0xD(139)(4) <= LUT_4bit_to_3bit(ChLLRxDI(292));
  CNStageIntLLRInputS0xD(177)(4) <= LUT_4bit_to_3bit(ChLLRxDI(292));
  CNStageIntLLRInputS0xD(257)(4) <= LUT_4bit_to_3bit(ChLLRxDI(292));
  CNStageIntLLRInputS0xD(313)(4) <= LUT_4bit_to_3bit(ChLLRxDI(292));
  CNStageIntLLRInputS0xD(367)(4) <= LUT_4bit_to_3bit(ChLLRxDI(292));
  CNStageIntLLRInputS0xD(17)(4) <= LUT_4bit_to_3bit(ChLLRxDI(293));
  CNStageIntLLRInputS0xD(77)(4) <= LUT_4bit_to_3bit(ChLLRxDI(293));
  CNStageIntLLRInputS0xD(113)(4) <= LUT_4bit_to_3bit(ChLLRxDI(293));
  CNStageIntLLRInputS0xD(197)(4) <= LUT_4bit_to_3bit(ChLLRxDI(293));
  CNStageIntLLRInputS0xD(306)(4) <= LUT_4bit_to_3bit(ChLLRxDI(293));
  CNStageIntLLRInputS0xD(354)(4) <= LUT_4bit_to_3bit(ChLLRxDI(293));
  CNStageIntLLRInputS0xD(16)(4) <= LUT_4bit_to_3bit(ChLLRxDI(294));
  CNStageIntLLRInputS0xD(73)(4) <= LUT_4bit_to_3bit(ChLLRxDI(294));
  CNStageIntLLRInputS0xD(123)(4) <= LUT_4bit_to_3bit(ChLLRxDI(294));
  CNStageIntLLRInputS0xD(196)(4) <= LUT_4bit_to_3bit(ChLLRxDI(294));
  CNStageIntLLRInputS0xD(258)(4) <= LUT_4bit_to_3bit(ChLLRxDI(294));
  CNStageIntLLRInputS0xD(284)(4) <= LUT_4bit_to_3bit(ChLLRxDI(294));
  CNStageIntLLRInputS0xD(373)(4) <= LUT_4bit_to_3bit(ChLLRxDI(294));
  CNStageIntLLRInputS0xD(15)(4) <= LUT_4bit_to_3bit(ChLLRxDI(295));
  CNStageIntLLRInputS0xD(92)(4) <= LUT_4bit_to_3bit(ChLLRxDI(295));
  CNStageIntLLRInputS0xD(117)(4) <= LUT_4bit_to_3bit(ChLLRxDI(295));
  CNStageIntLLRInputS0xD(175)(4) <= LUT_4bit_to_3bit(ChLLRxDI(295));
  CNStageIntLLRInputS0xD(346)(4) <= LUT_4bit_to_3bit(ChLLRxDI(295));
  CNStageIntLLRInputS0xD(14)(4) <= LUT_4bit_to_3bit(ChLLRxDI(296));
  CNStageIntLLRInputS0xD(55)(4) <= LUT_4bit_to_3bit(ChLLRxDI(296));
  CNStageIntLLRInputS0xD(121)(4) <= LUT_4bit_to_3bit(ChLLRxDI(296));
  CNStageIntLLRInputS0xD(208)(4) <= LUT_4bit_to_3bit(ChLLRxDI(296));
  CNStageIntLLRInputS0xD(286)(4) <= LUT_4bit_to_3bit(ChLLRxDI(296));
  CNStageIntLLRInputS0xD(343)(4) <= LUT_4bit_to_3bit(ChLLRxDI(296));
  CNStageIntLLRInputS0xD(13)(4) <= LUT_4bit_to_3bit(ChLLRxDI(297));
  CNStageIntLLRInputS0xD(56)(4) <= LUT_4bit_to_3bit(ChLLRxDI(297));
  CNStageIntLLRInputS0xD(111)(4) <= LUT_4bit_to_3bit(ChLLRxDI(297));
  CNStageIntLLRInputS0xD(211)(4) <= LUT_4bit_to_3bit(ChLLRxDI(297));
  CNStageIntLLRInputS0xD(277)(4) <= LUT_4bit_to_3bit(ChLLRxDI(297));
  CNStageIntLLRInputS0xD(290)(4) <= LUT_4bit_to_3bit(ChLLRxDI(297));
  CNStageIntLLRInputS0xD(358)(4) <= LUT_4bit_to_3bit(ChLLRxDI(297));
  CNStageIntLLRInputS0xD(12)(4) <= LUT_4bit_to_3bit(ChLLRxDI(298));
  CNStageIntLLRInputS0xD(91)(4) <= LUT_4bit_to_3bit(ChLLRxDI(298));
  CNStageIntLLRInputS0xD(148)(4) <= LUT_4bit_to_3bit(ChLLRxDI(298));
  CNStageIntLLRInputS0xD(198)(4) <= LUT_4bit_to_3bit(ChLLRxDI(298));
  CNStageIntLLRInputS0xD(262)(4) <= LUT_4bit_to_3bit(ChLLRxDI(298));
  CNStageIntLLRInputS0xD(282)(4) <= LUT_4bit_to_3bit(ChLLRxDI(298));
  CNStageIntLLRInputS0xD(351)(4) <= LUT_4bit_to_3bit(ChLLRxDI(298));
  CNStageIntLLRInputS0xD(83)(4) <= LUT_4bit_to_3bit(ChLLRxDI(299));
  CNStageIntLLRInputS0xD(130)(4) <= LUT_4bit_to_3bit(ChLLRxDI(299));
  CNStageIntLLRInputS0xD(176)(4) <= LUT_4bit_to_3bit(ChLLRxDI(299));
  CNStageIntLLRInputS0xD(264)(4) <= LUT_4bit_to_3bit(ChLLRxDI(299));
  CNStageIntLLRInputS0xD(314)(4) <= LUT_4bit_to_3bit(ChLLRxDI(299));
  CNStageIntLLRInputS0xD(11)(4) <= LUT_4bit_to_3bit(ChLLRxDI(300));
  CNStageIntLLRInputS0xD(99)(4) <= LUT_4bit_to_3bit(ChLLRxDI(300));
  CNStageIntLLRInputS0xD(143)(4) <= LUT_4bit_to_3bit(ChLLRxDI(300));
  CNStageIntLLRInputS0xD(195)(4) <= LUT_4bit_to_3bit(ChLLRxDI(300));
  CNStageIntLLRInputS0xD(299)(4) <= LUT_4bit_to_3bit(ChLLRxDI(300));
  CNStageIntLLRInputS0xD(335)(4) <= LUT_4bit_to_3bit(ChLLRxDI(300));
  CNStageIntLLRInputS0xD(10)(4) <= LUT_4bit_to_3bit(ChLLRxDI(301));
  CNStageIntLLRInputS0xD(103)(4) <= LUT_4bit_to_3bit(ChLLRxDI(301));
  CNStageIntLLRInputS0xD(154)(4) <= LUT_4bit_to_3bit(ChLLRxDI(301));
  CNStageIntLLRInputS0xD(220)(4) <= LUT_4bit_to_3bit(ChLLRxDI(301));
  CNStageIntLLRInputS0xD(270)(4) <= LUT_4bit_to_3bit(ChLLRxDI(301));
  CNStageIntLLRInputS0xD(309)(4) <= LUT_4bit_to_3bit(ChLLRxDI(301));
  CNStageIntLLRInputS0xD(9)(4) <= LUT_4bit_to_3bit(ChLLRxDI(302));
  CNStageIntLLRInputS0xD(110)(4) <= LUT_4bit_to_3bit(ChLLRxDI(302));
  CNStageIntLLRInputS0xD(124)(4) <= LUT_4bit_to_3bit(ChLLRxDI(302));
  CNStageIntLLRInputS0xD(206)(4) <= LUT_4bit_to_3bit(ChLLRxDI(302));
  CNStageIntLLRInputS0xD(227)(4) <= LUT_4bit_to_3bit(ChLLRxDI(302));
  CNStageIntLLRInputS0xD(321)(4) <= LUT_4bit_to_3bit(ChLLRxDI(302));
  CNStageIntLLRInputS0xD(8)(4) <= LUT_4bit_to_3bit(ChLLRxDI(303));
  CNStageIntLLRInputS0xD(102)(4) <= LUT_4bit_to_3bit(ChLLRxDI(303));
  CNStageIntLLRInputS0xD(112)(4) <= LUT_4bit_to_3bit(ChLLRxDI(303));
  CNStageIntLLRInputS0xD(178)(4) <= LUT_4bit_to_3bit(ChLLRxDI(303));
  CNStageIntLLRInputS0xD(235)(4) <= LUT_4bit_to_3bit(ChLLRxDI(303));
  CNStageIntLLRInputS0xD(293)(4) <= LUT_4bit_to_3bit(ChLLRxDI(303));
  CNStageIntLLRInputS0xD(382)(4) <= LUT_4bit_to_3bit(ChLLRxDI(303));
  CNStageIntLLRInputS0xD(7)(4) <= LUT_4bit_to_3bit(ChLLRxDI(304));
  CNStageIntLLRInputS0xD(97)(4) <= LUT_4bit_to_3bit(ChLLRxDI(304));
  CNStageIntLLRInputS0xD(157)(4) <= LUT_4bit_to_3bit(ChLLRxDI(304));
  CNStageIntLLRInputS0xD(222)(4) <= LUT_4bit_to_3bit(ChLLRxDI(304));
  CNStageIntLLRInputS0xD(263)(4) <= LUT_4bit_to_3bit(ChLLRxDI(304));
  CNStageIntLLRInputS0xD(283)(4) <= LUT_4bit_to_3bit(ChLLRxDI(304));
  CNStageIntLLRInputS0xD(359)(4) <= LUT_4bit_to_3bit(ChLLRxDI(304));
  CNStageIntLLRInputS0xD(6)(4) <= LUT_4bit_to_3bit(ChLLRxDI(305));
  CNStageIntLLRInputS0xD(80)(4) <= LUT_4bit_to_3bit(ChLLRxDI(305));
  CNStageIntLLRInputS0xD(115)(4) <= LUT_4bit_to_3bit(ChLLRxDI(305));
  CNStageIntLLRInputS0xD(209)(4) <= LUT_4bit_to_3bit(ChLLRxDI(305));
  CNStageIntLLRInputS0xD(276)(4) <= LUT_4bit_to_3bit(ChLLRxDI(305));
  CNStageIntLLRInputS0xD(323)(4) <= LUT_4bit_to_3bit(ChLLRxDI(305));
  CNStageIntLLRInputS0xD(342)(4) <= LUT_4bit_to_3bit(ChLLRxDI(305));
  CNStageIntLLRInputS0xD(5)(4) <= LUT_4bit_to_3bit(ChLLRxDI(306));
  CNStageIntLLRInputS0xD(87)(4) <= LUT_4bit_to_3bit(ChLLRxDI(306));
  CNStageIntLLRInputS0xD(136)(4) <= LUT_4bit_to_3bit(ChLLRxDI(306));
  CNStageIntLLRInputS0xD(174)(4) <= LUT_4bit_to_3bit(ChLLRxDI(306));
  CNStageIntLLRInputS0xD(4)(4) <= LUT_4bit_to_3bit(ChLLRxDI(307));
  CNStageIntLLRInputS0xD(107)(4) <= LUT_4bit_to_3bit(ChLLRxDI(307));
  CNStageIntLLRInputS0xD(145)(4) <= LUT_4bit_to_3bit(ChLLRxDI(307));
  CNStageIntLLRInputS0xD(202)(4) <= LUT_4bit_to_3bit(ChLLRxDI(307));
  CNStageIntLLRInputS0xD(230)(4) <= LUT_4bit_to_3bit(ChLLRxDI(307));
  CNStageIntLLRInputS0xD(302)(4) <= LUT_4bit_to_3bit(ChLLRxDI(307));
  CNStageIntLLRInputS0xD(366)(4) <= LUT_4bit_to_3bit(ChLLRxDI(307));
  CNStageIntLLRInputS0xD(140)(4) <= LUT_4bit_to_3bit(ChLLRxDI(308));
  CNStageIntLLRInputS0xD(199)(4) <= LUT_4bit_to_3bit(ChLLRxDI(308));
  CNStageIntLLRInputS0xD(251)(4) <= LUT_4bit_to_3bit(ChLLRxDI(308));
  CNStageIntLLRInputS0xD(311)(4) <= LUT_4bit_to_3bit(ChLLRxDI(308));
  CNStageIntLLRInputS0xD(336)(4) <= LUT_4bit_to_3bit(ChLLRxDI(308));
  CNStageIntLLRInputS0xD(3)(4) <= LUT_4bit_to_3bit(ChLLRxDI(309));
  CNStageIntLLRInputS0xD(86)(4) <= LUT_4bit_to_3bit(ChLLRxDI(309));
  CNStageIntLLRInputS0xD(146)(4) <= LUT_4bit_to_3bit(ChLLRxDI(309));
  CNStageIntLLRInputS0xD(214)(4) <= LUT_4bit_to_3bit(ChLLRxDI(309));
  CNStageIntLLRInputS0xD(265)(4) <= LUT_4bit_to_3bit(ChLLRxDI(309));
  CNStageIntLLRInputS0xD(307)(4) <= LUT_4bit_to_3bit(ChLLRxDI(309));
  CNStageIntLLRInputS0xD(2)(4) <= LUT_4bit_to_3bit(ChLLRxDI(310));
  CNStageIntLLRInputS0xD(65)(4) <= LUT_4bit_to_3bit(ChLLRxDI(310));
  CNStageIntLLRInputS0xD(135)(4) <= LUT_4bit_to_3bit(ChLLRxDI(310));
  CNStageIntLLRInputS0xD(261)(4) <= LUT_4bit_to_3bit(ChLLRxDI(310));
  CNStageIntLLRInputS0xD(312)(4) <= LUT_4bit_to_3bit(ChLLRxDI(310));
  CNStageIntLLRInputS0xD(369)(4) <= LUT_4bit_to_3bit(ChLLRxDI(310));
  CNStageIntLLRInputS0xD(1)(4) <= LUT_4bit_to_3bit(ChLLRxDI(311));
  CNStageIntLLRInputS0xD(68)(4) <= LUT_4bit_to_3bit(ChLLRxDI(311));
  CNStageIntLLRInputS0xD(160)(4) <= LUT_4bit_to_3bit(ChLLRxDI(311));
  CNStageIntLLRInputS0xD(225)(4) <= LUT_4bit_to_3bit(ChLLRxDI(311));
  CNStageIntLLRInputS0xD(301)(4) <= LUT_4bit_to_3bit(ChLLRxDI(311));
  CNStageIntLLRInputS0xD(0)(4) <= LUT_4bit_to_3bit(ChLLRxDI(312));
  CNStageIntLLRInputS0xD(108)(4) <= LUT_4bit_to_3bit(ChLLRxDI(312));
  CNStageIntLLRInputS0xD(167)(4) <= LUT_4bit_to_3bit(ChLLRxDI(312));
  CNStageIntLLRInputS0xD(246)(4) <= LUT_4bit_to_3bit(ChLLRxDI(312));
  CNStageIntLLRInputS0xD(326)(4) <= LUT_4bit_to_3bit(ChLLRxDI(312));
  CNStageIntLLRInputS0xD(348)(4) <= LUT_4bit_to_3bit(ChLLRxDI(312));
  CNStageIntLLRInputS0xD(150)(4) <= LUT_4bit_to_3bit(ChLLRxDI(313));
  CNStageIntLLRInputS0xD(188)(4) <= LUT_4bit_to_3bit(ChLLRxDI(313));
  CNStageIntLLRInputS0xD(247)(4) <= LUT_4bit_to_3bit(ChLLRxDI(313));
  CNStageIntLLRInputS0xD(356)(4) <= LUT_4bit_to_3bit(ChLLRxDI(313));
  CNStageIntLLRInputS0xD(191)(4) <= LUT_4bit_to_3bit(ChLLRxDI(314));
  CNStageIntLLRInputS0xD(278)(4) <= LUT_4bit_to_3bit(ChLLRxDI(314));
  CNStageIntLLRInputS0xD(316)(4) <= LUT_4bit_to_3bit(ChLLRxDI(314));
  CNStageIntLLRInputS0xD(352)(4) <= LUT_4bit_to_3bit(ChLLRxDI(314));
  CNStageIntLLRInputS0xD(78)(4) <= LUT_4bit_to_3bit(ChLLRxDI(315));
  CNStageIntLLRInputS0xD(119)(4) <= LUT_4bit_to_3bit(ChLLRxDI(315));
  CNStageIntLLRInputS0xD(183)(4) <= LUT_4bit_to_3bit(ChLLRxDI(315));
  CNStageIntLLRInputS0xD(271)(4) <= LUT_4bit_to_3bit(ChLLRxDI(315));
  CNStageIntLLRInputS0xD(318)(4) <= LUT_4bit_to_3bit(ChLLRxDI(315));
  CNStageIntLLRInputS0xD(357)(4) <= LUT_4bit_to_3bit(ChLLRxDI(315));
  CNStageIntLLRInputS0xD(61)(4) <= LUT_4bit_to_3bit(ChLLRxDI(316));
  CNStageIntLLRInputS0xD(158)(4) <= LUT_4bit_to_3bit(ChLLRxDI(316));
  CNStageIntLLRInputS0xD(234)(4) <= LUT_4bit_to_3bit(ChLLRxDI(316));
  CNStageIntLLRInputS0xD(288)(4) <= LUT_4bit_to_3bit(ChLLRxDI(316));
  CNStageIntLLRInputS0xD(347)(4) <= LUT_4bit_to_3bit(ChLLRxDI(316));
  CNStageIntLLRInputS0xD(88)(4) <= LUT_4bit_to_3bit(ChLLRxDI(317));
  CNStageIntLLRInputS0xD(238)(4) <= LUT_4bit_to_3bit(ChLLRxDI(317));
  CNStageIntLLRInputS0xD(324)(4) <= LUT_4bit_to_3bit(ChLLRxDI(317));
  CNStageIntLLRInputS0xD(372)(4) <= LUT_4bit_to_3bit(ChLLRxDI(317));
  CNStageIntLLRInputS0xD(120)(4) <= LUT_4bit_to_3bit(ChLLRxDI(318));
  CNStageIntLLRInputS0xD(210)(4) <= LUT_4bit_to_3bit(ChLLRxDI(318));
  CNStageIntLLRInputS0xD(279)(4) <= LUT_4bit_to_3bit(ChLLRxDI(318));
  CNStageIntLLRInputS0xD(379)(4) <= LUT_4bit_to_3bit(ChLLRxDI(318));
  CNStageIntLLRInputS0xD(52)(4) <= LUT_4bit_to_3bit(ChLLRxDI(319));
  CNStageIntLLRInputS0xD(66)(4) <= LUT_4bit_to_3bit(ChLLRxDI(319));
  CNStageIntLLRInputS0xD(151)(4) <= LUT_4bit_to_3bit(ChLLRxDI(319));
  CNStageIntLLRInputS0xD(221)(4) <= LUT_4bit_to_3bit(ChLLRxDI(319));
  CNStageIntLLRInputS0xD(237)(4) <= LUT_4bit_to_3bit(ChLLRxDI(319));
  CNStageIntLLRInputS0xD(289)(4) <= LUT_4bit_to_3bit(ChLLRxDI(319));
  CNStageIntLLRInputS0xD(361)(4) <= LUT_4bit_to_3bit(ChLLRxDI(319));
  CNStageIntLLRInputS0xD(53)(5) <= LUT_4bit_to_3bit(ChLLRxDI(320));
  CNStageIntLLRInputS0xD(126)(5) <= LUT_4bit_to_3bit(ChLLRxDI(320));
  CNStageIntLLRInputS0xD(196)(5) <= LUT_4bit_to_3bit(ChLLRxDI(320));
  CNStageIntLLRInputS0xD(295)(5) <= LUT_4bit_to_3bit(ChLLRxDI(320));
  CNStageIntLLRInputS0xD(338)(5) <= LUT_4bit_to_3bit(ChLLRxDI(320));
  CNStageIntLLRInputS0xD(51)(5) <= LUT_4bit_to_3bit(ChLLRxDI(321));
  CNStageIntLLRInputS0xD(65)(5) <= LUT_4bit_to_3bit(ChLLRxDI(321));
  CNStageIntLLRInputS0xD(150)(5) <= LUT_4bit_to_3bit(ChLLRxDI(321));
  CNStageIntLLRInputS0xD(220)(5) <= LUT_4bit_to_3bit(ChLLRxDI(321));
  CNStageIntLLRInputS0xD(236)(5) <= LUT_4bit_to_3bit(ChLLRxDI(321));
  CNStageIntLLRInputS0xD(288)(5) <= LUT_4bit_to_3bit(ChLLRxDI(321));
  CNStageIntLLRInputS0xD(360)(5) <= LUT_4bit_to_3bit(ChLLRxDI(321));
  CNStageIntLLRInputS0xD(50)(5) <= LUT_4bit_to_3bit(ChLLRxDI(322));
  CNStageIntLLRInputS0xD(84)(5) <= LUT_4bit_to_3bit(ChLLRxDI(322));
  CNStageIntLLRInputS0xD(165)(5) <= LUT_4bit_to_3bit(ChLLRxDI(322));
  CNStageIntLLRInputS0xD(231)(5) <= LUT_4bit_to_3bit(ChLLRxDI(322));
  CNStageIntLLRInputS0xD(316)(5) <= LUT_4bit_to_3bit(ChLLRxDI(322));
  CNStageIntLLRInputS0xD(362)(5) <= LUT_4bit_to_3bit(ChLLRxDI(322));
  CNStageIntLLRInputS0xD(56)(5) <= LUT_4bit_to_3bit(ChLLRxDI(323));
  CNStageIntLLRInputS0xD(136)(5) <= LUT_4bit_to_3bit(ChLLRxDI(323));
  CNStageIntLLRInputS0xD(184)(5) <= LUT_4bit_to_3bit(ChLLRxDI(323));
  CNStageIntLLRInputS0xD(268)(5) <= LUT_4bit_to_3bit(ChLLRxDI(323));
  CNStageIntLLRInputS0xD(330)(5) <= LUT_4bit_to_3bit(ChLLRxDI(323));
  CNStageIntLLRInputS0xD(49)(5) <= LUT_4bit_to_3bit(ChLLRxDI(324));
  CNStageIntLLRInputS0xD(109)(5) <= LUT_4bit_to_3bit(ChLLRxDI(324));
  CNStageIntLLRInputS0xD(113)(5) <= LUT_4bit_to_3bit(ChLLRxDI(324));
  CNStageIntLLRInputS0xD(223)(5) <= LUT_4bit_to_3bit(ChLLRxDI(324));
  CNStageIntLLRInputS0xD(273)(5) <= LUT_4bit_to_3bit(ChLLRxDI(324));
  CNStageIntLLRInputS0xD(302)(5) <= LUT_4bit_to_3bit(ChLLRxDI(324));
  CNStageIntLLRInputS0xD(369)(5) <= LUT_4bit_to_3bit(ChLLRxDI(324));
  CNStageIntLLRInputS0xD(48)(5) <= LUT_4bit_to_3bit(ChLLRxDI(325));
  CNStageIntLLRInputS0xD(70)(5) <= LUT_4bit_to_3bit(ChLLRxDI(325));
  CNStageIntLLRInputS0xD(137)(5) <= LUT_4bit_to_3bit(ChLLRxDI(325));
  CNStageIntLLRInputS0xD(185)(5) <= LUT_4bit_to_3bit(ChLLRxDI(325));
  CNStageIntLLRInputS0xD(242)(5) <= LUT_4bit_to_3bit(ChLLRxDI(325));
  CNStageIntLLRInputS0xD(284)(5) <= LUT_4bit_to_3bit(ChLLRxDI(325));
  CNStageIntLLRInputS0xD(382)(5) <= LUT_4bit_to_3bit(ChLLRxDI(325));
  CNStageIntLLRInputS0xD(47)(5) <= LUT_4bit_to_3bit(ChLLRxDI(326));
  CNStageIntLLRInputS0xD(62)(5) <= LUT_4bit_to_3bit(ChLLRxDI(326));
  CNStageIntLLRInputS0xD(203)(5) <= LUT_4bit_to_3bit(ChLLRxDI(326));
  CNStageIntLLRInputS0xD(241)(5) <= LUT_4bit_to_3bit(ChLLRxDI(326));
  CNStageIntLLRInputS0xD(304)(5) <= LUT_4bit_to_3bit(ChLLRxDI(326));
  CNStageIntLLRInputS0xD(46)(5) <= LUT_4bit_to_3bit(ChLLRxDI(327));
  CNStageIntLLRInputS0xD(94)(5) <= LUT_4bit_to_3bit(ChLLRxDI(327));
  CNStageIntLLRInputS0xD(148)(5) <= LUT_4bit_to_3bit(ChLLRxDI(327));
  CNStageIntLLRInputS0xD(211)(5) <= LUT_4bit_to_3bit(ChLLRxDI(327));
  CNStageIntLLRInputS0xD(272)(5) <= LUT_4bit_to_3bit(ChLLRxDI(327));
  CNStageIntLLRInputS0xD(318)(5) <= LUT_4bit_to_3bit(ChLLRxDI(327));
  CNStageIntLLRInputS0xD(361)(5) <= LUT_4bit_to_3bit(ChLLRxDI(327));
  CNStageIntLLRInputS0xD(45)(5) <= LUT_4bit_to_3bit(ChLLRxDI(328));
  CNStageIntLLRInputS0xD(103)(5) <= LUT_4bit_to_3bit(ChLLRxDI(328));
  CNStageIntLLRInputS0xD(168)(5) <= LUT_4bit_to_3bit(ChLLRxDI(328));
  CNStageIntLLRInputS0xD(314)(5) <= LUT_4bit_to_3bit(ChLLRxDI(328));
  CNStageIntLLRInputS0xD(377)(5) <= LUT_4bit_to_3bit(ChLLRxDI(328));
  CNStageIntLLRInputS0xD(44)(5) <= LUT_4bit_to_3bit(ChLLRxDI(329));
  CNStageIntLLRInputS0xD(97)(5) <= LUT_4bit_to_3bit(ChLLRxDI(329));
  CNStageIntLLRInputS0xD(131)(5) <= LUT_4bit_to_3bit(ChLLRxDI(329));
  CNStageIntLLRInputS0xD(212)(5) <= LUT_4bit_to_3bit(ChLLRxDI(329));
  CNStageIntLLRInputS0xD(255)(5) <= LUT_4bit_to_3bit(ChLLRxDI(329));
  CNStageIntLLRInputS0xD(280)(5) <= LUT_4bit_to_3bit(ChLLRxDI(329));
  CNStageIntLLRInputS0xD(348)(5) <= LUT_4bit_to_3bit(ChLLRxDI(329));
  CNStageIntLLRInputS0xD(43)(5) <= LUT_4bit_to_3bit(ChLLRxDI(330));
  CNStageIntLLRInputS0xD(101)(5) <= LUT_4bit_to_3bit(ChLLRxDI(330));
  CNStageIntLLRInputS0xD(132)(5) <= LUT_4bit_to_3bit(ChLLRxDI(330));
  CNStageIntLLRInputS0xD(202)(5) <= LUT_4bit_to_3bit(ChLLRxDI(330));
  CNStageIntLLRInputS0xD(243)(5) <= LUT_4bit_to_3bit(ChLLRxDI(330));
  CNStageIntLLRInputS0xD(42)(5) <= LUT_4bit_to_3bit(ChLLRxDI(331));
  CNStageIntLLRInputS0xD(92)(5) <= LUT_4bit_to_3bit(ChLLRxDI(331));
  CNStageIntLLRInputS0xD(167)(5) <= LUT_4bit_to_3bit(ChLLRxDI(331));
  CNStageIntLLRInputS0xD(172)(5) <= LUT_4bit_to_3bit(ChLLRxDI(331));
  CNStageIntLLRInputS0xD(350)(5) <= LUT_4bit_to_3bit(ChLLRxDI(331));
  CNStageIntLLRInputS0xD(41)(5) <= LUT_4bit_to_3bit(ChLLRxDI(332));
  CNStageIntLLRInputS0xD(71)(5) <= LUT_4bit_to_3bit(ChLLRxDI(332));
  CNStageIntLLRInputS0xD(158)(5) <= LUT_4bit_to_3bit(ChLLRxDI(332));
  CNStageIntLLRInputS0xD(179)(5) <= LUT_4bit_to_3bit(ChLLRxDI(332));
  CNStageIntLLRInputS0xD(240)(5) <= LUT_4bit_to_3bit(ChLLRxDI(332));
  CNStageIntLLRInputS0xD(363)(5) <= LUT_4bit_to_3bit(ChLLRxDI(332));
  CNStageIntLLRInputS0xD(108)(5) <= LUT_4bit_to_3bit(ChLLRxDI(333));
  CNStageIntLLRInputS0xD(117)(5) <= LUT_4bit_to_3bit(ChLLRxDI(333));
  CNStageIntLLRInputS0xD(215)(5) <= LUT_4bit_to_3bit(ChLLRxDI(333));
  CNStageIntLLRInputS0xD(265)(5) <= LUT_4bit_to_3bit(ChLLRxDI(333));
  CNStageIntLLRInputS0xD(324)(5) <= LUT_4bit_to_3bit(ChLLRxDI(333));
  CNStageIntLLRInputS0xD(359)(5) <= LUT_4bit_to_3bit(ChLLRxDI(333));
  CNStageIntLLRInputS0xD(40)(5) <= LUT_4bit_to_3bit(ChLLRxDI(334));
  CNStageIntLLRInputS0xD(66)(5) <= LUT_4bit_to_3bit(ChLLRxDI(334));
  CNStageIntLLRInputS0xD(217)(5) <= LUT_4bit_to_3bit(ChLLRxDI(334));
  CNStageIntLLRInputS0xD(286)(5) <= LUT_4bit_to_3bit(ChLLRxDI(334));
  CNStageIntLLRInputS0xD(380)(5) <= LUT_4bit_to_3bit(ChLLRxDI(334));
  CNStageIntLLRInputS0xD(39)(5) <= LUT_4bit_to_3bit(ChLLRxDI(335));
  CNStageIntLLRInputS0xD(78)(5) <= LUT_4bit_to_3bit(ChLLRxDI(335));
  CNStageIntLLRInputS0xD(170)(5) <= LUT_4bit_to_3bit(ChLLRxDI(335));
  CNStageIntLLRInputS0xD(189)(5) <= LUT_4bit_to_3bit(ChLLRxDI(335));
  CNStageIntLLRInputS0xD(274)(5) <= LUT_4bit_to_3bit(ChLLRxDI(335));
  CNStageIntLLRInputS0xD(291)(5) <= LUT_4bit_to_3bit(ChLLRxDI(335));
  CNStageIntLLRInputS0xD(343)(5) <= LUT_4bit_to_3bit(ChLLRxDI(335));
  CNStageIntLLRInputS0xD(38)(5) <= LUT_4bit_to_3bit(ChLLRxDI(336));
  CNStageIntLLRInputS0xD(104)(5) <= LUT_4bit_to_3bit(ChLLRxDI(336));
  CNStageIntLLRInputS0xD(121)(5) <= LUT_4bit_to_3bit(ChLLRxDI(336));
  CNStageIntLLRInputS0xD(267)(5) <= LUT_4bit_to_3bit(ChLLRxDI(336));
  CNStageIntLLRInputS0xD(332)(5) <= LUT_4bit_to_3bit(ChLLRxDI(336));
  CNStageIntLLRInputS0xD(344)(5) <= LUT_4bit_to_3bit(ChLLRxDI(336));
  CNStageIntLLRInputS0xD(37)(5) <= LUT_4bit_to_3bit(ChLLRxDI(337));
  CNStageIntLLRInputS0xD(93)(5) <= LUT_4bit_to_3bit(ChLLRxDI(337));
  CNStageIntLLRInputS0xD(115)(5) <= LUT_4bit_to_3bit(ChLLRxDI(337));
  CNStageIntLLRInputS0xD(183)(5) <= LUT_4bit_to_3bit(ChLLRxDI(337));
  CNStageIntLLRInputS0xD(253)(5) <= LUT_4bit_to_3bit(ChLLRxDI(337));
  CNStageIntLLRInputS0xD(290)(5) <= LUT_4bit_to_3bit(ChLLRxDI(337));
  CNStageIntLLRInputS0xD(379)(5) <= LUT_4bit_to_3bit(ChLLRxDI(337));
  CNStageIntLLRInputS0xD(36)(5) <= LUT_4bit_to_3bit(ChLLRxDI(338));
  CNStageIntLLRInputS0xD(80)(5) <= LUT_4bit_to_3bit(ChLLRxDI(338));
  CNStageIntLLRInputS0xD(155)(5) <= LUT_4bit_to_3bit(ChLLRxDI(338));
  CNStageIntLLRInputS0xD(190)(5) <= LUT_4bit_to_3bit(ChLLRxDI(338));
  CNStageIntLLRInputS0xD(370)(5) <= LUT_4bit_to_3bit(ChLLRxDI(338));
  CNStageIntLLRInputS0xD(35)(5) <= LUT_4bit_to_3bit(ChLLRxDI(339));
  CNStageIntLLRInputS0xD(96)(5) <= LUT_4bit_to_3bit(ChLLRxDI(339));
  CNStageIntLLRInputS0xD(163)(5) <= LUT_4bit_to_3bit(ChLLRxDI(339));
  CNStageIntLLRInputS0xD(216)(5) <= LUT_4bit_to_3bit(ChLLRxDI(339));
  CNStageIntLLRInputS0xD(247)(5) <= LUT_4bit_to_3bit(ChLLRxDI(339));
  CNStageIntLLRInputS0xD(322)(5) <= LUT_4bit_to_3bit(ChLLRxDI(339));
  CNStageIntLLRInputS0xD(34)(5) <= LUT_4bit_to_3bit(ChLLRxDI(340));
  CNStageIntLLRInputS0xD(58)(5) <= LUT_4bit_to_3bit(ChLLRxDI(340));
  CNStageIntLLRInputS0xD(127)(5) <= LUT_4bit_to_3bit(ChLLRxDI(340));
  CNStageIntLLRInputS0xD(178)(5) <= LUT_4bit_to_3bit(ChLLRxDI(340));
  CNStageIntLLRInputS0xD(245)(5) <= LUT_4bit_to_3bit(ChLLRxDI(340));
  CNStageIntLLRInputS0xD(334)(5) <= LUT_4bit_to_3bit(ChLLRxDI(340));
  CNStageIntLLRInputS0xD(33)(5) <= LUT_4bit_to_3bit(ChLLRxDI(341));
  CNStageIntLLRInputS0xD(68)(5) <= LUT_4bit_to_3bit(ChLLRxDI(341));
  CNStageIntLLRInputS0xD(125)(5) <= LUT_4bit_to_3bit(ChLLRxDI(341));
  CNStageIntLLRInputS0xD(204)(5) <= LUT_4bit_to_3bit(ChLLRxDI(341));
  CNStageIntLLRInputS0xD(258)(5) <= LUT_4bit_to_3bit(ChLLRxDI(341));
  CNStageIntLLRInputS0xD(296)(5) <= LUT_4bit_to_3bit(ChLLRxDI(341));
  CNStageIntLLRInputS0xD(32)(5) <= LUT_4bit_to_3bit(ChLLRxDI(342));
  CNStageIntLLRInputS0xD(63)(5) <= LUT_4bit_to_3bit(ChLLRxDI(342));
  CNStageIntLLRInputS0xD(161)(5) <= LUT_4bit_to_3bit(ChLLRxDI(342));
  CNStageIntLLRInputS0xD(251)(5) <= LUT_4bit_to_3bit(ChLLRxDI(342));
  CNStageIntLLRInputS0xD(294)(5) <= LUT_4bit_to_3bit(ChLLRxDI(342));
  CNStageIntLLRInputS0xD(31)(5) <= LUT_4bit_to_3bit(ChLLRxDI(343));
  CNStageIntLLRInputS0xD(69)(5) <= LUT_4bit_to_3bit(ChLLRxDI(343));
  CNStageIntLLRInputS0xD(140)(5) <= LUT_4bit_to_3bit(ChLLRxDI(343));
  CNStageIntLLRInputS0xD(206)(5) <= LUT_4bit_to_3bit(ChLLRxDI(343));
  CNStageIntLLRInputS0xD(228)(5) <= LUT_4bit_to_3bit(ChLLRxDI(343));
  CNStageIntLLRInputS0xD(327)(5) <= LUT_4bit_to_3bit(ChLLRxDI(343));
  CNStageIntLLRInputS0xD(30)(5) <= LUT_4bit_to_3bit(ChLLRxDI(344));
  CNStageIntLLRInputS0xD(57)(5) <= LUT_4bit_to_3bit(ChLLRxDI(344));
  CNStageIntLLRInputS0xD(143)(5) <= LUT_4bit_to_3bit(ChLLRxDI(344));
  CNStageIntLLRInputS0xD(218)(5) <= LUT_4bit_to_3bit(ChLLRxDI(344));
  CNStageIntLLRInputS0xD(238)(5) <= LUT_4bit_to_3bit(ChLLRxDI(344));
  CNStageIntLLRInputS0xD(307)(5) <= LUT_4bit_to_3bit(ChLLRxDI(344));
  CNStageIntLLRInputS0xD(367)(5) <= LUT_4bit_to_3bit(ChLLRxDI(344));
  CNStageIntLLRInputS0xD(29)(5) <= LUT_4bit_to_3bit(ChLLRxDI(345));
  CNStageIntLLRInputS0xD(83)(5) <= LUT_4bit_to_3bit(ChLLRxDI(345));
  CNStageIntLLRInputS0xD(128)(5) <= LUT_4bit_to_3bit(ChLLRxDI(345));
  CNStageIntLLRInputS0xD(232)(5) <= LUT_4bit_to_3bit(ChLLRxDI(345));
  CNStageIntLLRInputS0xD(309)(5) <= LUT_4bit_to_3bit(ChLLRxDI(345));
  CNStageIntLLRInputS0xD(375)(5) <= LUT_4bit_to_3bit(ChLLRxDI(345));
  CNStageIntLLRInputS0xD(28)(5) <= LUT_4bit_to_3bit(ChLLRxDI(346));
  CNStageIntLLRInputS0xD(89)(5) <= LUT_4bit_to_3bit(ChLLRxDI(346));
  CNStageIntLLRInputS0xD(162)(5) <= LUT_4bit_to_3bit(ChLLRxDI(346));
  CNStageIntLLRInputS0xD(181)(5) <= LUT_4bit_to_3bit(ChLLRxDI(346));
  CNStageIntLLRInputS0xD(235)(5) <= LUT_4bit_to_3bit(ChLLRxDI(346));
  CNStageIntLLRInputS0xD(297)(5) <= LUT_4bit_to_3bit(ChLLRxDI(346));
  CNStageIntLLRInputS0xD(339)(5) <= LUT_4bit_to_3bit(ChLLRxDI(346));
  CNStageIntLLRInputS0xD(27)(5) <= LUT_4bit_to_3bit(ChLLRxDI(347));
  CNStageIntLLRInputS0xD(73)(5) <= LUT_4bit_to_3bit(ChLLRxDI(347));
  CNStageIntLLRInputS0xD(124)(5) <= LUT_4bit_to_3bit(ChLLRxDI(347));
  CNStageIntLLRInputS0xD(199)(5) <= LUT_4bit_to_3bit(ChLLRxDI(347));
  CNStageIntLLRInputS0xD(225)(5) <= LUT_4bit_to_3bit(ChLLRxDI(347));
  CNStageIntLLRInputS0xD(328)(5) <= LUT_4bit_to_3bit(ChLLRxDI(347));
  CNStageIntLLRInputS0xD(337)(5) <= LUT_4bit_to_3bit(ChLLRxDI(347));
  CNStageIntLLRInputS0xD(26)(5) <= LUT_4bit_to_3bit(ChLLRxDI(348));
  CNStageIntLLRInputS0xD(75)(5) <= LUT_4bit_to_3bit(ChLLRxDI(348));
  CNStageIntLLRInputS0xD(152)(5) <= LUT_4bit_to_3bit(ChLLRxDI(348));
  CNStageIntLLRInputS0xD(200)(5) <= LUT_4bit_to_3bit(ChLLRxDI(348));
  CNStageIntLLRInputS0xD(259)(5) <= LUT_4bit_to_3bit(ChLLRxDI(348));
  CNStageIntLLRInputS0xD(293)(5) <= LUT_4bit_to_3bit(ChLLRxDI(348));
  CNStageIntLLRInputS0xD(373)(5) <= LUT_4bit_to_3bit(ChLLRxDI(348));
  CNStageIntLLRInputS0xD(25)(5) <= LUT_4bit_to_3bit(ChLLRxDI(349));
  CNStageIntLLRInputS0xD(99)(5) <= LUT_4bit_to_3bit(ChLLRxDI(349));
  CNStageIntLLRInputS0xD(180)(5) <= LUT_4bit_to_3bit(ChLLRxDI(349));
  CNStageIntLLRInputS0xD(244)(5) <= LUT_4bit_to_3bit(ChLLRxDI(349));
  CNStageIntLLRInputS0xD(319)(5) <= LUT_4bit_to_3bit(ChLLRxDI(349));
  CNStageIntLLRInputS0xD(352)(5) <= LUT_4bit_to_3bit(ChLLRxDI(349));
  CNStageIntLLRInputS0xD(24)(5) <= LUT_4bit_to_3bit(ChLLRxDI(350));
  CNStageIntLLRInputS0xD(81)(5) <= LUT_4bit_to_3bit(ChLLRxDI(350));
  CNStageIntLLRInputS0xD(164)(5) <= LUT_4bit_to_3bit(ChLLRxDI(350));
  CNStageIntLLRInputS0xD(171)(5) <= LUT_4bit_to_3bit(ChLLRxDI(350));
  CNStageIntLLRInputS0xD(254)(5) <= LUT_4bit_to_3bit(ChLLRxDI(350));
  CNStageIntLLRInputS0xD(303)(5) <= LUT_4bit_to_3bit(ChLLRxDI(350));
  CNStageIntLLRInputS0xD(23)(5) <= LUT_4bit_to_3bit(ChLLRxDI(351));
  CNStageIntLLRInputS0xD(154)(5) <= LUT_4bit_to_3bit(ChLLRxDI(351));
  CNStageIntLLRInputS0xD(188)(5) <= LUT_4bit_to_3bit(ChLLRxDI(351));
  CNStageIntLLRInputS0xD(266)(5) <= LUT_4bit_to_3bit(ChLLRxDI(351));
  CNStageIntLLRInputS0xD(329)(5) <= LUT_4bit_to_3bit(ChLLRxDI(351));
  CNStageIntLLRInputS0xD(340)(5) <= LUT_4bit_to_3bit(ChLLRxDI(351));
  CNStageIntLLRInputS0xD(22)(5) <= LUT_4bit_to_3bit(ChLLRxDI(352));
  CNStageIntLLRInputS0xD(100)(5) <= LUT_4bit_to_3bit(ChLLRxDI(352));
  CNStageIntLLRInputS0xD(141)(5) <= LUT_4bit_to_3bit(ChLLRxDI(352));
  CNStageIntLLRInputS0xD(192)(5) <= LUT_4bit_to_3bit(ChLLRxDI(352));
  CNStageIntLLRInputS0xD(239)(5) <= LUT_4bit_to_3bit(ChLLRxDI(352));
  CNStageIntLLRInputS0xD(321)(5) <= LUT_4bit_to_3bit(ChLLRxDI(352));
  CNStageIntLLRInputS0xD(374)(5) <= LUT_4bit_to_3bit(ChLLRxDI(352));
  CNStageIntLLRInputS0xD(21)(5) <= LUT_4bit_to_3bit(ChLLRxDI(353));
  CNStageIntLLRInputS0xD(74)(5) <= LUT_4bit_to_3bit(ChLLRxDI(353));
  CNStageIntLLRInputS0xD(160)(5) <= LUT_4bit_to_3bit(ChLLRxDI(353));
  CNStageIntLLRInputS0xD(224)(5) <= LUT_4bit_to_3bit(ChLLRxDI(353));
  CNStageIntLLRInputS0xD(227)(5) <= LUT_4bit_to_3bit(ChLLRxDI(353));
  CNStageIntLLRInputS0xD(336)(5) <= LUT_4bit_to_3bit(ChLLRxDI(353));
  CNStageIntLLRInputS0xD(20)(5) <= LUT_4bit_to_3bit(ChLLRxDI(354));
  CNStageIntLLRInputS0xD(88)(5) <= LUT_4bit_to_3bit(ChLLRxDI(354));
  CNStageIntLLRInputS0xD(133)(5) <= LUT_4bit_to_3bit(ChLLRxDI(354));
  CNStageIntLLRInputS0xD(191)(5) <= LUT_4bit_to_3bit(ChLLRxDI(354));
  CNStageIntLLRInputS0xD(326)(5) <= LUT_4bit_to_3bit(ChLLRxDI(354));
  CNStageIntLLRInputS0xD(364)(5) <= LUT_4bit_to_3bit(ChLLRxDI(354));
  CNStageIntLLRInputS0xD(19)(5) <= LUT_4bit_to_3bit(ChLLRxDI(355));
  CNStageIntLLRInputS0xD(59)(5) <= LUT_4bit_to_3bit(ChLLRxDI(355));
  CNStageIntLLRInputS0xD(130)(5) <= LUT_4bit_to_3bit(ChLLRxDI(355));
  CNStageIntLLRInputS0xD(186)(5) <= LUT_4bit_to_3bit(ChLLRxDI(355));
  CNStageIntLLRInputS0xD(230)(5) <= LUT_4bit_to_3bit(ChLLRxDI(355));
  CNStageIntLLRInputS0xD(300)(5) <= LUT_4bit_to_3bit(ChLLRxDI(355));
  CNStageIntLLRInputS0xD(349)(5) <= LUT_4bit_to_3bit(ChLLRxDI(355));
  CNStageIntLLRInputS0xD(18)(5) <= LUT_4bit_to_3bit(ChLLRxDI(356));
  CNStageIntLLRInputS0xD(95)(5) <= LUT_4bit_to_3bit(ChLLRxDI(356));
  CNStageIntLLRInputS0xD(146)(5) <= LUT_4bit_to_3bit(ChLLRxDI(356));
  CNStageIntLLRInputS0xD(222)(5) <= LUT_4bit_to_3bit(ChLLRxDI(356));
  CNStageIntLLRInputS0xD(299)(5) <= LUT_4bit_to_3bit(ChLLRxDI(356));
  CNStageIntLLRInputS0xD(376)(5) <= LUT_4bit_to_3bit(ChLLRxDI(356));
  CNStageIntLLRInputS0xD(17)(5) <= LUT_4bit_to_3bit(ChLLRxDI(357));
  CNStageIntLLRInputS0xD(61)(5) <= LUT_4bit_to_3bit(ChLLRxDI(357));
  CNStageIntLLRInputS0xD(138)(5) <= LUT_4bit_to_3bit(ChLLRxDI(357));
  CNStageIntLLRInputS0xD(176)(5) <= LUT_4bit_to_3bit(ChLLRxDI(357));
  CNStageIntLLRInputS0xD(256)(5) <= LUT_4bit_to_3bit(ChLLRxDI(357));
  CNStageIntLLRInputS0xD(312)(5) <= LUT_4bit_to_3bit(ChLLRxDI(357));
  CNStageIntLLRInputS0xD(366)(5) <= LUT_4bit_to_3bit(ChLLRxDI(357));
  CNStageIntLLRInputS0xD(16)(5) <= LUT_4bit_to_3bit(ChLLRxDI(358));
  CNStageIntLLRInputS0xD(76)(5) <= LUT_4bit_to_3bit(ChLLRxDI(358));
  CNStageIntLLRInputS0xD(112)(5) <= LUT_4bit_to_3bit(ChLLRxDI(358));
  CNStageIntLLRInputS0xD(252)(5) <= LUT_4bit_to_3bit(ChLLRxDI(358));
  CNStageIntLLRInputS0xD(305)(5) <= LUT_4bit_to_3bit(ChLLRxDI(358));
  CNStageIntLLRInputS0xD(353)(5) <= LUT_4bit_to_3bit(ChLLRxDI(358));
  CNStageIntLLRInputS0xD(15)(5) <= LUT_4bit_to_3bit(ChLLRxDI(359));
  CNStageIntLLRInputS0xD(72)(5) <= LUT_4bit_to_3bit(ChLLRxDI(359));
  CNStageIntLLRInputS0xD(122)(5) <= LUT_4bit_to_3bit(ChLLRxDI(359));
  CNStageIntLLRInputS0xD(195)(5) <= LUT_4bit_to_3bit(ChLLRxDI(359));
  CNStageIntLLRInputS0xD(257)(5) <= LUT_4bit_to_3bit(ChLLRxDI(359));
  CNStageIntLLRInputS0xD(283)(5) <= LUT_4bit_to_3bit(ChLLRxDI(359));
  CNStageIntLLRInputS0xD(372)(5) <= LUT_4bit_to_3bit(ChLLRxDI(359));
  CNStageIntLLRInputS0xD(14)(5) <= LUT_4bit_to_3bit(ChLLRxDI(360));
  CNStageIntLLRInputS0xD(91)(5) <= LUT_4bit_to_3bit(ChLLRxDI(360));
  CNStageIntLLRInputS0xD(116)(5) <= LUT_4bit_to_3bit(ChLLRxDI(360));
  CNStageIntLLRInputS0xD(174)(5) <= LUT_4bit_to_3bit(ChLLRxDI(360));
  CNStageIntLLRInputS0xD(248)(5) <= LUT_4bit_to_3bit(ChLLRxDI(360));
  CNStageIntLLRInputS0xD(292)(5) <= LUT_4bit_to_3bit(ChLLRxDI(360));
  CNStageIntLLRInputS0xD(345)(5) <= LUT_4bit_to_3bit(ChLLRxDI(360));
  CNStageIntLLRInputS0xD(13)(5) <= LUT_4bit_to_3bit(ChLLRxDI(361));
  CNStageIntLLRInputS0xD(54)(5) <= LUT_4bit_to_3bit(ChLLRxDI(361));
  CNStageIntLLRInputS0xD(120)(5) <= LUT_4bit_to_3bit(ChLLRxDI(361));
  CNStageIntLLRInputS0xD(207)(5) <= LUT_4bit_to_3bit(ChLLRxDI(361));
  CNStageIntLLRInputS0xD(271)(5) <= LUT_4bit_to_3bit(ChLLRxDI(361));
  CNStageIntLLRInputS0xD(285)(5) <= LUT_4bit_to_3bit(ChLLRxDI(361));
  CNStageIntLLRInputS0xD(342)(5) <= LUT_4bit_to_3bit(ChLLRxDI(361));
  CNStageIntLLRInputS0xD(12)(5) <= LUT_4bit_to_3bit(ChLLRxDI(362));
  CNStageIntLLRInputS0xD(55)(5) <= LUT_4bit_to_3bit(ChLLRxDI(362));
  CNStageIntLLRInputS0xD(169)(5) <= LUT_4bit_to_3bit(ChLLRxDI(362));
  CNStageIntLLRInputS0xD(210)(5) <= LUT_4bit_to_3bit(ChLLRxDI(362));
  CNStageIntLLRInputS0xD(276)(5) <= LUT_4bit_to_3bit(ChLLRxDI(362));
  CNStageIntLLRInputS0xD(289)(5) <= LUT_4bit_to_3bit(ChLLRxDI(362));
  CNStageIntLLRInputS0xD(357)(5) <= LUT_4bit_to_3bit(ChLLRxDI(362));
  CNStageIntLLRInputS0xD(90)(5) <= LUT_4bit_to_3bit(ChLLRxDI(363));
  CNStageIntLLRInputS0xD(147)(5) <= LUT_4bit_to_3bit(ChLLRxDI(363));
  CNStageIntLLRInputS0xD(197)(5) <= LUT_4bit_to_3bit(ChLLRxDI(363));
  CNStageIntLLRInputS0xD(261)(5) <= LUT_4bit_to_3bit(ChLLRxDI(363));
  CNStageIntLLRInputS0xD(281)(5) <= LUT_4bit_to_3bit(ChLLRxDI(363));
  CNStageIntLLRInputS0xD(11)(5) <= LUT_4bit_to_3bit(ChLLRxDI(364));
  CNStageIntLLRInputS0xD(82)(5) <= LUT_4bit_to_3bit(ChLLRxDI(364));
  CNStageIntLLRInputS0xD(129)(5) <= LUT_4bit_to_3bit(ChLLRxDI(364));
  CNStageIntLLRInputS0xD(175)(5) <= LUT_4bit_to_3bit(ChLLRxDI(364));
  CNStageIntLLRInputS0xD(263)(5) <= LUT_4bit_to_3bit(ChLLRxDI(364));
  CNStageIntLLRInputS0xD(313)(5) <= LUT_4bit_to_3bit(ChLLRxDI(364));
  CNStageIntLLRInputS0xD(10)(5) <= LUT_4bit_to_3bit(ChLLRxDI(365));
  CNStageIntLLRInputS0xD(98)(5) <= LUT_4bit_to_3bit(ChLLRxDI(365));
  CNStageIntLLRInputS0xD(142)(5) <= LUT_4bit_to_3bit(ChLLRxDI(365));
  CNStageIntLLRInputS0xD(194)(5) <= LUT_4bit_to_3bit(ChLLRxDI(365));
  CNStageIntLLRInputS0xD(234)(5) <= LUT_4bit_to_3bit(ChLLRxDI(365));
  CNStageIntLLRInputS0xD(298)(5) <= LUT_4bit_to_3bit(ChLLRxDI(365));
  CNStageIntLLRInputS0xD(9)(5) <= LUT_4bit_to_3bit(ChLLRxDI(366));
  CNStageIntLLRInputS0xD(102)(5) <= LUT_4bit_to_3bit(ChLLRxDI(366));
  CNStageIntLLRInputS0xD(153)(5) <= LUT_4bit_to_3bit(ChLLRxDI(366));
  CNStageIntLLRInputS0xD(219)(5) <= LUT_4bit_to_3bit(ChLLRxDI(366));
  CNStageIntLLRInputS0xD(269)(5) <= LUT_4bit_to_3bit(ChLLRxDI(366));
  CNStageIntLLRInputS0xD(308)(5) <= LUT_4bit_to_3bit(ChLLRxDI(366));
  CNStageIntLLRInputS0xD(8)(5) <= LUT_4bit_to_3bit(ChLLRxDI(367));
  CNStageIntLLRInputS0xD(110)(5) <= LUT_4bit_to_3bit(ChLLRxDI(367));
  CNStageIntLLRInputS0xD(123)(5) <= LUT_4bit_to_3bit(ChLLRxDI(367));
  CNStageIntLLRInputS0xD(205)(5) <= LUT_4bit_to_3bit(ChLLRxDI(367));
  CNStageIntLLRInputS0xD(226)(5) <= LUT_4bit_to_3bit(ChLLRxDI(367));
  CNStageIntLLRInputS0xD(320)(5) <= LUT_4bit_to_3bit(ChLLRxDI(367));
  CNStageIntLLRInputS0xD(333)(5) <= LUT_4bit_to_3bit(ChLLRxDI(367));
  CNStageIntLLRInputS0xD(7)(5) <= LUT_4bit_to_3bit(ChLLRxDI(368));
  CNStageIntLLRInputS0xD(177)(5) <= LUT_4bit_to_3bit(ChLLRxDI(368));
  CNStageIntLLRInputS0xD(381)(5) <= LUT_4bit_to_3bit(ChLLRxDI(368));
  CNStageIntLLRInputS0xD(6)(5) <= LUT_4bit_to_3bit(ChLLRxDI(369));
  CNStageIntLLRInputS0xD(156)(5) <= LUT_4bit_to_3bit(ChLLRxDI(369));
  CNStageIntLLRInputS0xD(221)(5) <= LUT_4bit_to_3bit(ChLLRxDI(369));
  CNStageIntLLRInputS0xD(262)(5) <= LUT_4bit_to_3bit(ChLLRxDI(369));
  CNStageIntLLRInputS0xD(358)(5) <= LUT_4bit_to_3bit(ChLLRxDI(369));
  CNStageIntLLRInputS0xD(5)(5) <= LUT_4bit_to_3bit(ChLLRxDI(370));
  CNStageIntLLRInputS0xD(114)(5) <= LUT_4bit_to_3bit(ChLLRxDI(370));
  CNStageIntLLRInputS0xD(208)(5) <= LUT_4bit_to_3bit(ChLLRxDI(370));
  CNStageIntLLRInputS0xD(275)(5) <= LUT_4bit_to_3bit(ChLLRxDI(370));
  CNStageIntLLRInputS0xD(341)(5) <= LUT_4bit_to_3bit(ChLLRxDI(370));
  CNStageIntLLRInputS0xD(4)(5) <= LUT_4bit_to_3bit(ChLLRxDI(371));
  CNStageIntLLRInputS0xD(135)(5) <= LUT_4bit_to_3bit(ChLLRxDI(371));
  CNStageIntLLRInputS0xD(173)(5) <= LUT_4bit_to_3bit(ChLLRxDI(371));
  CNStageIntLLRInputS0xD(249)(5) <= LUT_4bit_to_3bit(ChLLRxDI(371));
  CNStageIntLLRInputS0xD(354)(5) <= LUT_4bit_to_3bit(ChLLRxDI(371));
  CNStageIntLLRInputS0xD(106)(5) <= LUT_4bit_to_3bit(ChLLRxDI(372));
  CNStageIntLLRInputS0xD(144)(5) <= LUT_4bit_to_3bit(ChLLRxDI(372));
  CNStageIntLLRInputS0xD(201)(5) <= LUT_4bit_to_3bit(ChLLRxDI(372));
  CNStageIntLLRInputS0xD(229)(5) <= LUT_4bit_to_3bit(ChLLRxDI(372));
  CNStageIntLLRInputS0xD(301)(5) <= LUT_4bit_to_3bit(ChLLRxDI(372));
  CNStageIntLLRInputS0xD(365)(5) <= LUT_4bit_to_3bit(ChLLRxDI(372));
  CNStageIntLLRInputS0xD(3)(5) <= LUT_4bit_to_3bit(ChLLRxDI(373));
  CNStageIntLLRInputS0xD(139)(5) <= LUT_4bit_to_3bit(ChLLRxDI(373));
  CNStageIntLLRInputS0xD(250)(5) <= LUT_4bit_to_3bit(ChLLRxDI(373));
  CNStageIntLLRInputS0xD(310)(5) <= LUT_4bit_to_3bit(ChLLRxDI(373));
  CNStageIntLLRInputS0xD(335)(5) <= LUT_4bit_to_3bit(ChLLRxDI(373));
  CNStageIntLLRInputS0xD(2)(5) <= LUT_4bit_to_3bit(ChLLRxDI(374));
  CNStageIntLLRInputS0xD(85)(5) <= LUT_4bit_to_3bit(ChLLRxDI(374));
  CNStageIntLLRInputS0xD(145)(5) <= LUT_4bit_to_3bit(ChLLRxDI(374));
  CNStageIntLLRInputS0xD(213)(5) <= LUT_4bit_to_3bit(ChLLRxDI(374));
  CNStageIntLLRInputS0xD(264)(5) <= LUT_4bit_to_3bit(ChLLRxDI(374));
  CNStageIntLLRInputS0xD(306)(5) <= LUT_4bit_to_3bit(ChLLRxDI(374));
  CNStageIntLLRInputS0xD(383)(5) <= LUT_4bit_to_3bit(ChLLRxDI(374));
  CNStageIntLLRInputS0xD(1)(5) <= LUT_4bit_to_3bit(ChLLRxDI(375));
  CNStageIntLLRInputS0xD(64)(5) <= LUT_4bit_to_3bit(ChLLRxDI(375));
  CNStageIntLLRInputS0xD(134)(5) <= LUT_4bit_to_3bit(ChLLRxDI(375));
  CNStageIntLLRInputS0xD(260)(5) <= LUT_4bit_to_3bit(ChLLRxDI(375));
  CNStageIntLLRInputS0xD(311)(5) <= LUT_4bit_to_3bit(ChLLRxDI(375));
  CNStageIntLLRInputS0xD(368)(5) <= LUT_4bit_to_3bit(ChLLRxDI(375));
  CNStageIntLLRInputS0xD(0)(5) <= LUT_4bit_to_3bit(ChLLRxDI(376));
  CNStageIntLLRInputS0xD(67)(5) <= LUT_4bit_to_3bit(ChLLRxDI(376));
  CNStageIntLLRInputS0xD(159)(5) <= LUT_4bit_to_3bit(ChLLRxDI(376));
  CNStageIntLLRInputS0xD(278)(5) <= LUT_4bit_to_3bit(ChLLRxDI(376));
  CNStageIntLLRInputS0xD(107)(5) <= LUT_4bit_to_3bit(ChLLRxDI(377));
  CNStageIntLLRInputS0xD(166)(5) <= LUT_4bit_to_3bit(ChLLRxDI(377));
  CNStageIntLLRInputS0xD(193)(5) <= LUT_4bit_to_3bit(ChLLRxDI(377));
  CNStageIntLLRInputS0xD(325)(5) <= LUT_4bit_to_3bit(ChLLRxDI(377));
  CNStageIntLLRInputS0xD(347)(5) <= LUT_4bit_to_3bit(ChLLRxDI(377));
  CNStageIntLLRInputS0xD(86)(5) <= LUT_4bit_to_3bit(ChLLRxDI(378));
  CNStageIntLLRInputS0xD(149)(5) <= LUT_4bit_to_3bit(ChLLRxDI(378));
  CNStageIntLLRInputS0xD(187)(5) <= LUT_4bit_to_3bit(ChLLRxDI(378));
  CNStageIntLLRInputS0xD(246)(5) <= LUT_4bit_to_3bit(ChLLRxDI(378));
  CNStageIntLLRInputS0xD(331)(5) <= LUT_4bit_to_3bit(ChLLRxDI(378));
  CNStageIntLLRInputS0xD(355)(5) <= LUT_4bit_to_3bit(ChLLRxDI(378));
  CNStageIntLLRInputS0xD(105)(5) <= LUT_4bit_to_3bit(ChLLRxDI(379));
  CNStageIntLLRInputS0xD(151)(5) <= LUT_4bit_to_3bit(ChLLRxDI(379));
  CNStageIntLLRInputS0xD(277)(5) <= LUT_4bit_to_3bit(ChLLRxDI(379));
  CNStageIntLLRInputS0xD(315)(5) <= LUT_4bit_to_3bit(ChLLRxDI(379));
  CNStageIntLLRInputS0xD(351)(5) <= LUT_4bit_to_3bit(ChLLRxDI(379));
  CNStageIntLLRInputS0xD(77)(5) <= LUT_4bit_to_3bit(ChLLRxDI(380));
  CNStageIntLLRInputS0xD(118)(5) <= LUT_4bit_to_3bit(ChLLRxDI(380));
  CNStageIntLLRInputS0xD(182)(5) <= LUT_4bit_to_3bit(ChLLRxDI(380));
  CNStageIntLLRInputS0xD(270)(5) <= LUT_4bit_to_3bit(ChLLRxDI(380));
  CNStageIntLLRInputS0xD(317)(5) <= LUT_4bit_to_3bit(ChLLRxDI(380));
  CNStageIntLLRInputS0xD(356)(5) <= LUT_4bit_to_3bit(ChLLRxDI(380));
  CNStageIntLLRInputS0xD(60)(5) <= LUT_4bit_to_3bit(ChLLRxDI(381));
  CNStageIntLLRInputS0xD(157)(5) <= LUT_4bit_to_3bit(ChLLRxDI(381));
  CNStageIntLLRInputS0xD(214)(5) <= LUT_4bit_to_3bit(ChLLRxDI(381));
  CNStageIntLLRInputS0xD(233)(5) <= LUT_4bit_to_3bit(ChLLRxDI(381));
  CNStageIntLLRInputS0xD(287)(5) <= LUT_4bit_to_3bit(ChLLRxDI(381));
  CNStageIntLLRInputS0xD(346)(5) <= LUT_4bit_to_3bit(ChLLRxDI(381));
  CNStageIntLLRInputS0xD(87)(5) <= LUT_4bit_to_3bit(ChLLRxDI(382));
  CNStageIntLLRInputS0xD(111)(5) <= LUT_4bit_to_3bit(ChLLRxDI(382));
  CNStageIntLLRInputS0xD(198)(5) <= LUT_4bit_to_3bit(ChLLRxDI(382));
  CNStageIntLLRInputS0xD(237)(5) <= LUT_4bit_to_3bit(ChLLRxDI(382));
  CNStageIntLLRInputS0xD(323)(5) <= LUT_4bit_to_3bit(ChLLRxDI(382));
  CNStageIntLLRInputS0xD(371)(5) <= LUT_4bit_to_3bit(ChLLRxDI(382));
  CNStageIntLLRInputS0xD(52)(5) <= LUT_4bit_to_3bit(ChLLRxDI(383));
  CNStageIntLLRInputS0xD(79)(5) <= LUT_4bit_to_3bit(ChLLRxDI(383));
  CNStageIntLLRInputS0xD(119)(5) <= LUT_4bit_to_3bit(ChLLRxDI(383));
  CNStageIntLLRInputS0xD(209)(5) <= LUT_4bit_to_3bit(ChLLRxDI(383));
  CNStageIntLLRInputS0xD(279)(5) <= LUT_4bit_to_3bit(ChLLRxDI(383));
  CNStageIntLLRInputS0xD(282)(5) <= LUT_4bit_to_3bit(ChLLRxDI(383));
  CNStageIntLLRInputS0xD(378)(5) <= LUT_4bit_to_3bit(ChLLRxDI(383));

  -- Connect output channel LLRs of stages with input channel LLRs of following stages
  CNStageChLLRInputS0xD <= ChLLRxDI;
  VNStageChLLRInputS0xD <= CNStageChLLROutputS0xD;
  CNStageChLLRInputS1xD <= VNStageChLLROutputS0xD;
  VNStageChLLRInputS1xD <= CNStageChLLROutputS1xD;
  CNStageChLLRInputS2xD <= VNStageChLLROutputS1xD;
  VNStageChLLRInputS2xD <= CNStageChLLROutputS2xD;
  CNStageChLLRInputS3xD <= VNStageChLLROutputS2xD;
  VNStageChLLRInputS3xD <= CNStageChLLROutputS3xD;
  CNStageChLLRInputS4xD <= VNStageChLLROutputS3xD;
  VNStageChLLRInputS4xD <= CNStageChLLROutputS4xD;
  CNStageChLLRInputS5xD <= VNStageChLLROutputS4xD;
  VNStageChLLRInputS5xD <= CNStageChLLROutputS5xD;
  CNStageChLLRInputS6xD <= VNStageChLLROutputS5xD;
  VNStageChLLRInputS6xD <= CNStageChLLROutputS6xD;
  CNStageChLLRInputS7xD <= VNStageChLLROutputS6xD;
  VNStageChLLRInputS7xD <= CNStageChLLROutputS7xD;

-- Connect CN and VN stages

  -- Variable Nodes (Iteration 0)
  VNStageIntLLRInputS0xD(56)(0) <= CNStageIntLLROutputS0xD(0)(0);
  VNStageIntLLRInputS0xD(120)(0) <= CNStageIntLLROutputS0xD(0)(1);
  VNStageIntLLRInputS0xD(184)(0) <= CNStageIntLLROutputS0xD(0)(2);
  VNStageIntLLRInputS0xD(248)(0) <= CNStageIntLLROutputS0xD(0)(3);
  VNStageIntLLRInputS0xD(312)(0) <= CNStageIntLLROutputS0xD(0)(4);
  VNStageIntLLRInputS0xD(376)(0) <= CNStageIntLLROutputS0xD(0)(5);
  VNStageIntLLRInputS0xD(55)(0) <= CNStageIntLLROutputS0xD(1)(0);
  VNStageIntLLRInputS0xD(119)(0) <= CNStageIntLLROutputS0xD(1)(1);
  VNStageIntLLRInputS0xD(183)(0) <= CNStageIntLLROutputS0xD(1)(2);
  VNStageIntLLRInputS0xD(247)(0) <= CNStageIntLLROutputS0xD(1)(3);
  VNStageIntLLRInputS0xD(311)(0) <= CNStageIntLLROutputS0xD(1)(4);
  VNStageIntLLRInputS0xD(375)(0) <= CNStageIntLLROutputS0xD(1)(5);
  VNStageIntLLRInputS0xD(54)(0) <= CNStageIntLLROutputS0xD(2)(0);
  VNStageIntLLRInputS0xD(118)(0) <= CNStageIntLLROutputS0xD(2)(1);
  VNStageIntLLRInputS0xD(182)(0) <= CNStageIntLLROutputS0xD(2)(2);
  VNStageIntLLRInputS0xD(246)(0) <= CNStageIntLLROutputS0xD(2)(3);
  VNStageIntLLRInputS0xD(310)(0) <= CNStageIntLLROutputS0xD(2)(4);
  VNStageIntLLRInputS0xD(374)(0) <= CNStageIntLLROutputS0xD(2)(5);
  VNStageIntLLRInputS0xD(53)(0) <= CNStageIntLLROutputS0xD(3)(0);
  VNStageIntLLRInputS0xD(117)(0) <= CNStageIntLLROutputS0xD(3)(1);
  VNStageIntLLRInputS0xD(181)(0) <= CNStageIntLLROutputS0xD(3)(2);
  VNStageIntLLRInputS0xD(245)(0) <= CNStageIntLLROutputS0xD(3)(3);
  VNStageIntLLRInputS0xD(309)(0) <= CNStageIntLLROutputS0xD(3)(4);
  VNStageIntLLRInputS0xD(373)(0) <= CNStageIntLLROutputS0xD(3)(5);
  VNStageIntLLRInputS0xD(51)(0) <= CNStageIntLLROutputS0xD(4)(0);
  VNStageIntLLRInputS0xD(115)(0) <= CNStageIntLLROutputS0xD(4)(1);
  VNStageIntLLRInputS0xD(179)(0) <= CNStageIntLLROutputS0xD(4)(2);
  VNStageIntLLRInputS0xD(243)(0) <= CNStageIntLLROutputS0xD(4)(3);
  VNStageIntLLRInputS0xD(307)(0) <= CNStageIntLLROutputS0xD(4)(4);
  VNStageIntLLRInputS0xD(371)(0) <= CNStageIntLLROutputS0xD(4)(5);
  VNStageIntLLRInputS0xD(50)(0) <= CNStageIntLLROutputS0xD(5)(0);
  VNStageIntLLRInputS0xD(114)(0) <= CNStageIntLLROutputS0xD(5)(1);
  VNStageIntLLRInputS0xD(178)(0) <= CNStageIntLLROutputS0xD(5)(2);
  VNStageIntLLRInputS0xD(242)(0) <= CNStageIntLLROutputS0xD(5)(3);
  VNStageIntLLRInputS0xD(306)(0) <= CNStageIntLLROutputS0xD(5)(4);
  VNStageIntLLRInputS0xD(370)(0) <= CNStageIntLLROutputS0xD(5)(5);
  VNStageIntLLRInputS0xD(49)(0) <= CNStageIntLLROutputS0xD(6)(0);
  VNStageIntLLRInputS0xD(113)(0) <= CNStageIntLLROutputS0xD(6)(1);
  VNStageIntLLRInputS0xD(177)(0) <= CNStageIntLLROutputS0xD(6)(2);
  VNStageIntLLRInputS0xD(241)(0) <= CNStageIntLLROutputS0xD(6)(3);
  VNStageIntLLRInputS0xD(305)(0) <= CNStageIntLLROutputS0xD(6)(4);
  VNStageIntLLRInputS0xD(369)(0) <= CNStageIntLLROutputS0xD(6)(5);
  VNStageIntLLRInputS0xD(48)(0) <= CNStageIntLLROutputS0xD(7)(0);
  VNStageIntLLRInputS0xD(112)(0) <= CNStageIntLLROutputS0xD(7)(1);
  VNStageIntLLRInputS0xD(176)(0) <= CNStageIntLLROutputS0xD(7)(2);
  VNStageIntLLRInputS0xD(240)(0) <= CNStageIntLLROutputS0xD(7)(3);
  VNStageIntLLRInputS0xD(304)(0) <= CNStageIntLLROutputS0xD(7)(4);
  VNStageIntLLRInputS0xD(368)(0) <= CNStageIntLLROutputS0xD(7)(5);
  VNStageIntLLRInputS0xD(47)(0) <= CNStageIntLLROutputS0xD(8)(0);
  VNStageIntLLRInputS0xD(111)(0) <= CNStageIntLLROutputS0xD(8)(1);
  VNStageIntLLRInputS0xD(175)(0) <= CNStageIntLLROutputS0xD(8)(2);
  VNStageIntLLRInputS0xD(239)(0) <= CNStageIntLLROutputS0xD(8)(3);
  VNStageIntLLRInputS0xD(303)(0) <= CNStageIntLLROutputS0xD(8)(4);
  VNStageIntLLRInputS0xD(367)(0) <= CNStageIntLLROutputS0xD(8)(5);
  VNStageIntLLRInputS0xD(46)(0) <= CNStageIntLLROutputS0xD(9)(0);
  VNStageIntLLRInputS0xD(110)(0) <= CNStageIntLLROutputS0xD(9)(1);
  VNStageIntLLRInputS0xD(174)(0) <= CNStageIntLLROutputS0xD(9)(2);
  VNStageIntLLRInputS0xD(238)(0) <= CNStageIntLLROutputS0xD(9)(3);
  VNStageIntLLRInputS0xD(302)(0) <= CNStageIntLLROutputS0xD(9)(4);
  VNStageIntLLRInputS0xD(366)(0) <= CNStageIntLLROutputS0xD(9)(5);
  VNStageIntLLRInputS0xD(45)(0) <= CNStageIntLLROutputS0xD(10)(0);
  VNStageIntLLRInputS0xD(109)(0) <= CNStageIntLLROutputS0xD(10)(1);
  VNStageIntLLRInputS0xD(173)(0) <= CNStageIntLLROutputS0xD(10)(2);
  VNStageIntLLRInputS0xD(237)(0) <= CNStageIntLLROutputS0xD(10)(3);
  VNStageIntLLRInputS0xD(301)(0) <= CNStageIntLLROutputS0xD(10)(4);
  VNStageIntLLRInputS0xD(365)(0) <= CNStageIntLLROutputS0xD(10)(5);
  VNStageIntLLRInputS0xD(44)(0) <= CNStageIntLLROutputS0xD(11)(0);
  VNStageIntLLRInputS0xD(108)(0) <= CNStageIntLLROutputS0xD(11)(1);
  VNStageIntLLRInputS0xD(172)(0) <= CNStageIntLLROutputS0xD(11)(2);
  VNStageIntLLRInputS0xD(236)(0) <= CNStageIntLLROutputS0xD(11)(3);
  VNStageIntLLRInputS0xD(300)(0) <= CNStageIntLLROutputS0xD(11)(4);
  VNStageIntLLRInputS0xD(364)(0) <= CNStageIntLLROutputS0xD(11)(5);
  VNStageIntLLRInputS0xD(42)(0) <= CNStageIntLLROutputS0xD(12)(0);
  VNStageIntLLRInputS0xD(106)(0) <= CNStageIntLLROutputS0xD(12)(1);
  VNStageIntLLRInputS0xD(170)(0) <= CNStageIntLLROutputS0xD(12)(2);
  VNStageIntLLRInputS0xD(234)(0) <= CNStageIntLLROutputS0xD(12)(3);
  VNStageIntLLRInputS0xD(298)(0) <= CNStageIntLLROutputS0xD(12)(4);
  VNStageIntLLRInputS0xD(362)(0) <= CNStageIntLLROutputS0xD(12)(5);
  VNStageIntLLRInputS0xD(41)(0) <= CNStageIntLLROutputS0xD(13)(0);
  VNStageIntLLRInputS0xD(105)(0) <= CNStageIntLLROutputS0xD(13)(1);
  VNStageIntLLRInputS0xD(169)(0) <= CNStageIntLLROutputS0xD(13)(2);
  VNStageIntLLRInputS0xD(233)(0) <= CNStageIntLLROutputS0xD(13)(3);
  VNStageIntLLRInputS0xD(297)(0) <= CNStageIntLLROutputS0xD(13)(4);
  VNStageIntLLRInputS0xD(361)(0) <= CNStageIntLLROutputS0xD(13)(5);
  VNStageIntLLRInputS0xD(40)(0) <= CNStageIntLLROutputS0xD(14)(0);
  VNStageIntLLRInputS0xD(104)(0) <= CNStageIntLLROutputS0xD(14)(1);
  VNStageIntLLRInputS0xD(168)(0) <= CNStageIntLLROutputS0xD(14)(2);
  VNStageIntLLRInputS0xD(232)(0) <= CNStageIntLLROutputS0xD(14)(3);
  VNStageIntLLRInputS0xD(296)(0) <= CNStageIntLLROutputS0xD(14)(4);
  VNStageIntLLRInputS0xD(360)(0) <= CNStageIntLLROutputS0xD(14)(5);
  VNStageIntLLRInputS0xD(39)(0) <= CNStageIntLLROutputS0xD(15)(0);
  VNStageIntLLRInputS0xD(103)(0) <= CNStageIntLLROutputS0xD(15)(1);
  VNStageIntLLRInputS0xD(167)(0) <= CNStageIntLLROutputS0xD(15)(2);
  VNStageIntLLRInputS0xD(231)(0) <= CNStageIntLLROutputS0xD(15)(3);
  VNStageIntLLRInputS0xD(295)(0) <= CNStageIntLLROutputS0xD(15)(4);
  VNStageIntLLRInputS0xD(359)(0) <= CNStageIntLLROutputS0xD(15)(5);
  VNStageIntLLRInputS0xD(38)(0) <= CNStageIntLLROutputS0xD(16)(0);
  VNStageIntLLRInputS0xD(102)(0) <= CNStageIntLLROutputS0xD(16)(1);
  VNStageIntLLRInputS0xD(166)(0) <= CNStageIntLLROutputS0xD(16)(2);
  VNStageIntLLRInputS0xD(230)(0) <= CNStageIntLLROutputS0xD(16)(3);
  VNStageIntLLRInputS0xD(294)(0) <= CNStageIntLLROutputS0xD(16)(4);
  VNStageIntLLRInputS0xD(358)(0) <= CNStageIntLLROutputS0xD(16)(5);
  VNStageIntLLRInputS0xD(37)(0) <= CNStageIntLLROutputS0xD(17)(0);
  VNStageIntLLRInputS0xD(101)(0) <= CNStageIntLLROutputS0xD(17)(1);
  VNStageIntLLRInputS0xD(165)(0) <= CNStageIntLLROutputS0xD(17)(2);
  VNStageIntLLRInputS0xD(229)(0) <= CNStageIntLLROutputS0xD(17)(3);
  VNStageIntLLRInputS0xD(293)(0) <= CNStageIntLLROutputS0xD(17)(4);
  VNStageIntLLRInputS0xD(357)(0) <= CNStageIntLLROutputS0xD(17)(5);
  VNStageIntLLRInputS0xD(36)(0) <= CNStageIntLLROutputS0xD(18)(0);
  VNStageIntLLRInputS0xD(100)(0) <= CNStageIntLLROutputS0xD(18)(1);
  VNStageIntLLRInputS0xD(164)(0) <= CNStageIntLLROutputS0xD(18)(2);
  VNStageIntLLRInputS0xD(228)(0) <= CNStageIntLLROutputS0xD(18)(3);
  VNStageIntLLRInputS0xD(292)(0) <= CNStageIntLLROutputS0xD(18)(4);
  VNStageIntLLRInputS0xD(356)(0) <= CNStageIntLLROutputS0xD(18)(5);
  VNStageIntLLRInputS0xD(35)(0) <= CNStageIntLLROutputS0xD(19)(0);
  VNStageIntLLRInputS0xD(99)(0) <= CNStageIntLLROutputS0xD(19)(1);
  VNStageIntLLRInputS0xD(163)(0) <= CNStageIntLLROutputS0xD(19)(2);
  VNStageIntLLRInputS0xD(227)(0) <= CNStageIntLLROutputS0xD(19)(3);
  VNStageIntLLRInputS0xD(291)(0) <= CNStageIntLLROutputS0xD(19)(4);
  VNStageIntLLRInputS0xD(355)(0) <= CNStageIntLLROutputS0xD(19)(5);
  VNStageIntLLRInputS0xD(34)(0) <= CNStageIntLLROutputS0xD(20)(0);
  VNStageIntLLRInputS0xD(98)(0) <= CNStageIntLLROutputS0xD(20)(1);
  VNStageIntLLRInputS0xD(162)(0) <= CNStageIntLLROutputS0xD(20)(2);
  VNStageIntLLRInputS0xD(226)(0) <= CNStageIntLLROutputS0xD(20)(3);
  VNStageIntLLRInputS0xD(290)(0) <= CNStageIntLLROutputS0xD(20)(4);
  VNStageIntLLRInputS0xD(354)(0) <= CNStageIntLLROutputS0xD(20)(5);
  VNStageIntLLRInputS0xD(33)(0) <= CNStageIntLLROutputS0xD(21)(0);
  VNStageIntLLRInputS0xD(97)(0) <= CNStageIntLLROutputS0xD(21)(1);
  VNStageIntLLRInputS0xD(161)(0) <= CNStageIntLLROutputS0xD(21)(2);
  VNStageIntLLRInputS0xD(225)(0) <= CNStageIntLLROutputS0xD(21)(3);
  VNStageIntLLRInputS0xD(289)(0) <= CNStageIntLLROutputS0xD(21)(4);
  VNStageIntLLRInputS0xD(353)(0) <= CNStageIntLLROutputS0xD(21)(5);
  VNStageIntLLRInputS0xD(32)(0) <= CNStageIntLLROutputS0xD(22)(0);
  VNStageIntLLRInputS0xD(96)(0) <= CNStageIntLLROutputS0xD(22)(1);
  VNStageIntLLRInputS0xD(160)(0) <= CNStageIntLLROutputS0xD(22)(2);
  VNStageIntLLRInputS0xD(224)(0) <= CNStageIntLLROutputS0xD(22)(3);
  VNStageIntLLRInputS0xD(288)(0) <= CNStageIntLLROutputS0xD(22)(4);
  VNStageIntLLRInputS0xD(352)(0) <= CNStageIntLLROutputS0xD(22)(5);
  VNStageIntLLRInputS0xD(31)(0) <= CNStageIntLLROutputS0xD(23)(0);
  VNStageIntLLRInputS0xD(95)(0) <= CNStageIntLLROutputS0xD(23)(1);
  VNStageIntLLRInputS0xD(159)(0) <= CNStageIntLLROutputS0xD(23)(2);
  VNStageIntLLRInputS0xD(223)(0) <= CNStageIntLLROutputS0xD(23)(3);
  VNStageIntLLRInputS0xD(287)(0) <= CNStageIntLLROutputS0xD(23)(4);
  VNStageIntLLRInputS0xD(351)(0) <= CNStageIntLLROutputS0xD(23)(5);
  VNStageIntLLRInputS0xD(30)(0) <= CNStageIntLLROutputS0xD(24)(0);
  VNStageIntLLRInputS0xD(94)(0) <= CNStageIntLLROutputS0xD(24)(1);
  VNStageIntLLRInputS0xD(158)(0) <= CNStageIntLLROutputS0xD(24)(2);
  VNStageIntLLRInputS0xD(222)(0) <= CNStageIntLLROutputS0xD(24)(3);
  VNStageIntLLRInputS0xD(286)(0) <= CNStageIntLLROutputS0xD(24)(4);
  VNStageIntLLRInputS0xD(350)(0) <= CNStageIntLLROutputS0xD(24)(5);
  VNStageIntLLRInputS0xD(29)(0) <= CNStageIntLLROutputS0xD(25)(0);
  VNStageIntLLRInputS0xD(93)(0) <= CNStageIntLLROutputS0xD(25)(1);
  VNStageIntLLRInputS0xD(157)(0) <= CNStageIntLLROutputS0xD(25)(2);
  VNStageIntLLRInputS0xD(221)(0) <= CNStageIntLLROutputS0xD(25)(3);
  VNStageIntLLRInputS0xD(285)(0) <= CNStageIntLLROutputS0xD(25)(4);
  VNStageIntLLRInputS0xD(349)(0) <= CNStageIntLLROutputS0xD(25)(5);
  VNStageIntLLRInputS0xD(28)(0) <= CNStageIntLLROutputS0xD(26)(0);
  VNStageIntLLRInputS0xD(92)(0) <= CNStageIntLLROutputS0xD(26)(1);
  VNStageIntLLRInputS0xD(156)(0) <= CNStageIntLLROutputS0xD(26)(2);
  VNStageIntLLRInputS0xD(220)(0) <= CNStageIntLLROutputS0xD(26)(3);
  VNStageIntLLRInputS0xD(284)(0) <= CNStageIntLLROutputS0xD(26)(4);
  VNStageIntLLRInputS0xD(348)(0) <= CNStageIntLLROutputS0xD(26)(5);
  VNStageIntLLRInputS0xD(27)(0) <= CNStageIntLLROutputS0xD(27)(0);
  VNStageIntLLRInputS0xD(91)(0) <= CNStageIntLLROutputS0xD(27)(1);
  VNStageIntLLRInputS0xD(155)(0) <= CNStageIntLLROutputS0xD(27)(2);
  VNStageIntLLRInputS0xD(219)(0) <= CNStageIntLLROutputS0xD(27)(3);
  VNStageIntLLRInputS0xD(283)(0) <= CNStageIntLLROutputS0xD(27)(4);
  VNStageIntLLRInputS0xD(347)(0) <= CNStageIntLLROutputS0xD(27)(5);
  VNStageIntLLRInputS0xD(26)(0) <= CNStageIntLLROutputS0xD(28)(0);
  VNStageIntLLRInputS0xD(90)(0) <= CNStageIntLLROutputS0xD(28)(1);
  VNStageIntLLRInputS0xD(154)(0) <= CNStageIntLLROutputS0xD(28)(2);
  VNStageIntLLRInputS0xD(218)(0) <= CNStageIntLLROutputS0xD(28)(3);
  VNStageIntLLRInputS0xD(282)(0) <= CNStageIntLLROutputS0xD(28)(4);
  VNStageIntLLRInputS0xD(346)(0) <= CNStageIntLLROutputS0xD(28)(5);
  VNStageIntLLRInputS0xD(25)(0) <= CNStageIntLLROutputS0xD(29)(0);
  VNStageIntLLRInputS0xD(89)(0) <= CNStageIntLLROutputS0xD(29)(1);
  VNStageIntLLRInputS0xD(153)(0) <= CNStageIntLLROutputS0xD(29)(2);
  VNStageIntLLRInputS0xD(217)(0) <= CNStageIntLLROutputS0xD(29)(3);
  VNStageIntLLRInputS0xD(281)(0) <= CNStageIntLLROutputS0xD(29)(4);
  VNStageIntLLRInputS0xD(345)(0) <= CNStageIntLLROutputS0xD(29)(5);
  VNStageIntLLRInputS0xD(24)(0) <= CNStageIntLLROutputS0xD(30)(0);
  VNStageIntLLRInputS0xD(88)(0) <= CNStageIntLLROutputS0xD(30)(1);
  VNStageIntLLRInputS0xD(152)(0) <= CNStageIntLLROutputS0xD(30)(2);
  VNStageIntLLRInputS0xD(216)(0) <= CNStageIntLLROutputS0xD(30)(3);
  VNStageIntLLRInputS0xD(280)(0) <= CNStageIntLLROutputS0xD(30)(4);
  VNStageIntLLRInputS0xD(344)(0) <= CNStageIntLLROutputS0xD(30)(5);
  VNStageIntLLRInputS0xD(23)(0) <= CNStageIntLLROutputS0xD(31)(0);
  VNStageIntLLRInputS0xD(87)(0) <= CNStageIntLLROutputS0xD(31)(1);
  VNStageIntLLRInputS0xD(151)(0) <= CNStageIntLLROutputS0xD(31)(2);
  VNStageIntLLRInputS0xD(215)(0) <= CNStageIntLLROutputS0xD(31)(3);
  VNStageIntLLRInputS0xD(279)(0) <= CNStageIntLLROutputS0xD(31)(4);
  VNStageIntLLRInputS0xD(343)(0) <= CNStageIntLLROutputS0xD(31)(5);
  VNStageIntLLRInputS0xD(22)(0) <= CNStageIntLLROutputS0xD(32)(0);
  VNStageIntLLRInputS0xD(86)(0) <= CNStageIntLLROutputS0xD(32)(1);
  VNStageIntLLRInputS0xD(150)(0) <= CNStageIntLLROutputS0xD(32)(2);
  VNStageIntLLRInputS0xD(214)(0) <= CNStageIntLLROutputS0xD(32)(3);
  VNStageIntLLRInputS0xD(278)(0) <= CNStageIntLLROutputS0xD(32)(4);
  VNStageIntLLRInputS0xD(342)(0) <= CNStageIntLLROutputS0xD(32)(5);
  VNStageIntLLRInputS0xD(21)(0) <= CNStageIntLLROutputS0xD(33)(0);
  VNStageIntLLRInputS0xD(85)(0) <= CNStageIntLLROutputS0xD(33)(1);
  VNStageIntLLRInputS0xD(149)(0) <= CNStageIntLLROutputS0xD(33)(2);
  VNStageIntLLRInputS0xD(213)(0) <= CNStageIntLLROutputS0xD(33)(3);
  VNStageIntLLRInputS0xD(277)(0) <= CNStageIntLLROutputS0xD(33)(4);
  VNStageIntLLRInputS0xD(341)(0) <= CNStageIntLLROutputS0xD(33)(5);
  VNStageIntLLRInputS0xD(20)(0) <= CNStageIntLLROutputS0xD(34)(0);
  VNStageIntLLRInputS0xD(84)(0) <= CNStageIntLLROutputS0xD(34)(1);
  VNStageIntLLRInputS0xD(148)(0) <= CNStageIntLLROutputS0xD(34)(2);
  VNStageIntLLRInputS0xD(212)(0) <= CNStageIntLLROutputS0xD(34)(3);
  VNStageIntLLRInputS0xD(276)(0) <= CNStageIntLLROutputS0xD(34)(4);
  VNStageIntLLRInputS0xD(340)(0) <= CNStageIntLLROutputS0xD(34)(5);
  VNStageIntLLRInputS0xD(19)(0) <= CNStageIntLLROutputS0xD(35)(0);
  VNStageIntLLRInputS0xD(83)(0) <= CNStageIntLLROutputS0xD(35)(1);
  VNStageIntLLRInputS0xD(147)(0) <= CNStageIntLLROutputS0xD(35)(2);
  VNStageIntLLRInputS0xD(211)(0) <= CNStageIntLLROutputS0xD(35)(3);
  VNStageIntLLRInputS0xD(275)(0) <= CNStageIntLLROutputS0xD(35)(4);
  VNStageIntLLRInputS0xD(339)(0) <= CNStageIntLLROutputS0xD(35)(5);
  VNStageIntLLRInputS0xD(18)(0) <= CNStageIntLLROutputS0xD(36)(0);
  VNStageIntLLRInputS0xD(82)(0) <= CNStageIntLLROutputS0xD(36)(1);
  VNStageIntLLRInputS0xD(146)(0) <= CNStageIntLLROutputS0xD(36)(2);
  VNStageIntLLRInputS0xD(210)(0) <= CNStageIntLLROutputS0xD(36)(3);
  VNStageIntLLRInputS0xD(274)(0) <= CNStageIntLLROutputS0xD(36)(4);
  VNStageIntLLRInputS0xD(338)(0) <= CNStageIntLLROutputS0xD(36)(5);
  VNStageIntLLRInputS0xD(17)(0) <= CNStageIntLLROutputS0xD(37)(0);
  VNStageIntLLRInputS0xD(81)(0) <= CNStageIntLLROutputS0xD(37)(1);
  VNStageIntLLRInputS0xD(145)(0) <= CNStageIntLLROutputS0xD(37)(2);
  VNStageIntLLRInputS0xD(209)(0) <= CNStageIntLLROutputS0xD(37)(3);
  VNStageIntLLRInputS0xD(273)(0) <= CNStageIntLLROutputS0xD(37)(4);
  VNStageIntLLRInputS0xD(337)(0) <= CNStageIntLLROutputS0xD(37)(5);
  VNStageIntLLRInputS0xD(16)(0) <= CNStageIntLLROutputS0xD(38)(0);
  VNStageIntLLRInputS0xD(80)(0) <= CNStageIntLLROutputS0xD(38)(1);
  VNStageIntLLRInputS0xD(144)(0) <= CNStageIntLLROutputS0xD(38)(2);
  VNStageIntLLRInputS0xD(208)(0) <= CNStageIntLLROutputS0xD(38)(3);
  VNStageIntLLRInputS0xD(272)(0) <= CNStageIntLLROutputS0xD(38)(4);
  VNStageIntLLRInputS0xD(336)(0) <= CNStageIntLLROutputS0xD(38)(5);
  VNStageIntLLRInputS0xD(15)(0) <= CNStageIntLLROutputS0xD(39)(0);
  VNStageIntLLRInputS0xD(79)(0) <= CNStageIntLLROutputS0xD(39)(1);
  VNStageIntLLRInputS0xD(143)(0) <= CNStageIntLLROutputS0xD(39)(2);
  VNStageIntLLRInputS0xD(207)(0) <= CNStageIntLLROutputS0xD(39)(3);
  VNStageIntLLRInputS0xD(271)(0) <= CNStageIntLLROutputS0xD(39)(4);
  VNStageIntLLRInputS0xD(335)(0) <= CNStageIntLLROutputS0xD(39)(5);
  VNStageIntLLRInputS0xD(14)(0) <= CNStageIntLLROutputS0xD(40)(0);
  VNStageIntLLRInputS0xD(78)(0) <= CNStageIntLLROutputS0xD(40)(1);
  VNStageIntLLRInputS0xD(142)(0) <= CNStageIntLLROutputS0xD(40)(2);
  VNStageIntLLRInputS0xD(206)(0) <= CNStageIntLLROutputS0xD(40)(3);
  VNStageIntLLRInputS0xD(270)(0) <= CNStageIntLLROutputS0xD(40)(4);
  VNStageIntLLRInputS0xD(334)(0) <= CNStageIntLLROutputS0xD(40)(5);
  VNStageIntLLRInputS0xD(12)(0) <= CNStageIntLLROutputS0xD(41)(0);
  VNStageIntLLRInputS0xD(76)(0) <= CNStageIntLLROutputS0xD(41)(1);
  VNStageIntLLRInputS0xD(140)(0) <= CNStageIntLLROutputS0xD(41)(2);
  VNStageIntLLRInputS0xD(204)(0) <= CNStageIntLLROutputS0xD(41)(3);
  VNStageIntLLRInputS0xD(268)(0) <= CNStageIntLLROutputS0xD(41)(4);
  VNStageIntLLRInputS0xD(332)(0) <= CNStageIntLLROutputS0xD(41)(5);
  VNStageIntLLRInputS0xD(11)(0) <= CNStageIntLLROutputS0xD(42)(0);
  VNStageIntLLRInputS0xD(75)(0) <= CNStageIntLLROutputS0xD(42)(1);
  VNStageIntLLRInputS0xD(139)(0) <= CNStageIntLLROutputS0xD(42)(2);
  VNStageIntLLRInputS0xD(203)(0) <= CNStageIntLLROutputS0xD(42)(3);
  VNStageIntLLRInputS0xD(267)(0) <= CNStageIntLLROutputS0xD(42)(4);
  VNStageIntLLRInputS0xD(331)(0) <= CNStageIntLLROutputS0xD(42)(5);
  VNStageIntLLRInputS0xD(10)(0) <= CNStageIntLLROutputS0xD(43)(0);
  VNStageIntLLRInputS0xD(74)(0) <= CNStageIntLLROutputS0xD(43)(1);
  VNStageIntLLRInputS0xD(138)(0) <= CNStageIntLLROutputS0xD(43)(2);
  VNStageIntLLRInputS0xD(202)(0) <= CNStageIntLLROutputS0xD(43)(3);
  VNStageIntLLRInputS0xD(266)(0) <= CNStageIntLLROutputS0xD(43)(4);
  VNStageIntLLRInputS0xD(330)(0) <= CNStageIntLLROutputS0xD(43)(5);
  VNStageIntLLRInputS0xD(9)(0) <= CNStageIntLLROutputS0xD(44)(0);
  VNStageIntLLRInputS0xD(73)(0) <= CNStageIntLLROutputS0xD(44)(1);
  VNStageIntLLRInputS0xD(137)(0) <= CNStageIntLLROutputS0xD(44)(2);
  VNStageIntLLRInputS0xD(201)(0) <= CNStageIntLLROutputS0xD(44)(3);
  VNStageIntLLRInputS0xD(265)(0) <= CNStageIntLLROutputS0xD(44)(4);
  VNStageIntLLRInputS0xD(329)(0) <= CNStageIntLLROutputS0xD(44)(5);
  VNStageIntLLRInputS0xD(8)(0) <= CNStageIntLLROutputS0xD(45)(0);
  VNStageIntLLRInputS0xD(72)(0) <= CNStageIntLLROutputS0xD(45)(1);
  VNStageIntLLRInputS0xD(136)(0) <= CNStageIntLLROutputS0xD(45)(2);
  VNStageIntLLRInputS0xD(200)(0) <= CNStageIntLLROutputS0xD(45)(3);
  VNStageIntLLRInputS0xD(264)(0) <= CNStageIntLLROutputS0xD(45)(4);
  VNStageIntLLRInputS0xD(328)(0) <= CNStageIntLLROutputS0xD(45)(5);
  VNStageIntLLRInputS0xD(7)(0) <= CNStageIntLLROutputS0xD(46)(0);
  VNStageIntLLRInputS0xD(71)(0) <= CNStageIntLLROutputS0xD(46)(1);
  VNStageIntLLRInputS0xD(135)(0) <= CNStageIntLLROutputS0xD(46)(2);
  VNStageIntLLRInputS0xD(199)(0) <= CNStageIntLLROutputS0xD(46)(3);
  VNStageIntLLRInputS0xD(263)(0) <= CNStageIntLLROutputS0xD(46)(4);
  VNStageIntLLRInputS0xD(327)(0) <= CNStageIntLLROutputS0xD(46)(5);
  VNStageIntLLRInputS0xD(6)(0) <= CNStageIntLLROutputS0xD(47)(0);
  VNStageIntLLRInputS0xD(70)(0) <= CNStageIntLLROutputS0xD(47)(1);
  VNStageIntLLRInputS0xD(134)(0) <= CNStageIntLLROutputS0xD(47)(2);
  VNStageIntLLRInputS0xD(198)(0) <= CNStageIntLLROutputS0xD(47)(3);
  VNStageIntLLRInputS0xD(262)(0) <= CNStageIntLLROutputS0xD(47)(4);
  VNStageIntLLRInputS0xD(326)(0) <= CNStageIntLLROutputS0xD(47)(5);
  VNStageIntLLRInputS0xD(5)(0) <= CNStageIntLLROutputS0xD(48)(0);
  VNStageIntLLRInputS0xD(69)(0) <= CNStageIntLLROutputS0xD(48)(1);
  VNStageIntLLRInputS0xD(133)(0) <= CNStageIntLLROutputS0xD(48)(2);
  VNStageIntLLRInputS0xD(197)(0) <= CNStageIntLLROutputS0xD(48)(3);
  VNStageIntLLRInputS0xD(261)(0) <= CNStageIntLLROutputS0xD(48)(4);
  VNStageIntLLRInputS0xD(325)(0) <= CNStageIntLLROutputS0xD(48)(5);
  VNStageIntLLRInputS0xD(4)(0) <= CNStageIntLLROutputS0xD(49)(0);
  VNStageIntLLRInputS0xD(68)(0) <= CNStageIntLLROutputS0xD(49)(1);
  VNStageIntLLRInputS0xD(132)(0) <= CNStageIntLLROutputS0xD(49)(2);
  VNStageIntLLRInputS0xD(196)(0) <= CNStageIntLLROutputS0xD(49)(3);
  VNStageIntLLRInputS0xD(260)(0) <= CNStageIntLLROutputS0xD(49)(4);
  VNStageIntLLRInputS0xD(324)(0) <= CNStageIntLLROutputS0xD(49)(5);
  VNStageIntLLRInputS0xD(2)(0) <= CNStageIntLLROutputS0xD(50)(0);
  VNStageIntLLRInputS0xD(66)(0) <= CNStageIntLLROutputS0xD(50)(1);
  VNStageIntLLRInputS0xD(130)(0) <= CNStageIntLLROutputS0xD(50)(2);
  VNStageIntLLRInputS0xD(194)(0) <= CNStageIntLLROutputS0xD(50)(3);
  VNStageIntLLRInputS0xD(258)(0) <= CNStageIntLLROutputS0xD(50)(4);
  VNStageIntLLRInputS0xD(322)(0) <= CNStageIntLLROutputS0xD(50)(5);
  VNStageIntLLRInputS0xD(1)(0) <= CNStageIntLLROutputS0xD(51)(0);
  VNStageIntLLRInputS0xD(65)(0) <= CNStageIntLLROutputS0xD(51)(1);
  VNStageIntLLRInputS0xD(129)(0) <= CNStageIntLLROutputS0xD(51)(2);
  VNStageIntLLRInputS0xD(193)(0) <= CNStageIntLLROutputS0xD(51)(3);
  VNStageIntLLRInputS0xD(257)(0) <= CNStageIntLLROutputS0xD(51)(4);
  VNStageIntLLRInputS0xD(321)(0) <= CNStageIntLLROutputS0xD(51)(5);
  VNStageIntLLRInputS0xD(63)(0) <= CNStageIntLLROutputS0xD(52)(0);
  VNStageIntLLRInputS0xD(127)(0) <= CNStageIntLLROutputS0xD(52)(1);
  VNStageIntLLRInputS0xD(191)(0) <= CNStageIntLLROutputS0xD(52)(2);
  VNStageIntLLRInputS0xD(255)(0) <= CNStageIntLLROutputS0xD(52)(3);
  VNStageIntLLRInputS0xD(319)(0) <= CNStageIntLLROutputS0xD(52)(4);
  VNStageIntLLRInputS0xD(383)(0) <= CNStageIntLLROutputS0xD(52)(5);
  VNStageIntLLRInputS0xD(0)(0) <= CNStageIntLLROutputS0xD(53)(0);
  VNStageIntLLRInputS0xD(64)(0) <= CNStageIntLLROutputS0xD(53)(1);
  VNStageIntLLRInputS0xD(128)(0) <= CNStageIntLLROutputS0xD(53)(2);
  VNStageIntLLRInputS0xD(192)(0) <= CNStageIntLLROutputS0xD(53)(3);
  VNStageIntLLRInputS0xD(256)(0) <= CNStageIntLLROutputS0xD(53)(4);
  VNStageIntLLRInputS0xD(320)(0) <= CNStageIntLLROutputS0xD(53)(5);
  VNStageIntLLRInputS0xD(42)(1) <= CNStageIntLLROutputS0xD(54)(0);
  VNStageIntLLRInputS0xD(112)(1) <= CNStageIntLLROutputS0xD(54)(1);
  VNStageIntLLRInputS0xD(182)(1) <= CNStageIntLLROutputS0xD(54)(2);
  VNStageIntLLRInputS0xD(203)(1) <= CNStageIntLLROutputS0xD(54)(3);
  VNStageIntLLRInputS0xD(259)(0) <= CNStageIntLLROutputS0xD(54)(4);
  VNStageIntLLRInputS0xD(361)(1) <= CNStageIntLLROutputS0xD(54)(5);
  VNStageIntLLRInputS0xD(41)(1) <= CNStageIntLLROutputS0xD(55)(0);
  VNStageIntLLRInputS0xD(117)(1) <= CNStageIntLLROutputS0xD(55)(1);
  VNStageIntLLRInputS0xD(138)(1) <= CNStageIntLLROutputS0xD(55)(2);
  VNStageIntLLRInputS0xD(194)(1) <= CNStageIntLLROutputS0xD(55)(3);
  VNStageIntLLRInputS0xD(296)(1) <= CNStageIntLLROutputS0xD(55)(4);
  VNStageIntLLRInputS0xD(362)(1) <= CNStageIntLLROutputS0xD(55)(5);
  VNStageIntLLRInputS0xD(40)(1) <= CNStageIntLLROutputS0xD(56)(0);
  VNStageIntLLRInputS0xD(73)(1) <= CNStageIntLLROutputS0xD(56)(1);
  VNStageIntLLRInputS0xD(129)(1) <= CNStageIntLLROutputS0xD(56)(2);
  VNStageIntLLRInputS0xD(231)(1) <= CNStageIntLLROutputS0xD(56)(3);
  VNStageIntLLRInputS0xD(297)(1) <= CNStageIntLLROutputS0xD(56)(4);
  VNStageIntLLRInputS0xD(323)(0) <= CNStageIntLLROutputS0xD(56)(5);
  VNStageIntLLRInputS0xD(39)(1) <= CNStageIntLLROutputS0xD(57)(0);
  VNStageIntLLRInputS0xD(127)(1) <= CNStageIntLLROutputS0xD(57)(1);
  VNStageIntLLRInputS0xD(166)(1) <= CNStageIntLLROutputS0xD(57)(2);
  VNStageIntLLRInputS0xD(232)(1) <= CNStageIntLLROutputS0xD(57)(3);
  VNStageIntLLRInputS0xD(258)(1) <= CNStageIntLLROutputS0xD(57)(4);
  VNStageIntLLRInputS0xD(344)(1) <= CNStageIntLLROutputS0xD(57)(5);
  VNStageIntLLRInputS0xD(38)(1) <= CNStageIntLLROutputS0xD(58)(0);
  VNStageIntLLRInputS0xD(101)(1) <= CNStageIntLLROutputS0xD(58)(1);
  VNStageIntLLRInputS0xD(167)(1) <= CNStageIntLLROutputS0xD(58)(2);
  VNStageIntLLRInputS0xD(193)(1) <= CNStageIntLLROutputS0xD(58)(3);
  VNStageIntLLRInputS0xD(279)(1) <= CNStageIntLLROutputS0xD(58)(4);
  VNStageIntLLRInputS0xD(340)(1) <= CNStageIntLLROutputS0xD(58)(5);
  VNStageIntLLRInputS0xD(37)(1) <= CNStageIntLLROutputS0xD(59)(0);
  VNStageIntLLRInputS0xD(102)(1) <= CNStageIntLLROutputS0xD(59)(1);
  VNStageIntLLRInputS0xD(191)(1) <= CNStageIntLLROutputS0xD(59)(2);
  VNStageIntLLRInputS0xD(214)(1) <= CNStageIntLLROutputS0xD(59)(3);
  VNStageIntLLRInputS0xD(275)(1) <= CNStageIntLLROutputS0xD(59)(4);
  VNStageIntLLRInputS0xD(355)(1) <= CNStageIntLLROutputS0xD(59)(5);
  VNStageIntLLRInputS0xD(36)(1) <= CNStageIntLLROutputS0xD(60)(0);
  VNStageIntLLRInputS0xD(126)(0) <= CNStageIntLLROutputS0xD(60)(1);
  VNStageIntLLRInputS0xD(149)(1) <= CNStageIntLLROutputS0xD(60)(2);
  VNStageIntLLRInputS0xD(210)(1) <= CNStageIntLLROutputS0xD(60)(3);
  VNStageIntLLRInputS0xD(290)(1) <= CNStageIntLLROutputS0xD(60)(4);
  VNStageIntLLRInputS0xD(381)(0) <= CNStageIntLLROutputS0xD(60)(5);
  VNStageIntLLRInputS0xD(35)(1) <= CNStageIntLLROutputS0xD(61)(0);
  VNStageIntLLRInputS0xD(84)(1) <= CNStageIntLLROutputS0xD(61)(1);
  VNStageIntLLRInputS0xD(145)(1) <= CNStageIntLLROutputS0xD(61)(2);
  VNStageIntLLRInputS0xD(225)(1) <= CNStageIntLLROutputS0xD(61)(3);
  VNStageIntLLRInputS0xD(316)(0) <= CNStageIntLLROutputS0xD(61)(4);
  VNStageIntLLRInputS0xD(357)(1) <= CNStageIntLLROutputS0xD(61)(5);
  VNStageIntLLRInputS0xD(34)(1) <= CNStageIntLLROutputS0xD(62)(0);
  VNStageIntLLRInputS0xD(80)(1) <= CNStageIntLLROutputS0xD(62)(1);
  VNStageIntLLRInputS0xD(160)(1) <= CNStageIntLLROutputS0xD(62)(2);
  VNStageIntLLRInputS0xD(251)(0) <= CNStageIntLLROutputS0xD(62)(3);
  VNStageIntLLRInputS0xD(292)(1) <= CNStageIntLLROutputS0xD(62)(4);
  VNStageIntLLRInputS0xD(326)(1) <= CNStageIntLLROutputS0xD(62)(5);
  VNStageIntLLRInputS0xD(33)(1) <= CNStageIntLLROutputS0xD(63)(0);
  VNStageIntLLRInputS0xD(95)(1) <= CNStageIntLLROutputS0xD(63)(1);
  VNStageIntLLRInputS0xD(186)(0) <= CNStageIntLLROutputS0xD(63)(2);
  VNStageIntLLRInputS0xD(227)(1) <= CNStageIntLLROutputS0xD(63)(3);
  VNStageIntLLRInputS0xD(261)(1) <= CNStageIntLLROutputS0xD(63)(4);
  VNStageIntLLRInputS0xD(342)(1) <= CNStageIntLLROutputS0xD(63)(5);
  VNStageIntLLRInputS0xD(32)(1) <= CNStageIntLLROutputS0xD(64)(0);
  VNStageIntLLRInputS0xD(121)(0) <= CNStageIntLLROutputS0xD(64)(1);
  VNStageIntLLRInputS0xD(162)(1) <= CNStageIntLLROutputS0xD(64)(2);
  VNStageIntLLRInputS0xD(196)(1) <= CNStageIntLLROutputS0xD(64)(3);
  VNStageIntLLRInputS0xD(277)(1) <= CNStageIntLLROutputS0xD(64)(4);
  VNStageIntLLRInputS0xD(375)(1) <= CNStageIntLLROutputS0xD(64)(5);
  VNStageIntLLRInputS0xD(31)(1) <= CNStageIntLLROutputS0xD(65)(0);
  VNStageIntLLRInputS0xD(97)(1) <= CNStageIntLLROutputS0xD(65)(1);
  VNStageIntLLRInputS0xD(131)(0) <= CNStageIntLLROutputS0xD(65)(2);
  VNStageIntLLRInputS0xD(212)(1) <= CNStageIntLLROutputS0xD(65)(3);
  VNStageIntLLRInputS0xD(310)(1) <= CNStageIntLLROutputS0xD(65)(4);
  VNStageIntLLRInputS0xD(321)(1) <= CNStageIntLLROutputS0xD(65)(5);
  VNStageIntLLRInputS0xD(30)(1) <= CNStageIntLLROutputS0xD(66)(0);
  VNStageIntLLRInputS0xD(66)(1) <= CNStageIntLLROutputS0xD(66)(1);
  VNStageIntLLRInputS0xD(147)(1) <= CNStageIntLLROutputS0xD(66)(2);
  VNStageIntLLRInputS0xD(245)(1) <= CNStageIntLLROutputS0xD(66)(3);
  VNStageIntLLRInputS0xD(319)(1) <= CNStageIntLLROutputS0xD(66)(4);
  VNStageIntLLRInputS0xD(334)(1) <= CNStageIntLLROutputS0xD(66)(5);
  VNStageIntLLRInputS0xD(29)(1) <= CNStageIntLLROutputS0xD(67)(0);
  VNStageIntLLRInputS0xD(82)(1) <= CNStageIntLLROutputS0xD(67)(1);
  VNStageIntLLRInputS0xD(180)(0) <= CNStageIntLLROutputS0xD(67)(2);
  VNStageIntLLRInputS0xD(254)(0) <= CNStageIntLLROutputS0xD(67)(3);
  VNStageIntLLRInputS0xD(269)(0) <= CNStageIntLLROutputS0xD(67)(4);
  VNStageIntLLRInputS0xD(376)(1) <= CNStageIntLLROutputS0xD(67)(5);
  VNStageIntLLRInputS0xD(28)(1) <= CNStageIntLLROutputS0xD(68)(0);
  VNStageIntLLRInputS0xD(115)(1) <= CNStageIntLLROutputS0xD(68)(1);
  VNStageIntLLRInputS0xD(189)(0) <= CNStageIntLLROutputS0xD(68)(2);
  VNStageIntLLRInputS0xD(204)(1) <= CNStageIntLLROutputS0xD(68)(3);
  VNStageIntLLRInputS0xD(311)(1) <= CNStageIntLLROutputS0xD(68)(4);
  VNStageIntLLRInputS0xD(341)(1) <= CNStageIntLLROutputS0xD(68)(5);
  VNStageIntLLRInputS0xD(27)(1) <= CNStageIntLLROutputS0xD(69)(0);
  VNStageIntLLRInputS0xD(124)(0) <= CNStageIntLLROutputS0xD(69)(1);
  VNStageIntLLRInputS0xD(139)(1) <= CNStageIntLLROutputS0xD(69)(2);
  VNStageIntLLRInputS0xD(246)(1) <= CNStageIntLLROutputS0xD(69)(3);
  VNStageIntLLRInputS0xD(276)(1) <= CNStageIntLLROutputS0xD(69)(4);
  VNStageIntLLRInputS0xD(343)(1) <= CNStageIntLLROutputS0xD(69)(5);
  VNStageIntLLRInputS0xD(26)(1) <= CNStageIntLLROutputS0xD(70)(0);
  VNStageIntLLRInputS0xD(74)(1) <= CNStageIntLLROutputS0xD(70)(1);
  VNStageIntLLRInputS0xD(181)(1) <= CNStageIntLLROutputS0xD(70)(2);
  VNStageIntLLRInputS0xD(211)(1) <= CNStageIntLLROutputS0xD(70)(3);
  VNStageIntLLRInputS0xD(278)(1) <= CNStageIntLLROutputS0xD(70)(4);
  VNStageIntLLRInputS0xD(325)(1) <= CNStageIntLLROutputS0xD(70)(5);
  VNStageIntLLRInputS0xD(25)(1) <= CNStageIntLLROutputS0xD(71)(0);
  VNStageIntLLRInputS0xD(116)(0) <= CNStageIntLLROutputS0xD(71)(1);
  VNStageIntLLRInputS0xD(146)(1) <= CNStageIntLLROutputS0xD(71)(2);
  VNStageIntLLRInputS0xD(213)(1) <= CNStageIntLLROutputS0xD(71)(3);
  VNStageIntLLRInputS0xD(260)(1) <= CNStageIntLLROutputS0xD(71)(4);
  VNStageIntLLRInputS0xD(332)(1) <= CNStageIntLLROutputS0xD(71)(5);
  VNStageIntLLRInputS0xD(24)(1) <= CNStageIntLLROutputS0xD(72)(0);
  VNStageIntLLRInputS0xD(81)(1) <= CNStageIntLLROutputS0xD(72)(1);
  VNStageIntLLRInputS0xD(148)(1) <= CNStageIntLLROutputS0xD(72)(2);
  VNStageIntLLRInputS0xD(195)(0) <= CNStageIntLLROutputS0xD(72)(3);
  VNStageIntLLRInputS0xD(267)(1) <= CNStageIntLLROutputS0xD(72)(4);
  VNStageIntLLRInputS0xD(359)(1) <= CNStageIntLLROutputS0xD(72)(5);
  VNStageIntLLRInputS0xD(23)(1) <= CNStageIntLLROutputS0xD(73)(0);
  VNStageIntLLRInputS0xD(83)(1) <= CNStageIntLLROutputS0xD(73)(1);
  VNStageIntLLRInputS0xD(130)(1) <= CNStageIntLLROutputS0xD(73)(2);
  VNStageIntLLRInputS0xD(202)(1) <= CNStageIntLLROutputS0xD(73)(3);
  VNStageIntLLRInputS0xD(294)(1) <= CNStageIntLLROutputS0xD(73)(4);
  VNStageIntLLRInputS0xD(347)(1) <= CNStageIntLLROutputS0xD(73)(5);
  VNStageIntLLRInputS0xD(22)(1) <= CNStageIntLLROutputS0xD(74)(0);
  VNStageIntLLRInputS0xD(65)(1) <= CNStageIntLLROutputS0xD(74)(1);
  VNStageIntLLRInputS0xD(137)(1) <= CNStageIntLLROutputS0xD(74)(2);
  VNStageIntLLRInputS0xD(229)(1) <= CNStageIntLLROutputS0xD(74)(3);
  VNStageIntLLRInputS0xD(282)(1) <= CNStageIntLLROutputS0xD(74)(4);
  VNStageIntLLRInputS0xD(353)(1) <= CNStageIntLLROutputS0xD(74)(5);
  VNStageIntLLRInputS0xD(21)(1) <= CNStageIntLLROutputS0xD(75)(0);
  VNStageIntLLRInputS0xD(72)(1) <= CNStageIntLLROutputS0xD(75)(1);
  VNStageIntLLRInputS0xD(164)(1) <= CNStageIntLLROutputS0xD(75)(2);
  VNStageIntLLRInputS0xD(217)(1) <= CNStageIntLLROutputS0xD(75)(3);
  VNStageIntLLRInputS0xD(288)(1) <= CNStageIntLLROutputS0xD(75)(4);
  VNStageIntLLRInputS0xD(348)(1) <= CNStageIntLLROutputS0xD(75)(5);
  VNStageIntLLRInputS0xD(20)(1) <= CNStageIntLLROutputS0xD(76)(0);
  VNStageIntLLRInputS0xD(99)(1) <= CNStageIntLLROutputS0xD(76)(1);
  VNStageIntLLRInputS0xD(152)(1) <= CNStageIntLLROutputS0xD(76)(2);
  VNStageIntLLRInputS0xD(223)(1) <= CNStageIntLLROutputS0xD(76)(3);
  VNStageIntLLRInputS0xD(283)(1) <= CNStageIntLLROutputS0xD(76)(4);
  VNStageIntLLRInputS0xD(358)(1) <= CNStageIntLLROutputS0xD(76)(5);
  VNStageIntLLRInputS0xD(19)(1) <= CNStageIntLLROutputS0xD(77)(0);
  VNStageIntLLRInputS0xD(87)(1) <= CNStageIntLLROutputS0xD(77)(1);
  VNStageIntLLRInputS0xD(158)(1) <= CNStageIntLLROutputS0xD(77)(2);
  VNStageIntLLRInputS0xD(218)(1) <= CNStageIntLLROutputS0xD(77)(3);
  VNStageIntLLRInputS0xD(293)(1) <= CNStageIntLLROutputS0xD(77)(4);
  VNStageIntLLRInputS0xD(380)(0) <= CNStageIntLLROutputS0xD(77)(5);
  VNStageIntLLRInputS0xD(18)(1) <= CNStageIntLLROutputS0xD(78)(0);
  VNStageIntLLRInputS0xD(93)(1) <= CNStageIntLLROutputS0xD(78)(1);
  VNStageIntLLRInputS0xD(153)(1) <= CNStageIntLLROutputS0xD(78)(2);
  VNStageIntLLRInputS0xD(228)(1) <= CNStageIntLLROutputS0xD(78)(3);
  VNStageIntLLRInputS0xD(315)(0) <= CNStageIntLLROutputS0xD(78)(4);
  VNStageIntLLRInputS0xD(335)(1) <= CNStageIntLLROutputS0xD(78)(5);
  VNStageIntLLRInputS0xD(17)(1) <= CNStageIntLLROutputS0xD(79)(0);
  VNStageIntLLRInputS0xD(88)(1) <= CNStageIntLLROutputS0xD(79)(1);
  VNStageIntLLRInputS0xD(163)(1) <= CNStageIntLLROutputS0xD(79)(2);
  VNStageIntLLRInputS0xD(250)(0) <= CNStageIntLLROutputS0xD(79)(3);
  VNStageIntLLRInputS0xD(270)(1) <= CNStageIntLLROutputS0xD(79)(4);
  VNStageIntLLRInputS0xD(383)(1) <= CNStageIntLLROutputS0xD(79)(5);
  VNStageIntLLRInputS0xD(15)(1) <= CNStageIntLLROutputS0xD(80)(0);
  VNStageIntLLRInputS0xD(120)(1) <= CNStageIntLLROutputS0xD(80)(1);
  VNStageIntLLRInputS0xD(140)(1) <= CNStageIntLLROutputS0xD(80)(2);
  VNStageIntLLRInputS0xD(253)(0) <= CNStageIntLLROutputS0xD(80)(3);
  VNStageIntLLRInputS0xD(305)(1) <= CNStageIntLLROutputS0xD(80)(4);
  VNStageIntLLRInputS0xD(338)(1) <= CNStageIntLLROutputS0xD(80)(5);
  VNStageIntLLRInputS0xD(14)(1) <= CNStageIntLLROutputS0xD(81)(0);
  VNStageIntLLRInputS0xD(75)(1) <= CNStageIntLLROutputS0xD(81)(1);
  VNStageIntLLRInputS0xD(188)(0) <= CNStageIntLLROutputS0xD(81)(2);
  VNStageIntLLRInputS0xD(240)(1) <= CNStageIntLLROutputS0xD(81)(3);
  VNStageIntLLRInputS0xD(273)(1) <= CNStageIntLLROutputS0xD(81)(4);
  VNStageIntLLRInputS0xD(350)(1) <= CNStageIntLLROutputS0xD(81)(5);
  VNStageIntLLRInputS0xD(13)(0) <= CNStageIntLLROutputS0xD(82)(0);
  VNStageIntLLRInputS0xD(123)(0) <= CNStageIntLLROutputS0xD(82)(1);
  VNStageIntLLRInputS0xD(175)(1) <= CNStageIntLLROutputS0xD(82)(2);
  VNStageIntLLRInputS0xD(208)(1) <= CNStageIntLLROutputS0xD(82)(3);
  VNStageIntLLRInputS0xD(285)(1) <= CNStageIntLLROutputS0xD(82)(4);
  VNStageIntLLRInputS0xD(364)(1) <= CNStageIntLLROutputS0xD(82)(5);
  VNStageIntLLRInputS0xD(12)(1) <= CNStageIntLLROutputS0xD(83)(0);
  VNStageIntLLRInputS0xD(110)(1) <= CNStageIntLLROutputS0xD(83)(1);
  VNStageIntLLRInputS0xD(143)(1) <= CNStageIntLLROutputS0xD(83)(2);
  VNStageIntLLRInputS0xD(220)(1) <= CNStageIntLLROutputS0xD(83)(3);
  VNStageIntLLRInputS0xD(299)(0) <= CNStageIntLLROutputS0xD(83)(4);
  VNStageIntLLRInputS0xD(345)(1) <= CNStageIntLLROutputS0xD(83)(5);
  VNStageIntLLRInputS0xD(11)(1) <= CNStageIntLLROutputS0xD(84)(0);
  VNStageIntLLRInputS0xD(78)(1) <= CNStageIntLLROutputS0xD(84)(1);
  VNStageIntLLRInputS0xD(155)(1) <= CNStageIntLLROutputS0xD(84)(2);
  VNStageIntLLRInputS0xD(234)(1) <= CNStageIntLLROutputS0xD(84)(3);
  VNStageIntLLRInputS0xD(280)(1) <= CNStageIntLLROutputS0xD(84)(4);
  VNStageIntLLRInputS0xD(322)(1) <= CNStageIntLLROutputS0xD(84)(5);
  VNStageIntLLRInputS0xD(10)(1) <= CNStageIntLLROutputS0xD(85)(0);
  VNStageIntLLRInputS0xD(90)(1) <= CNStageIntLLROutputS0xD(85)(1);
  VNStageIntLLRInputS0xD(169)(1) <= CNStageIntLLROutputS0xD(85)(2);
  VNStageIntLLRInputS0xD(215)(1) <= CNStageIntLLROutputS0xD(85)(3);
  VNStageIntLLRInputS0xD(257)(1) <= CNStageIntLLROutputS0xD(85)(4);
  VNStageIntLLRInputS0xD(374)(1) <= CNStageIntLLROutputS0xD(85)(5);
  VNStageIntLLRInputS0xD(9)(1) <= CNStageIntLLROutputS0xD(86)(0);
  VNStageIntLLRInputS0xD(104)(1) <= CNStageIntLLROutputS0xD(86)(1);
  VNStageIntLLRInputS0xD(150)(1) <= CNStageIntLLROutputS0xD(86)(2);
  VNStageIntLLRInputS0xD(255)(1) <= CNStageIntLLROutputS0xD(86)(3);
  VNStageIntLLRInputS0xD(309)(1) <= CNStageIntLLROutputS0xD(86)(4);
  VNStageIntLLRInputS0xD(378)(0) <= CNStageIntLLROutputS0xD(86)(5);
  VNStageIntLLRInputS0xD(7)(1) <= CNStageIntLLROutputS0xD(87)(0);
  VNStageIntLLRInputS0xD(125)(0) <= CNStageIntLLROutputS0xD(87)(1);
  VNStageIntLLRInputS0xD(179)(1) <= CNStageIntLLROutputS0xD(87)(2);
  VNStageIntLLRInputS0xD(248)(1) <= CNStageIntLLROutputS0xD(87)(3);
  VNStageIntLLRInputS0xD(306)(1) <= CNStageIntLLROutputS0xD(87)(4);
  VNStageIntLLRInputS0xD(382)(0) <= CNStageIntLLROutputS0xD(87)(5);
  VNStageIntLLRInputS0xD(6)(1) <= CNStageIntLLROutputS0xD(88)(0);
  VNStageIntLLRInputS0xD(114)(1) <= CNStageIntLLROutputS0xD(88)(1);
  VNStageIntLLRInputS0xD(183)(1) <= CNStageIntLLROutputS0xD(88)(2);
  VNStageIntLLRInputS0xD(241)(1) <= CNStageIntLLROutputS0xD(88)(3);
  VNStageIntLLRInputS0xD(317)(0) <= CNStageIntLLROutputS0xD(88)(4);
  VNStageIntLLRInputS0xD(354)(1) <= CNStageIntLLROutputS0xD(88)(5);
  VNStageIntLLRInputS0xD(5)(1) <= CNStageIntLLROutputS0xD(89)(0);
  VNStageIntLLRInputS0xD(118)(1) <= CNStageIntLLROutputS0xD(89)(1);
  VNStageIntLLRInputS0xD(176)(1) <= CNStageIntLLROutputS0xD(89)(2);
  VNStageIntLLRInputS0xD(252)(0) <= CNStageIntLLROutputS0xD(89)(3);
  VNStageIntLLRInputS0xD(289)(1) <= CNStageIntLLROutputS0xD(89)(4);
  VNStageIntLLRInputS0xD(346)(1) <= CNStageIntLLROutputS0xD(89)(5);
  VNStageIntLLRInputS0xD(4)(1) <= CNStageIntLLROutputS0xD(90)(0);
  VNStageIntLLRInputS0xD(111)(1) <= CNStageIntLLROutputS0xD(90)(1);
  VNStageIntLLRInputS0xD(187)(0) <= CNStageIntLLROutputS0xD(90)(2);
  VNStageIntLLRInputS0xD(224)(1) <= CNStageIntLLROutputS0xD(90)(3);
  VNStageIntLLRInputS0xD(281)(1) <= CNStageIntLLROutputS0xD(90)(4);
  VNStageIntLLRInputS0xD(363)(0) <= CNStageIntLLROutputS0xD(90)(5);
  VNStageIntLLRInputS0xD(3)(0) <= CNStageIntLLROutputS0xD(91)(0);
  VNStageIntLLRInputS0xD(122)(0) <= CNStageIntLLROutputS0xD(91)(1);
  VNStageIntLLRInputS0xD(159)(1) <= CNStageIntLLROutputS0xD(91)(2);
  VNStageIntLLRInputS0xD(216)(1) <= CNStageIntLLROutputS0xD(91)(3);
  VNStageIntLLRInputS0xD(298)(1) <= CNStageIntLLROutputS0xD(91)(4);
  VNStageIntLLRInputS0xD(360)(1) <= CNStageIntLLROutputS0xD(91)(5);
  VNStageIntLLRInputS0xD(2)(1) <= CNStageIntLLROutputS0xD(92)(0);
  VNStageIntLLRInputS0xD(94)(1) <= CNStageIntLLROutputS0xD(92)(1);
  VNStageIntLLRInputS0xD(151)(1) <= CNStageIntLLROutputS0xD(92)(2);
  VNStageIntLLRInputS0xD(233)(1) <= CNStageIntLLROutputS0xD(92)(3);
  VNStageIntLLRInputS0xD(295)(1) <= CNStageIntLLROutputS0xD(92)(4);
  VNStageIntLLRInputS0xD(331)(1) <= CNStageIntLLROutputS0xD(92)(5);
  VNStageIntLLRInputS0xD(63)(1) <= CNStageIntLLROutputS0xD(93)(0);
  VNStageIntLLRInputS0xD(103)(1) <= CNStageIntLLROutputS0xD(93)(1);
  VNStageIntLLRInputS0xD(165)(1) <= CNStageIntLLROutputS0xD(93)(2);
  VNStageIntLLRInputS0xD(201)(1) <= CNStageIntLLROutputS0xD(93)(3);
  VNStageIntLLRInputS0xD(286)(1) <= CNStageIntLLROutputS0xD(93)(4);
  VNStageIntLLRInputS0xD(337)(1) <= CNStageIntLLROutputS0xD(93)(5);
  VNStageIntLLRInputS0xD(62)(0) <= CNStageIntLLROutputS0xD(94)(0);
  VNStageIntLLRInputS0xD(100)(1) <= CNStageIntLLROutputS0xD(94)(1);
  VNStageIntLLRInputS0xD(136)(1) <= CNStageIntLLROutputS0xD(94)(2);
  VNStageIntLLRInputS0xD(221)(1) <= CNStageIntLLROutputS0xD(94)(3);
  VNStageIntLLRInputS0xD(272)(1) <= CNStageIntLLROutputS0xD(94)(4);
  VNStageIntLLRInputS0xD(327)(1) <= CNStageIntLLROutputS0xD(94)(5);
  VNStageIntLLRInputS0xD(61)(0) <= CNStageIntLLROutputS0xD(95)(0);
  VNStageIntLLRInputS0xD(71)(1) <= CNStageIntLLROutputS0xD(95)(1);
  VNStageIntLLRInputS0xD(156)(1) <= CNStageIntLLROutputS0xD(95)(2);
  VNStageIntLLRInputS0xD(207)(1) <= CNStageIntLLROutputS0xD(95)(3);
  VNStageIntLLRInputS0xD(262)(1) <= CNStageIntLLROutputS0xD(95)(4);
  VNStageIntLLRInputS0xD(356)(1) <= CNStageIntLLROutputS0xD(95)(5);
  VNStageIntLLRInputS0xD(60)(0) <= CNStageIntLLROutputS0xD(96)(0);
  VNStageIntLLRInputS0xD(91)(1) <= CNStageIntLLROutputS0xD(96)(1);
  VNStageIntLLRInputS0xD(142)(1) <= CNStageIntLLROutputS0xD(96)(2);
  VNStageIntLLRInputS0xD(197)(1) <= CNStageIntLLROutputS0xD(96)(3);
  VNStageIntLLRInputS0xD(291)(1) <= CNStageIntLLROutputS0xD(96)(4);
  VNStageIntLLRInputS0xD(339)(1) <= CNStageIntLLROutputS0xD(96)(5);
  VNStageIntLLRInputS0xD(58)(0) <= CNStageIntLLROutputS0xD(97)(0);
  VNStageIntLLRInputS0xD(67)(0) <= CNStageIntLLROutputS0xD(97)(1);
  VNStageIntLLRInputS0xD(161)(1) <= CNStageIntLLROutputS0xD(97)(2);
  VNStageIntLLRInputS0xD(209)(1) <= CNStageIntLLROutputS0xD(97)(3);
  VNStageIntLLRInputS0xD(304)(1) <= CNStageIntLLROutputS0xD(97)(4);
  VNStageIntLLRInputS0xD(329)(1) <= CNStageIntLLROutputS0xD(97)(5);
  VNStageIntLLRInputS0xD(57)(0) <= CNStageIntLLROutputS0xD(98)(0);
  VNStageIntLLRInputS0xD(96)(1) <= CNStageIntLLROutputS0xD(98)(1);
  VNStageIntLLRInputS0xD(144)(1) <= CNStageIntLLROutputS0xD(98)(2);
  VNStageIntLLRInputS0xD(239)(1) <= CNStageIntLLROutputS0xD(98)(3);
  VNStageIntLLRInputS0xD(264)(1) <= CNStageIntLLROutputS0xD(98)(4);
  VNStageIntLLRInputS0xD(365)(1) <= CNStageIntLLROutputS0xD(98)(5);
  VNStageIntLLRInputS0xD(56)(1) <= CNStageIntLLROutputS0xD(99)(0);
  VNStageIntLLRInputS0xD(79)(1) <= CNStageIntLLROutputS0xD(99)(1);
  VNStageIntLLRInputS0xD(174)(1) <= CNStageIntLLROutputS0xD(99)(2);
  VNStageIntLLRInputS0xD(199)(1) <= CNStageIntLLROutputS0xD(99)(3);
  VNStageIntLLRInputS0xD(300)(1) <= CNStageIntLLROutputS0xD(99)(4);
  VNStageIntLLRInputS0xD(349)(1) <= CNStageIntLLROutputS0xD(99)(5);
  VNStageIntLLRInputS0xD(55)(1) <= CNStageIntLLROutputS0xD(100)(0);
  VNStageIntLLRInputS0xD(109)(1) <= CNStageIntLLROutputS0xD(100)(1);
  VNStageIntLLRInputS0xD(134)(1) <= CNStageIntLLROutputS0xD(100)(2);
  VNStageIntLLRInputS0xD(235)(0) <= CNStageIntLLROutputS0xD(100)(3);
  VNStageIntLLRInputS0xD(284)(1) <= CNStageIntLLROutputS0xD(100)(4);
  VNStageIntLLRInputS0xD(352)(1) <= CNStageIntLLROutputS0xD(100)(5);
  VNStageIntLLRInputS0xD(54)(1) <= CNStageIntLLROutputS0xD(101)(0);
  VNStageIntLLRInputS0xD(69)(1) <= CNStageIntLLROutputS0xD(101)(1);
  VNStageIntLLRInputS0xD(170)(1) <= CNStageIntLLROutputS0xD(101)(2);
  VNStageIntLLRInputS0xD(219)(1) <= CNStageIntLLROutputS0xD(101)(3);
  VNStageIntLLRInputS0xD(287)(1) <= CNStageIntLLROutputS0xD(101)(4);
  VNStageIntLLRInputS0xD(330)(1) <= CNStageIntLLROutputS0xD(101)(5);
  VNStageIntLLRInputS0xD(52)(0) <= CNStageIntLLROutputS0xD(102)(0);
  VNStageIntLLRInputS0xD(89)(1) <= CNStageIntLLROutputS0xD(102)(1);
  VNStageIntLLRInputS0xD(157)(1) <= CNStageIntLLROutputS0xD(102)(2);
  VNStageIntLLRInputS0xD(200)(1) <= CNStageIntLLROutputS0xD(102)(3);
  VNStageIntLLRInputS0xD(303)(1) <= CNStageIntLLROutputS0xD(102)(4);
  VNStageIntLLRInputS0xD(366)(1) <= CNStageIntLLROutputS0xD(102)(5);
  VNStageIntLLRInputS0xD(51)(1) <= CNStageIntLLROutputS0xD(103)(0);
  VNStageIntLLRInputS0xD(92)(1) <= CNStageIntLLROutputS0xD(103)(1);
  VNStageIntLLRInputS0xD(135)(1) <= CNStageIntLLROutputS0xD(103)(2);
  VNStageIntLLRInputS0xD(238)(1) <= CNStageIntLLROutputS0xD(103)(3);
  VNStageIntLLRInputS0xD(301)(1) <= CNStageIntLLROutputS0xD(103)(4);
  VNStageIntLLRInputS0xD(328)(1) <= CNStageIntLLROutputS0xD(103)(5);
  VNStageIntLLRInputS0xD(50)(1) <= CNStageIntLLROutputS0xD(104)(0);
  VNStageIntLLRInputS0xD(70)(1) <= CNStageIntLLROutputS0xD(104)(1);
  VNStageIntLLRInputS0xD(173)(1) <= CNStageIntLLROutputS0xD(104)(2);
  VNStageIntLLRInputS0xD(236)(1) <= CNStageIntLLROutputS0xD(104)(3);
  VNStageIntLLRInputS0xD(263)(1) <= CNStageIntLLROutputS0xD(104)(4);
  VNStageIntLLRInputS0xD(336)(1) <= CNStageIntLLROutputS0xD(104)(5);
  VNStageIntLLRInputS0xD(49)(1) <= CNStageIntLLROutputS0xD(105)(0);
  VNStageIntLLRInputS0xD(108)(1) <= CNStageIntLLROutputS0xD(105)(1);
  VNStageIntLLRInputS0xD(171)(0) <= CNStageIntLLROutputS0xD(105)(2);
  VNStageIntLLRInputS0xD(198)(1) <= CNStageIntLLROutputS0xD(105)(3);
  VNStageIntLLRInputS0xD(271)(1) <= CNStageIntLLROutputS0xD(105)(4);
  VNStageIntLLRInputS0xD(379)(0) <= CNStageIntLLROutputS0xD(105)(5);
  VNStageIntLLRInputS0xD(46)(1) <= CNStageIntLLROutputS0xD(106)(0);
  VNStageIntLLRInputS0xD(76)(1) <= CNStageIntLLROutputS0xD(106)(1);
  VNStageIntLLRInputS0xD(184)(1) <= CNStageIntLLROutputS0xD(106)(2);
  VNStageIntLLRInputS0xD(243)(1) <= CNStageIntLLROutputS0xD(106)(3);
  VNStageIntLLRInputS0xD(256)(1) <= CNStageIntLLROutputS0xD(106)(4);
  VNStageIntLLRInputS0xD(372)(0) <= CNStageIntLLROutputS0xD(106)(5);
  VNStageIntLLRInputS0xD(45)(1) <= CNStageIntLLROutputS0xD(107)(0);
  VNStageIntLLRInputS0xD(119)(1) <= CNStageIntLLROutputS0xD(107)(1);
  VNStageIntLLRInputS0xD(178)(1) <= CNStageIntLLROutputS0xD(107)(2);
  VNStageIntLLRInputS0xD(192)(1) <= CNStageIntLLROutputS0xD(107)(3);
  VNStageIntLLRInputS0xD(307)(1) <= CNStageIntLLROutputS0xD(107)(4);
  VNStageIntLLRInputS0xD(377)(0) <= CNStageIntLLROutputS0xD(107)(5);
  VNStageIntLLRInputS0xD(44)(1) <= CNStageIntLLROutputS0xD(108)(0);
  VNStageIntLLRInputS0xD(113)(1) <= CNStageIntLLROutputS0xD(108)(1);
  VNStageIntLLRInputS0xD(128)(1) <= CNStageIntLLROutputS0xD(108)(2);
  VNStageIntLLRInputS0xD(242)(1) <= CNStageIntLLROutputS0xD(108)(3);
  VNStageIntLLRInputS0xD(312)(1) <= CNStageIntLLROutputS0xD(108)(4);
  VNStageIntLLRInputS0xD(333)(0) <= CNStageIntLLROutputS0xD(108)(5);
  VNStageIntLLRInputS0xD(43)(0) <= CNStageIntLLROutputS0xD(109)(0);
  VNStageIntLLRInputS0xD(64)(1) <= CNStageIntLLROutputS0xD(109)(1);
  VNStageIntLLRInputS0xD(177)(1) <= CNStageIntLLROutputS0xD(109)(2);
  VNStageIntLLRInputS0xD(247)(1) <= CNStageIntLLROutputS0xD(109)(3);
  VNStageIntLLRInputS0xD(268)(1) <= CNStageIntLLROutputS0xD(109)(4);
  VNStageIntLLRInputS0xD(324)(1) <= CNStageIntLLROutputS0xD(109)(5);
  VNStageIntLLRInputS0xD(0)(1) <= CNStageIntLLROutputS0xD(110)(0);
  VNStageIntLLRInputS0xD(107)(0) <= CNStageIntLLROutputS0xD(110)(1);
  VNStageIntLLRInputS0xD(172)(1) <= CNStageIntLLROutputS0xD(110)(2);
  VNStageIntLLRInputS0xD(237)(1) <= CNStageIntLLROutputS0xD(110)(3);
  VNStageIntLLRInputS0xD(302)(1) <= CNStageIntLLROutputS0xD(110)(4);
  VNStageIntLLRInputS0xD(367)(1) <= CNStageIntLLROutputS0xD(110)(5);
  VNStageIntLLRInputS0xD(32)(2) <= CNStageIntLLROutputS0xD(111)(0);
  VNStageIntLLRInputS0xD(117)(2) <= CNStageIntLLROutputS0xD(111)(1);
  VNStageIntLLRInputS0xD(136)(2) <= CNStageIntLLROutputS0xD(111)(2);
  VNStageIntLLRInputS0xD(198)(2) <= CNStageIntLLROutputS0xD(111)(3);
  VNStageIntLLRInputS0xD(297)(2) <= CNStageIntLLROutputS0xD(111)(4);
  VNStageIntLLRInputS0xD(382)(1) <= CNStageIntLLROutputS0xD(111)(5);
  VNStageIntLLRInputS0xD(30)(2) <= CNStageIntLLROutputS0xD(112)(0);
  VNStageIntLLRInputS0xD(68)(1) <= CNStageIntLLROutputS0xD(112)(1);
  VNStageIntLLRInputS0xD(167)(2) <= CNStageIntLLROutputS0xD(112)(2);
  VNStageIntLLRInputS0xD(252)(1) <= CNStageIntLLROutputS0xD(112)(3);
  VNStageIntLLRInputS0xD(303)(2) <= CNStageIntLLROutputS0xD(112)(4);
  VNStageIntLLRInputS0xD(358)(2) <= CNStageIntLLROutputS0xD(112)(5);
  VNStageIntLLRInputS0xD(29)(2) <= CNStageIntLLROutputS0xD(113)(0);
  VNStageIntLLRInputS0xD(102)(2) <= CNStageIntLLROutputS0xD(113)(1);
  VNStageIntLLRInputS0xD(187)(1) <= CNStageIntLLROutputS0xD(113)(2);
  VNStageIntLLRInputS0xD(238)(2) <= CNStageIntLLROutputS0xD(113)(3);
  VNStageIntLLRInputS0xD(293)(2) <= CNStageIntLLROutputS0xD(113)(4);
  VNStageIntLLRInputS0xD(324)(2) <= CNStageIntLLROutputS0xD(113)(5);
  VNStageIntLLRInputS0xD(28)(2) <= CNStageIntLLROutputS0xD(114)(0);
  VNStageIntLLRInputS0xD(122)(1) <= CNStageIntLLROutputS0xD(114)(1);
  VNStageIntLLRInputS0xD(173)(2) <= CNStageIntLLROutputS0xD(114)(2);
  VNStageIntLLRInputS0xD(228)(2) <= CNStageIntLLROutputS0xD(114)(3);
  VNStageIntLLRInputS0xD(259)(1) <= CNStageIntLLROutputS0xD(114)(4);
  VNStageIntLLRInputS0xD(370)(1) <= CNStageIntLLROutputS0xD(114)(5);
  VNStageIntLLRInputS0xD(27)(2) <= CNStageIntLLROutputS0xD(115)(0);
  VNStageIntLLRInputS0xD(108)(2) <= CNStageIntLLROutputS0xD(115)(1);
  VNStageIntLLRInputS0xD(163)(2) <= CNStageIntLLROutputS0xD(115)(2);
  VNStageIntLLRInputS0xD(194)(2) <= CNStageIntLLROutputS0xD(115)(3);
  VNStageIntLLRInputS0xD(305)(2) <= CNStageIntLLROutputS0xD(115)(4);
  VNStageIntLLRInputS0xD(337)(2) <= CNStageIntLLROutputS0xD(115)(5);
  VNStageIntLLRInputS0xD(26)(2) <= CNStageIntLLROutputS0xD(116)(0);
  VNStageIntLLRInputS0xD(98)(1) <= CNStageIntLLROutputS0xD(116)(1);
  VNStageIntLLRInputS0xD(129)(2) <= CNStageIntLLROutputS0xD(116)(2);
  VNStageIntLLRInputS0xD(240)(2) <= CNStageIntLLROutputS0xD(116)(3);
  VNStageIntLLRInputS0xD(272)(2) <= CNStageIntLLROutputS0xD(116)(4);
  VNStageIntLLRInputS0xD(360)(2) <= CNStageIntLLROutputS0xD(116)(5);
  VNStageIntLLRInputS0xD(25)(2) <= CNStageIntLLROutputS0xD(117)(0);
  VNStageIntLLRInputS0xD(127)(2) <= CNStageIntLLROutputS0xD(117)(1);
  VNStageIntLLRInputS0xD(175)(2) <= CNStageIntLLROutputS0xD(117)(2);
  VNStageIntLLRInputS0xD(207)(2) <= CNStageIntLLROutputS0xD(117)(3);
  VNStageIntLLRInputS0xD(295)(2) <= CNStageIntLLROutputS0xD(117)(4);
  VNStageIntLLRInputS0xD(333)(1) <= CNStageIntLLROutputS0xD(117)(5);
  VNStageIntLLRInputS0xD(24)(2) <= CNStageIntLLROutputS0xD(118)(0);
  VNStageIntLLRInputS0xD(110)(2) <= CNStageIntLLROutputS0xD(118)(1);
  VNStageIntLLRInputS0xD(142)(2) <= CNStageIntLLROutputS0xD(118)(2);
  VNStageIntLLRInputS0xD(230)(1) <= CNStageIntLLROutputS0xD(118)(3);
  VNStageIntLLRInputS0xD(268)(2) <= CNStageIntLLROutputS0xD(118)(4);
  VNStageIntLLRInputS0xD(380)(1) <= CNStageIntLLROutputS0xD(118)(5);
  VNStageIntLLRInputS0xD(23)(2) <= CNStageIntLLROutputS0xD(119)(0);
  VNStageIntLLRInputS0xD(77)(0) <= CNStageIntLLROutputS0xD(119)(1);
  VNStageIntLLRInputS0xD(165)(2) <= CNStageIntLLROutputS0xD(119)(2);
  VNStageIntLLRInputS0xD(203)(2) <= CNStageIntLLROutputS0xD(119)(3);
  VNStageIntLLRInputS0xD(315)(1) <= CNStageIntLLROutputS0xD(119)(4);
  VNStageIntLLRInputS0xD(383)(2) <= CNStageIntLLROutputS0xD(119)(5);
  VNStageIntLLRInputS0xD(22)(2) <= CNStageIntLLROutputS0xD(120)(0);
  VNStageIntLLRInputS0xD(100)(2) <= CNStageIntLLROutputS0xD(120)(1);
  VNStageIntLLRInputS0xD(138)(2) <= CNStageIntLLROutputS0xD(120)(2);
  VNStageIntLLRInputS0xD(250)(1) <= CNStageIntLLROutputS0xD(120)(3);
  VNStageIntLLRInputS0xD(318)(0) <= CNStageIntLLROutputS0xD(120)(4);
  VNStageIntLLRInputS0xD(361)(2) <= CNStageIntLLROutputS0xD(120)(5);
  VNStageIntLLRInputS0xD(21)(2) <= CNStageIntLLROutputS0xD(121)(0);
  VNStageIntLLRInputS0xD(73)(2) <= CNStageIntLLROutputS0xD(121)(1);
  VNStageIntLLRInputS0xD(185)(0) <= CNStageIntLLROutputS0xD(121)(2);
  VNStageIntLLRInputS0xD(253)(1) <= CNStageIntLLROutputS0xD(121)(3);
  VNStageIntLLRInputS0xD(296)(2) <= CNStageIntLLROutputS0xD(121)(4);
  VNStageIntLLRInputS0xD(336)(2) <= CNStageIntLLROutputS0xD(121)(5);
  VNStageIntLLRInputS0xD(19)(2) <= CNStageIntLLROutputS0xD(122)(0);
  VNStageIntLLRInputS0xD(123)(1) <= CNStageIntLLROutputS0xD(122)(1);
  VNStageIntLLRInputS0xD(166)(2) <= CNStageIntLLROutputS0xD(122)(2);
  VNStageIntLLRInputS0xD(206)(1) <= CNStageIntLLROutputS0xD(122)(3);
  VNStageIntLLRInputS0xD(269)(1) <= CNStageIntLLROutputS0xD(122)(4);
  VNStageIntLLRInputS0xD(359)(2) <= CNStageIntLLROutputS0xD(122)(5);
  VNStageIntLLRInputS0xD(18)(2) <= CNStageIntLLROutputS0xD(123)(0);
  VNStageIntLLRInputS0xD(101)(2) <= CNStageIntLLROutputS0xD(123)(1);
  VNStageIntLLRInputS0xD(141)(0) <= CNStageIntLLROutputS0xD(123)(2);
  VNStageIntLLRInputS0xD(204)(2) <= CNStageIntLLROutputS0xD(123)(3);
  VNStageIntLLRInputS0xD(294)(2) <= CNStageIntLLROutputS0xD(123)(4);
  VNStageIntLLRInputS0xD(367)(2) <= CNStageIntLLROutputS0xD(123)(5);
  VNStageIntLLRInputS0xD(17)(2) <= CNStageIntLLROutputS0xD(124)(0);
  VNStageIntLLRInputS0xD(76)(2) <= CNStageIntLLROutputS0xD(124)(1);
  VNStageIntLLRInputS0xD(139)(2) <= CNStageIntLLROutputS0xD(124)(2);
  VNStageIntLLRInputS0xD(229)(2) <= CNStageIntLLROutputS0xD(124)(3);
  VNStageIntLLRInputS0xD(302)(2) <= CNStageIntLLROutputS0xD(124)(4);
  VNStageIntLLRInputS0xD(347)(2) <= CNStageIntLLROutputS0xD(124)(5);
  VNStageIntLLRInputS0xD(16)(1) <= CNStageIntLLROutputS0xD(125)(0);
  VNStageIntLLRInputS0xD(74)(2) <= CNStageIntLLROutputS0xD(125)(1);
  VNStageIntLLRInputS0xD(164)(2) <= CNStageIntLLROutputS0xD(125)(2);
  VNStageIntLLRInputS0xD(237)(2) <= CNStageIntLLROutputS0xD(125)(3);
  VNStageIntLLRInputS0xD(282)(2) <= CNStageIntLLROutputS0xD(125)(4);
  VNStageIntLLRInputS0xD(341)(2) <= CNStageIntLLROutputS0xD(125)(5);
  VNStageIntLLRInputS0xD(15)(2) <= CNStageIntLLROutputS0xD(126)(0);
  VNStageIntLLRInputS0xD(99)(2) <= CNStageIntLLROutputS0xD(126)(1);
  VNStageIntLLRInputS0xD(172)(2) <= CNStageIntLLROutputS0xD(126)(2);
  VNStageIntLLRInputS0xD(217)(2) <= CNStageIntLLROutputS0xD(126)(3);
  VNStageIntLLRInputS0xD(276)(2) <= CNStageIntLLROutputS0xD(126)(4);
  VNStageIntLLRInputS0xD(320)(1) <= CNStageIntLLROutputS0xD(126)(5);
  VNStageIntLLRInputS0xD(14)(2) <= CNStageIntLLROutputS0xD(127)(0);
  VNStageIntLLRInputS0xD(107)(1) <= CNStageIntLLROutputS0xD(127)(1);
  VNStageIntLLRInputS0xD(152)(2) <= CNStageIntLLROutputS0xD(127)(2);
  VNStageIntLLRInputS0xD(211)(2) <= CNStageIntLLROutputS0xD(127)(3);
  VNStageIntLLRInputS0xD(256)(2) <= CNStageIntLLROutputS0xD(127)(4);
  VNStageIntLLRInputS0xD(340)(2) <= CNStageIntLLROutputS0xD(127)(5);
  VNStageIntLLRInputS0xD(13)(1) <= CNStageIntLLROutputS0xD(128)(0);
  VNStageIntLLRInputS0xD(87)(2) <= CNStageIntLLROutputS0xD(128)(1);
  VNStageIntLLRInputS0xD(146)(2) <= CNStageIntLLROutputS0xD(128)(2);
  VNStageIntLLRInputS0xD(192)(2) <= CNStageIntLLROutputS0xD(128)(3);
  VNStageIntLLRInputS0xD(275)(2) <= CNStageIntLLROutputS0xD(128)(4);
  VNStageIntLLRInputS0xD(345)(2) <= CNStageIntLLROutputS0xD(128)(5);
  VNStageIntLLRInputS0xD(12)(2) <= CNStageIntLLROutputS0xD(129)(0);
  VNStageIntLLRInputS0xD(81)(2) <= CNStageIntLLROutputS0xD(129)(1);
  VNStageIntLLRInputS0xD(128)(2) <= CNStageIntLLROutputS0xD(129)(2);
  VNStageIntLLRInputS0xD(210)(2) <= CNStageIntLLROutputS0xD(129)(3);
  VNStageIntLLRInputS0xD(280)(2) <= CNStageIntLLROutputS0xD(129)(4);
  VNStageIntLLRInputS0xD(364)(2) <= CNStageIntLLROutputS0xD(129)(5);
  VNStageIntLLRInputS0xD(11)(2) <= CNStageIntLLROutputS0xD(130)(0);
  VNStageIntLLRInputS0xD(64)(2) <= CNStageIntLLROutputS0xD(130)(1);
  VNStageIntLLRInputS0xD(145)(2) <= CNStageIntLLROutputS0xD(130)(2);
  VNStageIntLLRInputS0xD(215)(2) <= CNStageIntLLROutputS0xD(130)(3);
  VNStageIntLLRInputS0xD(299)(1) <= CNStageIntLLROutputS0xD(130)(4);
  VNStageIntLLRInputS0xD(355)(2) <= CNStageIntLLROutputS0xD(130)(5);
  VNStageIntLLRInputS0xD(10)(2) <= CNStageIntLLROutputS0xD(131)(0);
  VNStageIntLLRInputS0xD(80)(2) <= CNStageIntLLROutputS0xD(131)(1);
  VNStageIntLLRInputS0xD(150)(2) <= CNStageIntLLROutputS0xD(131)(2);
  VNStageIntLLRInputS0xD(234)(2) <= CNStageIntLLROutputS0xD(131)(3);
  VNStageIntLLRInputS0xD(290)(2) <= CNStageIntLLROutputS0xD(131)(4);
  VNStageIntLLRInputS0xD(329)(2) <= CNStageIntLLROutputS0xD(131)(5);
  VNStageIntLLRInputS0xD(9)(2) <= CNStageIntLLROutputS0xD(132)(0);
  VNStageIntLLRInputS0xD(85)(1) <= CNStageIntLLROutputS0xD(132)(1);
  VNStageIntLLRInputS0xD(169)(2) <= CNStageIntLLROutputS0xD(132)(2);
  VNStageIntLLRInputS0xD(225)(2) <= CNStageIntLLROutputS0xD(132)(3);
  VNStageIntLLRInputS0xD(264)(2) <= CNStageIntLLROutputS0xD(132)(4);
  VNStageIntLLRInputS0xD(330)(2) <= CNStageIntLLROutputS0xD(132)(5);
  VNStageIntLLRInputS0xD(8)(1) <= CNStageIntLLROutputS0xD(133)(0);
  VNStageIntLLRInputS0xD(104)(2) <= CNStageIntLLROutputS0xD(133)(1);
  VNStageIntLLRInputS0xD(160)(2) <= CNStageIntLLROutputS0xD(133)(2);
  VNStageIntLLRInputS0xD(199)(2) <= CNStageIntLLROutputS0xD(133)(3);
  VNStageIntLLRInputS0xD(265)(1) <= CNStageIntLLROutputS0xD(133)(4);
  VNStageIntLLRInputS0xD(354)(2) <= CNStageIntLLROutputS0xD(133)(5);
  VNStageIntLLRInputS0xD(7)(2) <= CNStageIntLLROutputS0xD(134)(0);
  VNStageIntLLRInputS0xD(95)(2) <= CNStageIntLLROutputS0xD(134)(1);
  VNStageIntLLRInputS0xD(134)(2) <= CNStageIntLLROutputS0xD(134)(2);
  VNStageIntLLRInputS0xD(200)(2) <= CNStageIntLLROutputS0xD(134)(3);
  VNStageIntLLRInputS0xD(289)(2) <= CNStageIntLLROutputS0xD(134)(4);
  VNStageIntLLRInputS0xD(375)(2) <= CNStageIntLLROutputS0xD(134)(5);
  VNStageIntLLRInputS0xD(6)(2) <= CNStageIntLLROutputS0xD(135)(0);
  VNStageIntLLRInputS0xD(69)(2) <= CNStageIntLLROutputS0xD(135)(1);
  VNStageIntLLRInputS0xD(135)(2) <= CNStageIntLLROutputS0xD(135)(2);
  VNStageIntLLRInputS0xD(224)(2) <= CNStageIntLLROutputS0xD(135)(3);
  VNStageIntLLRInputS0xD(310)(2) <= CNStageIntLLROutputS0xD(135)(4);
  VNStageIntLLRInputS0xD(371)(1) <= CNStageIntLLROutputS0xD(135)(5);
  VNStageIntLLRInputS0xD(5)(2) <= CNStageIntLLROutputS0xD(136)(0);
  VNStageIntLLRInputS0xD(70)(2) <= CNStageIntLLROutputS0xD(136)(1);
  VNStageIntLLRInputS0xD(159)(2) <= CNStageIntLLROutputS0xD(136)(2);
  VNStageIntLLRInputS0xD(245)(2) <= CNStageIntLLROutputS0xD(136)(3);
  VNStageIntLLRInputS0xD(306)(2) <= CNStageIntLLROutputS0xD(136)(4);
  VNStageIntLLRInputS0xD(323)(1) <= CNStageIntLLROutputS0xD(136)(5);
  VNStageIntLLRInputS0xD(3)(1) <= CNStageIntLLROutputS0xD(137)(0);
  VNStageIntLLRInputS0xD(115)(2) <= CNStageIntLLROutputS0xD(137)(1);
  VNStageIntLLRInputS0xD(176)(2) <= CNStageIntLLROutputS0xD(137)(2);
  VNStageIntLLRInputS0xD(193)(2) <= CNStageIntLLROutputS0xD(137)(3);
  VNStageIntLLRInputS0xD(284)(2) <= CNStageIntLLROutputS0xD(137)(4);
  VNStageIntLLRInputS0xD(325)(2) <= CNStageIntLLROutputS0xD(137)(5);
  VNStageIntLLRInputS0xD(2)(2) <= CNStageIntLLROutputS0xD(138)(0);
  VNStageIntLLRInputS0xD(111)(2) <= CNStageIntLLROutputS0xD(138)(1);
  VNStageIntLLRInputS0xD(191)(2) <= CNStageIntLLROutputS0xD(138)(2);
  VNStageIntLLRInputS0xD(219)(2) <= CNStageIntLLROutputS0xD(138)(3);
  VNStageIntLLRInputS0xD(260)(2) <= CNStageIntLLROutputS0xD(138)(4);
  VNStageIntLLRInputS0xD(357)(2) <= CNStageIntLLROutputS0xD(138)(5);
  VNStageIntLLRInputS0xD(1)(1) <= CNStageIntLLROutputS0xD(139)(0);
  VNStageIntLLRInputS0xD(126)(1) <= CNStageIntLLROutputS0xD(139)(1);
  VNStageIntLLRInputS0xD(154)(1) <= CNStageIntLLROutputS0xD(139)(2);
  VNStageIntLLRInputS0xD(195)(1) <= CNStageIntLLROutputS0xD(139)(3);
  VNStageIntLLRInputS0xD(292)(2) <= CNStageIntLLROutputS0xD(139)(4);
  VNStageIntLLRInputS0xD(373)(1) <= CNStageIntLLROutputS0xD(139)(5);
  VNStageIntLLRInputS0xD(63)(2) <= CNStageIntLLROutputS0xD(140)(0);
  VNStageIntLLRInputS0xD(89)(2) <= CNStageIntLLROutputS0xD(140)(1);
  VNStageIntLLRInputS0xD(130)(2) <= CNStageIntLLROutputS0xD(140)(2);
  VNStageIntLLRInputS0xD(227)(2) <= CNStageIntLLROutputS0xD(140)(3);
  VNStageIntLLRInputS0xD(308)(0) <= CNStageIntLLROutputS0xD(140)(4);
  VNStageIntLLRInputS0xD(343)(2) <= CNStageIntLLROutputS0xD(140)(5);
  VNStageIntLLRInputS0xD(62)(1) <= CNStageIntLLROutputS0xD(141)(0);
  VNStageIntLLRInputS0xD(65)(2) <= CNStageIntLLROutputS0xD(141)(1);
  VNStageIntLLRInputS0xD(162)(2) <= CNStageIntLLROutputS0xD(141)(2);
  VNStageIntLLRInputS0xD(243)(2) <= CNStageIntLLROutputS0xD(141)(3);
  VNStageIntLLRInputS0xD(278)(2) <= CNStageIntLLROutputS0xD(141)(4);
  VNStageIntLLRInputS0xD(352)(2) <= CNStageIntLLROutputS0xD(141)(5);
  VNStageIntLLRInputS0xD(61)(1) <= CNStageIntLLROutputS0xD(142)(0);
  VNStageIntLLRInputS0xD(97)(2) <= CNStageIntLLROutputS0xD(142)(1);
  VNStageIntLLRInputS0xD(178)(2) <= CNStageIntLLROutputS0xD(142)(2);
  VNStageIntLLRInputS0xD(213)(2) <= CNStageIntLLROutputS0xD(142)(3);
  VNStageIntLLRInputS0xD(287)(2) <= CNStageIntLLROutputS0xD(142)(4);
  VNStageIntLLRInputS0xD(365)(2) <= CNStageIntLLROutputS0xD(142)(5);
  VNStageIntLLRInputS0xD(60)(1) <= CNStageIntLLROutputS0xD(143)(0);
  VNStageIntLLRInputS0xD(113)(2) <= CNStageIntLLROutputS0xD(143)(1);
  VNStageIntLLRInputS0xD(148)(2) <= CNStageIntLLROutputS0xD(143)(2);
  VNStageIntLLRInputS0xD(222)(1) <= CNStageIntLLROutputS0xD(143)(3);
  VNStageIntLLRInputS0xD(300)(2) <= CNStageIntLLROutputS0xD(143)(4);
  VNStageIntLLRInputS0xD(344)(2) <= CNStageIntLLROutputS0xD(143)(5);
  VNStageIntLLRInputS0xD(59)(0) <= CNStageIntLLROutputS0xD(144)(0);
  VNStageIntLLRInputS0xD(83)(2) <= CNStageIntLLROutputS0xD(144)(1);
  VNStageIntLLRInputS0xD(157)(2) <= CNStageIntLLROutputS0xD(144)(2);
  VNStageIntLLRInputS0xD(235)(1) <= CNStageIntLLROutputS0xD(144)(3);
  VNStageIntLLRInputS0xD(279)(2) <= CNStageIntLLROutputS0xD(144)(4);
  VNStageIntLLRInputS0xD(372)(1) <= CNStageIntLLROutputS0xD(144)(5);
  VNStageIntLLRInputS0xD(58)(1) <= CNStageIntLLROutputS0xD(145)(0);
  VNStageIntLLRInputS0xD(92)(2) <= CNStageIntLLROutputS0xD(145)(1);
  VNStageIntLLRInputS0xD(170)(2) <= CNStageIntLLROutputS0xD(145)(2);
  VNStageIntLLRInputS0xD(214)(2) <= CNStageIntLLROutputS0xD(145)(3);
  VNStageIntLLRInputS0xD(307)(2) <= CNStageIntLLROutputS0xD(145)(4);
  VNStageIntLLRInputS0xD(374)(2) <= CNStageIntLLROutputS0xD(145)(5);
  VNStageIntLLRInputS0xD(57)(1) <= CNStageIntLLROutputS0xD(146)(0);
  VNStageIntLLRInputS0xD(105)(1) <= CNStageIntLLROutputS0xD(146)(1);
  VNStageIntLLRInputS0xD(149)(2) <= CNStageIntLLROutputS0xD(146)(2);
  VNStageIntLLRInputS0xD(242)(2) <= CNStageIntLLROutputS0xD(146)(3);
  VNStageIntLLRInputS0xD(309)(2) <= CNStageIntLLROutputS0xD(146)(4);
  VNStageIntLLRInputS0xD(356)(2) <= CNStageIntLLROutputS0xD(146)(5);
  VNStageIntLLRInputS0xD(56)(2) <= CNStageIntLLROutputS0xD(147)(0);
  VNStageIntLLRInputS0xD(84)(2) <= CNStageIntLLROutputS0xD(147)(1);
  VNStageIntLLRInputS0xD(177)(2) <= CNStageIntLLROutputS0xD(147)(2);
  VNStageIntLLRInputS0xD(244)(0) <= CNStageIntLLROutputS0xD(147)(3);
  VNStageIntLLRInputS0xD(291)(2) <= CNStageIntLLROutputS0xD(147)(4);
  VNStageIntLLRInputS0xD(363)(1) <= CNStageIntLLROutputS0xD(147)(5);
  VNStageIntLLRInputS0xD(55)(2) <= CNStageIntLLROutputS0xD(148)(0);
  VNStageIntLLRInputS0xD(112)(2) <= CNStageIntLLROutputS0xD(148)(1);
  VNStageIntLLRInputS0xD(179)(2) <= CNStageIntLLROutputS0xD(148)(2);
  VNStageIntLLRInputS0xD(226)(1) <= CNStageIntLLROutputS0xD(148)(3);
  VNStageIntLLRInputS0xD(298)(2) <= CNStageIntLLROutputS0xD(148)(4);
  VNStageIntLLRInputS0xD(327)(2) <= CNStageIntLLROutputS0xD(148)(5);
  VNStageIntLLRInputS0xD(54)(2) <= CNStageIntLLROutputS0xD(149)(0);
  VNStageIntLLRInputS0xD(114)(2) <= CNStageIntLLROutputS0xD(149)(1);
  VNStageIntLLRInputS0xD(161)(2) <= CNStageIntLLROutputS0xD(149)(2);
  VNStageIntLLRInputS0xD(233)(2) <= CNStageIntLLROutputS0xD(149)(3);
  VNStageIntLLRInputS0xD(262)(2) <= CNStageIntLLROutputS0xD(149)(4);
  VNStageIntLLRInputS0xD(378)(1) <= CNStageIntLLROutputS0xD(149)(5);
  VNStageIntLLRInputS0xD(53)(1) <= CNStageIntLLROutputS0xD(150)(0);
  VNStageIntLLRInputS0xD(96)(2) <= CNStageIntLLROutputS0xD(150)(1);
  VNStageIntLLRInputS0xD(168)(1) <= CNStageIntLLROutputS0xD(150)(2);
  VNStageIntLLRInputS0xD(197)(2) <= CNStageIntLLROutputS0xD(150)(3);
  VNStageIntLLRInputS0xD(313)(0) <= CNStageIntLLROutputS0xD(150)(4);
  VNStageIntLLRInputS0xD(321)(2) <= CNStageIntLLROutputS0xD(150)(5);
  VNStageIntLLRInputS0xD(52)(1) <= CNStageIntLLROutputS0xD(151)(0);
  VNStageIntLLRInputS0xD(103)(2) <= CNStageIntLLROutputS0xD(151)(1);
  VNStageIntLLRInputS0xD(132)(1) <= CNStageIntLLROutputS0xD(151)(2);
  VNStageIntLLRInputS0xD(248)(2) <= CNStageIntLLROutputS0xD(151)(3);
  VNStageIntLLRInputS0xD(319)(2) <= CNStageIntLLROutputS0xD(151)(4);
  VNStageIntLLRInputS0xD(379)(1) <= CNStageIntLLROutputS0xD(151)(5);
  VNStageIntLLRInputS0xD(50)(2) <= CNStageIntLLROutputS0xD(152)(0);
  VNStageIntLLRInputS0xD(118)(2) <= CNStageIntLLROutputS0xD(152)(1);
  VNStageIntLLRInputS0xD(189)(1) <= CNStageIntLLROutputS0xD(152)(2);
  VNStageIntLLRInputS0xD(249)(0) <= CNStageIntLLROutputS0xD(152)(3);
  VNStageIntLLRInputS0xD(261)(2) <= CNStageIntLLROutputS0xD(152)(4);
  VNStageIntLLRInputS0xD(348)(2) <= CNStageIntLLROutputS0xD(152)(5);
  VNStageIntLLRInputS0xD(49)(2) <= CNStageIntLLROutputS0xD(153)(0);
  VNStageIntLLRInputS0xD(124)(1) <= CNStageIntLLROutputS0xD(153)(1);
  VNStageIntLLRInputS0xD(184)(2) <= CNStageIntLLROutputS0xD(153)(2);
  VNStageIntLLRInputS0xD(196)(2) <= CNStageIntLLROutputS0xD(153)(3);
  VNStageIntLLRInputS0xD(283)(2) <= CNStageIntLLROutputS0xD(153)(4);
  VNStageIntLLRInputS0xD(366)(2) <= CNStageIntLLROutputS0xD(153)(5);
  VNStageIntLLRInputS0xD(48)(1) <= CNStageIntLLROutputS0xD(154)(0);
  VNStageIntLLRInputS0xD(119)(2) <= CNStageIntLLROutputS0xD(154)(1);
  VNStageIntLLRInputS0xD(131)(1) <= CNStageIntLLROutputS0xD(154)(2);
  VNStageIntLLRInputS0xD(218)(2) <= CNStageIntLLROutputS0xD(154)(3);
  VNStageIntLLRInputS0xD(301)(2) <= CNStageIntLLROutputS0xD(154)(4);
  VNStageIntLLRInputS0xD(351)(1) <= CNStageIntLLROutputS0xD(154)(5);
  VNStageIntLLRInputS0xD(47)(1) <= CNStageIntLLROutputS0xD(155)(0);
  VNStageIntLLRInputS0xD(66)(2) <= CNStageIntLLROutputS0xD(155)(1);
  VNStageIntLLRInputS0xD(153)(2) <= CNStageIntLLROutputS0xD(155)(2);
  VNStageIntLLRInputS0xD(236)(2) <= CNStageIntLLROutputS0xD(155)(3);
  VNStageIntLLRInputS0xD(286)(2) <= CNStageIntLLROutputS0xD(155)(4);
  VNStageIntLLRInputS0xD(338)(2) <= CNStageIntLLROutputS0xD(155)(5);
  VNStageIntLLRInputS0xD(46)(2) <= CNStageIntLLROutputS0xD(156)(0);
  VNStageIntLLRInputS0xD(88)(2) <= CNStageIntLLROutputS0xD(156)(1);
  VNStageIntLLRInputS0xD(171)(1) <= CNStageIntLLROutputS0xD(156)(2);
  VNStageIntLLRInputS0xD(221)(2) <= CNStageIntLLROutputS0xD(156)(3);
  VNStageIntLLRInputS0xD(273)(2) <= CNStageIntLLROutputS0xD(156)(4);
  VNStageIntLLRInputS0xD(369)(1) <= CNStageIntLLROutputS0xD(156)(5);
  VNStageIntLLRInputS0xD(45)(2) <= CNStageIntLLROutputS0xD(157)(0);
  VNStageIntLLRInputS0xD(106)(1) <= CNStageIntLLROutputS0xD(157)(1);
  VNStageIntLLRInputS0xD(156)(2) <= CNStageIntLLROutputS0xD(157)(2);
  VNStageIntLLRInputS0xD(208)(2) <= CNStageIntLLROutputS0xD(157)(3);
  VNStageIntLLRInputS0xD(304)(2) <= CNStageIntLLROutputS0xD(157)(4);
  VNStageIntLLRInputS0xD(381)(1) <= CNStageIntLLROutputS0xD(157)(5);
  VNStageIntLLRInputS0xD(44)(2) <= CNStageIntLLROutputS0xD(158)(0);
  VNStageIntLLRInputS0xD(91)(2) <= CNStageIntLLROutputS0xD(158)(1);
  VNStageIntLLRInputS0xD(143)(2) <= CNStageIntLLROutputS0xD(158)(2);
  VNStageIntLLRInputS0xD(239)(2) <= CNStageIntLLROutputS0xD(158)(3);
  VNStageIntLLRInputS0xD(316)(1) <= CNStageIntLLROutputS0xD(158)(4);
  VNStageIntLLRInputS0xD(332)(2) <= CNStageIntLLROutputS0xD(158)(5);
  VNStageIntLLRInputS0xD(43)(1) <= CNStageIntLLROutputS0xD(159)(0);
  VNStageIntLLRInputS0xD(78)(2) <= CNStageIntLLROutputS0xD(159)(1);
  VNStageIntLLRInputS0xD(174)(2) <= CNStageIntLLROutputS0xD(159)(2);
  VNStageIntLLRInputS0xD(251)(1) <= CNStageIntLLROutputS0xD(159)(3);
  VNStageIntLLRInputS0xD(267)(2) <= CNStageIntLLROutputS0xD(159)(4);
  VNStageIntLLRInputS0xD(376)(2) <= CNStageIntLLROutputS0xD(159)(5);
  VNStageIntLLRInputS0xD(42)(2) <= CNStageIntLLROutputS0xD(160)(0);
  VNStageIntLLRInputS0xD(109)(2) <= CNStageIntLLROutputS0xD(160)(1);
  VNStageIntLLRInputS0xD(186)(1) <= CNStageIntLLROutputS0xD(160)(2);
  VNStageIntLLRInputS0xD(202)(2) <= CNStageIntLLROutputS0xD(160)(3);
  VNStageIntLLRInputS0xD(311)(2) <= CNStageIntLLROutputS0xD(160)(4);
  VNStageIntLLRInputS0xD(353)(2) <= CNStageIntLLROutputS0xD(160)(5);
  VNStageIntLLRInputS0xD(41)(2) <= CNStageIntLLROutputS0xD(161)(0);
  VNStageIntLLRInputS0xD(121)(1) <= CNStageIntLLROutputS0xD(161)(1);
  VNStageIntLLRInputS0xD(137)(2) <= CNStageIntLLROutputS0xD(161)(2);
  VNStageIntLLRInputS0xD(246)(2) <= CNStageIntLLROutputS0xD(161)(3);
  VNStageIntLLRInputS0xD(288)(2) <= CNStageIntLLROutputS0xD(161)(4);
  VNStageIntLLRInputS0xD(342)(2) <= CNStageIntLLROutputS0xD(161)(5);
  VNStageIntLLRInputS0xD(40)(2) <= CNStageIntLLROutputS0xD(162)(0);
  VNStageIntLLRInputS0xD(72)(2) <= CNStageIntLLROutputS0xD(162)(1);
  VNStageIntLLRInputS0xD(181)(2) <= CNStageIntLLROutputS0xD(162)(2);
  VNStageIntLLRInputS0xD(223)(2) <= CNStageIntLLROutputS0xD(162)(3);
  VNStageIntLLRInputS0xD(277)(2) <= CNStageIntLLROutputS0xD(162)(4);
  VNStageIntLLRInputS0xD(346)(2) <= CNStageIntLLROutputS0xD(162)(5);
  VNStageIntLLRInputS0xD(39)(2) <= CNStageIntLLROutputS0xD(163)(0);
  VNStageIntLLRInputS0xD(116)(1) <= CNStageIntLLROutputS0xD(163)(1);
  VNStageIntLLRInputS0xD(158)(2) <= CNStageIntLLROutputS0xD(163)(2);
  VNStageIntLLRInputS0xD(212)(2) <= CNStageIntLLROutputS0xD(163)(3);
  VNStageIntLLRInputS0xD(281)(2) <= CNStageIntLLROutputS0xD(163)(4);
  VNStageIntLLRInputS0xD(339)(2) <= CNStageIntLLROutputS0xD(163)(5);
  VNStageIntLLRInputS0xD(38)(2) <= CNStageIntLLROutputS0xD(164)(0);
  VNStageIntLLRInputS0xD(93)(2) <= CNStageIntLLROutputS0xD(164)(1);
  VNStageIntLLRInputS0xD(147)(2) <= CNStageIntLLROutputS0xD(164)(2);
  VNStageIntLLRInputS0xD(216)(2) <= CNStageIntLLROutputS0xD(164)(3);
  VNStageIntLLRInputS0xD(274)(1) <= CNStageIntLLROutputS0xD(164)(4);
  VNStageIntLLRInputS0xD(350)(2) <= CNStageIntLLROutputS0xD(164)(5);
  VNStageIntLLRInputS0xD(37)(2) <= CNStageIntLLROutputS0xD(165)(0);
  VNStageIntLLRInputS0xD(82)(2) <= CNStageIntLLROutputS0xD(165)(1);
  VNStageIntLLRInputS0xD(151)(2) <= CNStageIntLLROutputS0xD(165)(2);
  VNStageIntLLRInputS0xD(209)(2) <= CNStageIntLLROutputS0xD(165)(3);
  VNStageIntLLRInputS0xD(285)(2) <= CNStageIntLLROutputS0xD(165)(4);
  VNStageIntLLRInputS0xD(322)(2) <= CNStageIntLLROutputS0xD(165)(5);
  VNStageIntLLRInputS0xD(36)(2) <= CNStageIntLLROutputS0xD(166)(0);
  VNStageIntLLRInputS0xD(86)(1) <= CNStageIntLLROutputS0xD(166)(1);
  VNStageIntLLRInputS0xD(144)(2) <= CNStageIntLLROutputS0xD(166)(2);
  VNStageIntLLRInputS0xD(220)(2) <= CNStageIntLLROutputS0xD(166)(3);
  VNStageIntLLRInputS0xD(257)(2) <= CNStageIntLLROutputS0xD(166)(4);
  VNStageIntLLRInputS0xD(377)(1) <= CNStageIntLLROutputS0xD(166)(5);
  VNStageIntLLRInputS0xD(35)(2) <= CNStageIntLLROutputS0xD(167)(0);
  VNStageIntLLRInputS0xD(79)(2) <= CNStageIntLLROutputS0xD(167)(1);
  VNStageIntLLRInputS0xD(155)(2) <= CNStageIntLLROutputS0xD(167)(2);
  VNStageIntLLRInputS0xD(255)(2) <= CNStageIntLLROutputS0xD(167)(3);
  VNStageIntLLRInputS0xD(312)(2) <= CNStageIntLLROutputS0xD(167)(4);
  VNStageIntLLRInputS0xD(331)(2) <= CNStageIntLLROutputS0xD(167)(5);
  VNStageIntLLRInputS0xD(34)(2) <= CNStageIntLLROutputS0xD(168)(0);
  VNStageIntLLRInputS0xD(90)(2) <= CNStageIntLLROutputS0xD(168)(1);
  VNStageIntLLRInputS0xD(190)(0) <= CNStageIntLLROutputS0xD(168)(2);
  VNStageIntLLRInputS0xD(247)(2) <= CNStageIntLLROutputS0xD(168)(3);
  VNStageIntLLRInputS0xD(266)(1) <= CNStageIntLLROutputS0xD(168)(4);
  VNStageIntLLRInputS0xD(328)(2) <= CNStageIntLLROutputS0xD(168)(5);
  VNStageIntLLRInputS0xD(33)(2) <= CNStageIntLLROutputS0xD(169)(0);
  VNStageIntLLRInputS0xD(125)(1) <= CNStageIntLLROutputS0xD(169)(1);
  VNStageIntLLRInputS0xD(182)(2) <= CNStageIntLLROutputS0xD(169)(2);
  VNStageIntLLRInputS0xD(201)(2) <= CNStageIntLLROutputS0xD(169)(3);
  VNStageIntLLRInputS0xD(263)(2) <= CNStageIntLLROutputS0xD(169)(4);
  VNStageIntLLRInputS0xD(362)(2) <= CNStageIntLLROutputS0xD(169)(5);
  VNStageIntLLRInputS0xD(0)(2) <= CNStageIntLLROutputS0xD(170)(0);
  VNStageIntLLRInputS0xD(75)(2) <= CNStageIntLLROutputS0xD(170)(1);
  VNStageIntLLRInputS0xD(140)(2) <= CNStageIntLLROutputS0xD(170)(2);
  VNStageIntLLRInputS0xD(205)(0) <= CNStageIntLLROutputS0xD(170)(3);
  VNStageIntLLRInputS0xD(270)(2) <= CNStageIntLLROutputS0xD(170)(4);
  VNStageIntLLRInputS0xD(335)(2) <= CNStageIntLLROutputS0xD(170)(5);
  VNStageIntLLRInputS0xD(62)(2) <= CNStageIntLLROutputS0xD(171)(0);
  VNStageIntLLRInputS0xD(109)(3) <= CNStageIntLLROutputS0xD(171)(1);
  VNStageIntLLRInputS0xD(161)(3) <= CNStageIntLLROutputS0xD(171)(2);
  VNStageIntLLRInputS0xD(194)(3) <= CNStageIntLLROutputS0xD(171)(3);
  VNStageIntLLRInputS0xD(271)(2) <= CNStageIntLLROutputS0xD(171)(4);
  VNStageIntLLRInputS0xD(350)(3) <= CNStageIntLLROutputS0xD(171)(5);
  VNStageIntLLRInputS0xD(61)(2) <= CNStageIntLLROutputS0xD(172)(0);
  VNStageIntLLRInputS0xD(96)(3) <= CNStageIntLLROutputS0xD(172)(1);
  VNStageIntLLRInputS0xD(129)(3) <= CNStageIntLLROutputS0xD(172)(2);
  VNStageIntLLRInputS0xD(206)(2) <= CNStageIntLLROutputS0xD(172)(3);
  VNStageIntLLRInputS0xD(285)(3) <= CNStageIntLLROutputS0xD(172)(4);
  VNStageIntLLRInputS0xD(331)(3) <= CNStageIntLLROutputS0xD(172)(5);
  VNStageIntLLRInputS0xD(60)(2) <= CNStageIntLLROutputS0xD(173)(0);
  VNStageIntLLRInputS0xD(127)(3) <= CNStageIntLLROutputS0xD(173)(1);
  VNStageIntLLRInputS0xD(141)(1) <= CNStageIntLLROutputS0xD(173)(2);
  VNStageIntLLRInputS0xD(220)(3) <= CNStageIntLLROutputS0xD(173)(3);
  VNStageIntLLRInputS0xD(266)(2) <= CNStageIntLLROutputS0xD(173)(4);
  VNStageIntLLRInputS0xD(371)(2) <= CNStageIntLLROutputS0xD(173)(5);
  VNStageIntLLRInputS0xD(59)(1) <= CNStageIntLLROutputS0xD(174)(0);
  VNStageIntLLRInputS0xD(76)(3) <= CNStageIntLLROutputS0xD(174)(1);
  VNStageIntLLRInputS0xD(155)(3) <= CNStageIntLLROutputS0xD(174)(2);
  VNStageIntLLRInputS0xD(201)(3) <= CNStageIntLLROutputS0xD(174)(3);
  VNStageIntLLRInputS0xD(306)(3) <= CNStageIntLLROutputS0xD(174)(4);
  VNStageIntLLRInputS0xD(360)(3) <= CNStageIntLLROutputS0xD(174)(5);
  VNStageIntLLRInputS0xD(58)(2) <= CNStageIntLLROutputS0xD(175)(0);
  VNStageIntLLRInputS0xD(90)(3) <= CNStageIntLLROutputS0xD(175)(1);
  VNStageIntLLRInputS0xD(136)(3) <= CNStageIntLLROutputS0xD(175)(2);
  VNStageIntLLRInputS0xD(241)(2) <= CNStageIntLLROutputS0xD(175)(3);
  VNStageIntLLRInputS0xD(295)(3) <= CNStageIntLLROutputS0xD(175)(4);
  VNStageIntLLRInputS0xD(364)(3) <= CNStageIntLLROutputS0xD(175)(5);
  VNStageIntLLRInputS0xD(57)(2) <= CNStageIntLLROutputS0xD(176)(0);
  VNStageIntLLRInputS0xD(71)(2) <= CNStageIntLLROutputS0xD(176)(1);
  VNStageIntLLRInputS0xD(176)(3) <= CNStageIntLLROutputS0xD(176)(2);
  VNStageIntLLRInputS0xD(230)(2) <= CNStageIntLLROutputS0xD(176)(3);
  VNStageIntLLRInputS0xD(299)(2) <= CNStageIntLLROutputS0xD(176)(4);
  VNStageIntLLRInputS0xD(357)(3) <= CNStageIntLLROutputS0xD(176)(5);
  VNStageIntLLRInputS0xD(56)(3) <= CNStageIntLLROutputS0xD(177)(0);
  VNStageIntLLRInputS0xD(111)(3) <= CNStageIntLLROutputS0xD(177)(1);
  VNStageIntLLRInputS0xD(165)(3) <= CNStageIntLLROutputS0xD(177)(2);
  VNStageIntLLRInputS0xD(234)(3) <= CNStageIntLLROutputS0xD(177)(3);
  VNStageIntLLRInputS0xD(292)(3) <= CNStageIntLLROutputS0xD(177)(4);
  VNStageIntLLRInputS0xD(368)(1) <= CNStageIntLLROutputS0xD(177)(5);
  VNStageIntLLRInputS0xD(55)(3) <= CNStageIntLLROutputS0xD(178)(0);
  VNStageIntLLRInputS0xD(100)(3) <= CNStageIntLLROutputS0xD(178)(1);
  VNStageIntLLRInputS0xD(169)(3) <= CNStageIntLLROutputS0xD(178)(2);
  VNStageIntLLRInputS0xD(227)(3) <= CNStageIntLLROutputS0xD(178)(3);
  VNStageIntLLRInputS0xD(303)(3) <= CNStageIntLLROutputS0xD(178)(4);
  VNStageIntLLRInputS0xD(340)(3) <= CNStageIntLLROutputS0xD(178)(5);
  VNStageIntLLRInputS0xD(54)(3) <= CNStageIntLLROutputS0xD(179)(0);
  VNStageIntLLRInputS0xD(104)(3) <= CNStageIntLLROutputS0xD(179)(1);
  VNStageIntLLRInputS0xD(162)(3) <= CNStageIntLLROutputS0xD(179)(2);
  VNStageIntLLRInputS0xD(238)(3) <= CNStageIntLLROutputS0xD(179)(3);
  VNStageIntLLRInputS0xD(275)(3) <= CNStageIntLLROutputS0xD(179)(4);
  VNStageIntLLRInputS0xD(332)(3) <= CNStageIntLLROutputS0xD(179)(5);
  VNStageIntLLRInputS0xD(53)(2) <= CNStageIntLLROutputS0xD(180)(0);
  VNStageIntLLRInputS0xD(97)(3) <= CNStageIntLLROutputS0xD(180)(1);
  VNStageIntLLRInputS0xD(173)(3) <= CNStageIntLLROutputS0xD(180)(2);
  VNStageIntLLRInputS0xD(210)(3) <= CNStageIntLLROutputS0xD(180)(3);
  VNStageIntLLRInputS0xD(267)(3) <= CNStageIntLLROutputS0xD(180)(4);
  VNStageIntLLRInputS0xD(349)(2) <= CNStageIntLLROutputS0xD(180)(5);
  VNStageIntLLRInputS0xD(52)(2) <= CNStageIntLLROutputS0xD(181)(0);
  VNStageIntLLRInputS0xD(108)(3) <= CNStageIntLLROutputS0xD(181)(1);
  VNStageIntLLRInputS0xD(145)(3) <= CNStageIntLLROutputS0xD(181)(2);
  VNStageIntLLRInputS0xD(202)(3) <= CNStageIntLLROutputS0xD(181)(3);
  VNStageIntLLRInputS0xD(284)(3) <= CNStageIntLLROutputS0xD(181)(4);
  VNStageIntLLRInputS0xD(346)(3) <= CNStageIntLLROutputS0xD(181)(5);
  VNStageIntLLRInputS0xD(51)(2) <= CNStageIntLLROutputS0xD(182)(0);
  VNStageIntLLRInputS0xD(80)(3) <= CNStageIntLLROutputS0xD(182)(1);
  VNStageIntLLRInputS0xD(137)(3) <= CNStageIntLLROutputS0xD(182)(2);
  VNStageIntLLRInputS0xD(219)(3) <= CNStageIntLLROutputS0xD(182)(3);
  VNStageIntLLRInputS0xD(281)(3) <= CNStageIntLLROutputS0xD(182)(4);
  VNStageIntLLRInputS0xD(380)(2) <= CNStageIntLLROutputS0xD(182)(5);
  VNStageIntLLRInputS0xD(50)(3) <= CNStageIntLLROutputS0xD(183)(0);
  VNStageIntLLRInputS0xD(72)(3) <= CNStageIntLLROutputS0xD(183)(1);
  VNStageIntLLRInputS0xD(154)(2) <= CNStageIntLLROutputS0xD(183)(2);
  VNStageIntLLRInputS0xD(216)(3) <= CNStageIntLLROutputS0xD(183)(3);
  VNStageIntLLRInputS0xD(315)(2) <= CNStageIntLLROutputS0xD(183)(4);
  VNStageIntLLRInputS0xD(337)(3) <= CNStageIntLLROutputS0xD(183)(5);
  VNStageIntLLRInputS0xD(49)(3) <= CNStageIntLLROutputS0xD(184)(0);
  VNStageIntLLRInputS0xD(89)(3) <= CNStageIntLLROutputS0xD(184)(1);
  VNStageIntLLRInputS0xD(151)(3) <= CNStageIntLLROutputS0xD(184)(2);
  VNStageIntLLRInputS0xD(250)(2) <= CNStageIntLLROutputS0xD(184)(3);
  VNStageIntLLRInputS0xD(272)(3) <= CNStageIntLLROutputS0xD(184)(4);
  VNStageIntLLRInputS0xD(323)(2) <= CNStageIntLLROutputS0xD(184)(5);
  VNStageIntLLRInputS0xD(46)(3) <= CNStageIntLLROutputS0xD(185)(0);
  VNStageIntLLRInputS0xD(77)(1) <= CNStageIntLLROutputS0xD(185)(1);
  VNStageIntLLRInputS0xD(191)(3) <= CNStageIntLLROutputS0xD(185)(2);
  VNStageIntLLRInputS0xD(246)(3) <= CNStageIntLLROutputS0xD(185)(3);
  VNStageIntLLRInputS0xD(277)(3) <= CNStageIntLLROutputS0xD(185)(4);
  VNStageIntLLRInputS0xD(325)(3) <= CNStageIntLLROutputS0xD(185)(5);
  VNStageIntLLRInputS0xD(45)(3) <= CNStageIntLLROutputS0xD(186)(0);
  VNStageIntLLRInputS0xD(126)(2) <= CNStageIntLLROutputS0xD(186)(1);
  VNStageIntLLRInputS0xD(181)(3) <= CNStageIntLLROutputS0xD(186)(2);
  VNStageIntLLRInputS0xD(212)(3) <= CNStageIntLLROutputS0xD(186)(3);
  VNStageIntLLRInputS0xD(260)(3) <= CNStageIntLLROutputS0xD(186)(4);
  VNStageIntLLRInputS0xD(355)(3) <= CNStageIntLLROutputS0xD(186)(5);
  VNStageIntLLRInputS0xD(44)(3) <= CNStageIntLLROutputS0xD(187)(0);
  VNStageIntLLRInputS0xD(116)(2) <= CNStageIntLLROutputS0xD(187)(1);
  VNStageIntLLRInputS0xD(147)(3) <= CNStageIntLLROutputS0xD(187)(2);
  VNStageIntLLRInputS0xD(195)(2) <= CNStageIntLLROutputS0xD(187)(3);
  VNStageIntLLRInputS0xD(290)(3) <= CNStageIntLLROutputS0xD(187)(4);
  VNStageIntLLRInputS0xD(378)(2) <= CNStageIntLLROutputS0xD(187)(5);
  VNStageIntLLRInputS0xD(43)(2) <= CNStageIntLLROutputS0xD(188)(0);
  VNStageIntLLRInputS0xD(82)(3) <= CNStageIntLLROutputS0xD(188)(1);
  VNStageIntLLRInputS0xD(130)(3) <= CNStageIntLLROutputS0xD(188)(2);
  VNStageIntLLRInputS0xD(225)(3) <= CNStageIntLLROutputS0xD(188)(3);
  VNStageIntLLRInputS0xD(313)(1) <= CNStageIntLLROutputS0xD(188)(4);
  VNStageIntLLRInputS0xD(351)(2) <= CNStageIntLLROutputS0xD(188)(5);
  VNStageIntLLRInputS0xD(42)(3) <= CNStageIntLLROutputS0xD(189)(0);
  VNStageIntLLRInputS0xD(65)(3) <= CNStageIntLLROutputS0xD(189)(1);
  VNStageIntLLRInputS0xD(160)(3) <= CNStageIntLLROutputS0xD(189)(2);
  VNStageIntLLRInputS0xD(248)(3) <= CNStageIntLLROutputS0xD(189)(3);
  VNStageIntLLRInputS0xD(286)(3) <= CNStageIntLLROutputS0xD(189)(4);
  VNStageIntLLRInputS0xD(335)(3) <= CNStageIntLLROutputS0xD(189)(5);
  VNStageIntLLRInputS0xD(41)(3) <= CNStageIntLLROutputS0xD(190)(0);
  VNStageIntLLRInputS0xD(95)(3) <= CNStageIntLLROutputS0xD(190)(1);
  VNStageIntLLRInputS0xD(183)(2) <= CNStageIntLLROutputS0xD(190)(2);
  VNStageIntLLRInputS0xD(221)(3) <= CNStageIntLLROutputS0xD(190)(3);
  VNStageIntLLRInputS0xD(270)(3) <= CNStageIntLLROutputS0xD(190)(4);
  VNStageIntLLRInputS0xD(338)(3) <= CNStageIntLLROutputS0xD(190)(5);
  VNStageIntLLRInputS0xD(39)(3) <= CNStageIntLLROutputS0xD(191)(0);
  VNStageIntLLRInputS0xD(91)(3) <= CNStageIntLLROutputS0xD(191)(1);
  VNStageIntLLRInputS0xD(140)(3) <= CNStageIntLLROutputS0xD(191)(2);
  VNStageIntLLRInputS0xD(208)(3) <= CNStageIntLLROutputS0xD(191)(3);
  VNStageIntLLRInputS0xD(314)(0) <= CNStageIntLLROutputS0xD(191)(4);
  VNStageIntLLRInputS0xD(354)(3) <= CNStageIntLLROutputS0xD(191)(5);
  VNStageIntLLRInputS0xD(38)(3) <= CNStageIntLLROutputS0xD(192)(0);
  VNStageIntLLRInputS0xD(75)(3) <= CNStageIntLLROutputS0xD(192)(1);
  VNStageIntLLRInputS0xD(143)(3) <= CNStageIntLLROutputS0xD(192)(2);
  VNStageIntLLRInputS0xD(249)(1) <= CNStageIntLLROutputS0xD(192)(3);
  VNStageIntLLRInputS0xD(289)(3) <= CNStageIntLLROutputS0xD(192)(4);
  VNStageIntLLRInputS0xD(352)(3) <= CNStageIntLLROutputS0xD(192)(5);
  VNStageIntLLRInputS0xD(37)(3) <= CNStageIntLLROutputS0xD(193)(0);
  VNStageIntLLRInputS0xD(78)(3) <= CNStageIntLLROutputS0xD(193)(1);
  VNStageIntLLRInputS0xD(184)(3) <= CNStageIntLLROutputS0xD(193)(2);
  VNStageIntLLRInputS0xD(224)(3) <= CNStageIntLLROutputS0xD(193)(3);
  VNStageIntLLRInputS0xD(287)(3) <= CNStageIntLLROutputS0xD(193)(4);
  VNStageIntLLRInputS0xD(377)(2) <= CNStageIntLLROutputS0xD(193)(5);
  VNStageIntLLRInputS0xD(35)(3) <= CNStageIntLLROutputS0xD(194)(0);
  VNStageIntLLRInputS0xD(94)(2) <= CNStageIntLLROutputS0xD(194)(1);
  VNStageIntLLRInputS0xD(157)(3) <= CNStageIntLLROutputS0xD(194)(2);
  VNStageIntLLRInputS0xD(247)(3) <= CNStageIntLLROutputS0xD(194)(3);
  VNStageIntLLRInputS0xD(257)(3) <= CNStageIntLLROutputS0xD(194)(4);
  VNStageIntLLRInputS0xD(365)(3) <= CNStageIntLLROutputS0xD(194)(5);
  VNStageIntLLRInputS0xD(34)(3) <= CNStageIntLLROutputS0xD(195)(0);
  VNStageIntLLRInputS0xD(92)(3) <= CNStageIntLLROutputS0xD(195)(1);
  VNStageIntLLRInputS0xD(182)(3) <= CNStageIntLLROutputS0xD(195)(2);
  VNStageIntLLRInputS0xD(255)(3) <= CNStageIntLLROutputS0xD(195)(3);
  VNStageIntLLRInputS0xD(300)(3) <= CNStageIntLLROutputS0xD(195)(4);
  VNStageIntLLRInputS0xD(359)(3) <= CNStageIntLLROutputS0xD(195)(5);
  VNStageIntLLRInputS0xD(33)(3) <= CNStageIntLLROutputS0xD(196)(0);
  VNStageIntLLRInputS0xD(117)(3) <= CNStageIntLLROutputS0xD(196)(1);
  VNStageIntLLRInputS0xD(190)(1) <= CNStageIntLLROutputS0xD(196)(2);
  VNStageIntLLRInputS0xD(235)(2) <= CNStageIntLLROutputS0xD(196)(3);
  VNStageIntLLRInputS0xD(294)(3) <= CNStageIntLLROutputS0xD(196)(4);
  VNStageIntLLRInputS0xD(320)(2) <= CNStageIntLLROutputS0xD(196)(5);
  VNStageIntLLRInputS0xD(31)(2) <= CNStageIntLLROutputS0xD(197)(0);
  VNStageIntLLRInputS0xD(105)(2) <= CNStageIntLLROutputS0xD(197)(1);
  VNStageIntLLRInputS0xD(164)(3) <= CNStageIntLLROutputS0xD(197)(2);
  VNStageIntLLRInputS0xD(192)(3) <= CNStageIntLLROutputS0xD(197)(3);
  VNStageIntLLRInputS0xD(293)(3) <= CNStageIntLLROutputS0xD(197)(4);
  VNStageIntLLRInputS0xD(363)(2) <= CNStageIntLLROutputS0xD(197)(5);
  VNStageIntLLRInputS0xD(30)(3) <= CNStageIntLLROutputS0xD(198)(0);
  VNStageIntLLRInputS0xD(99)(3) <= CNStageIntLLROutputS0xD(198)(1);
  VNStageIntLLRInputS0xD(128)(3) <= CNStageIntLLROutputS0xD(198)(2);
  VNStageIntLLRInputS0xD(228)(3) <= CNStageIntLLROutputS0xD(198)(3);
  VNStageIntLLRInputS0xD(298)(3) <= CNStageIntLLROutputS0xD(198)(4);
  VNStageIntLLRInputS0xD(382)(2) <= CNStageIntLLROutputS0xD(198)(5);
  VNStageIntLLRInputS0xD(28)(3) <= CNStageIntLLROutputS0xD(199)(0);
  VNStageIntLLRInputS0xD(98)(2) <= CNStageIntLLROutputS0xD(199)(1);
  VNStageIntLLRInputS0xD(168)(2) <= CNStageIntLLROutputS0xD(199)(2);
  VNStageIntLLRInputS0xD(252)(2) <= CNStageIntLLROutputS0xD(199)(3);
  VNStageIntLLRInputS0xD(308)(1) <= CNStageIntLLROutputS0xD(199)(4);
  VNStageIntLLRInputS0xD(347)(3) <= CNStageIntLLROutputS0xD(199)(5);
  VNStageIntLLRInputS0xD(27)(3) <= CNStageIntLLROutputS0xD(200)(0);
  VNStageIntLLRInputS0xD(103)(3) <= CNStageIntLLROutputS0xD(200)(1);
  VNStageIntLLRInputS0xD(187)(2) <= CNStageIntLLROutputS0xD(200)(2);
  VNStageIntLLRInputS0xD(243)(3) <= CNStageIntLLROutputS0xD(200)(3);
  VNStageIntLLRInputS0xD(282)(3) <= CNStageIntLLROutputS0xD(200)(4);
  VNStageIntLLRInputS0xD(348)(3) <= CNStageIntLLROutputS0xD(200)(5);
  VNStageIntLLRInputS0xD(26)(3) <= CNStageIntLLROutputS0xD(201)(0);
  VNStageIntLLRInputS0xD(122)(2) <= CNStageIntLLROutputS0xD(201)(1);
  VNStageIntLLRInputS0xD(178)(3) <= CNStageIntLLROutputS0xD(201)(2);
  VNStageIntLLRInputS0xD(217)(3) <= CNStageIntLLROutputS0xD(201)(3);
  VNStageIntLLRInputS0xD(283)(3) <= CNStageIntLLROutputS0xD(201)(4);
  VNStageIntLLRInputS0xD(372)(2) <= CNStageIntLLROutputS0xD(201)(5);
  VNStageIntLLRInputS0xD(25)(3) <= CNStageIntLLROutputS0xD(202)(0);
  VNStageIntLLRInputS0xD(113)(3) <= CNStageIntLLROutputS0xD(202)(1);
  VNStageIntLLRInputS0xD(152)(3) <= CNStageIntLLROutputS0xD(202)(2);
  VNStageIntLLRInputS0xD(218)(3) <= CNStageIntLLROutputS0xD(202)(3);
  VNStageIntLLRInputS0xD(307)(3) <= CNStageIntLLROutputS0xD(202)(4);
  VNStageIntLLRInputS0xD(330)(3) <= CNStageIntLLROutputS0xD(202)(5);
  VNStageIntLLRInputS0xD(24)(3) <= CNStageIntLLROutputS0xD(203)(0);
  VNStageIntLLRInputS0xD(87)(3) <= CNStageIntLLROutputS0xD(203)(1);
  VNStageIntLLRInputS0xD(153)(3) <= CNStageIntLLROutputS0xD(203)(2);
  VNStageIntLLRInputS0xD(242)(3) <= CNStageIntLLROutputS0xD(203)(3);
  VNStageIntLLRInputS0xD(265)(2) <= CNStageIntLLROutputS0xD(203)(4);
  VNStageIntLLRInputS0xD(326)(2) <= CNStageIntLLROutputS0xD(203)(5);
  VNStageIntLLRInputS0xD(23)(3) <= CNStageIntLLROutputS0xD(204)(0);
  VNStageIntLLRInputS0xD(88)(3) <= CNStageIntLLROutputS0xD(204)(1);
  VNStageIntLLRInputS0xD(177)(3) <= CNStageIntLLROutputS0xD(204)(2);
  VNStageIntLLRInputS0xD(200)(3) <= CNStageIntLLROutputS0xD(204)(3);
  VNStageIntLLRInputS0xD(261)(3) <= CNStageIntLLROutputS0xD(204)(4);
  VNStageIntLLRInputS0xD(341)(3) <= CNStageIntLLROutputS0xD(204)(5);
  VNStageIntLLRInputS0xD(22)(3) <= CNStageIntLLROutputS0xD(205)(0);
  VNStageIntLLRInputS0xD(112)(3) <= CNStageIntLLROutputS0xD(205)(1);
  VNStageIntLLRInputS0xD(135)(3) <= CNStageIntLLROutputS0xD(205)(2);
  VNStageIntLLRInputS0xD(196)(3) <= CNStageIntLLROutputS0xD(205)(3);
  VNStageIntLLRInputS0xD(276)(3) <= CNStageIntLLROutputS0xD(205)(4);
  VNStageIntLLRInputS0xD(367)(3) <= CNStageIntLLROutputS0xD(205)(5);
  VNStageIntLLRInputS0xD(21)(3) <= CNStageIntLLROutputS0xD(206)(0);
  VNStageIntLLRInputS0xD(70)(3) <= CNStageIntLLROutputS0xD(206)(1);
  VNStageIntLLRInputS0xD(131)(2) <= CNStageIntLLROutputS0xD(206)(2);
  VNStageIntLLRInputS0xD(211)(3) <= CNStageIntLLROutputS0xD(206)(3);
  VNStageIntLLRInputS0xD(302)(3) <= CNStageIntLLROutputS0xD(206)(4);
  VNStageIntLLRInputS0xD(343)(3) <= CNStageIntLLROutputS0xD(206)(5);
  VNStageIntLLRInputS0xD(18)(3) <= CNStageIntLLROutputS0xD(207)(0);
  VNStageIntLLRInputS0xD(107)(2) <= CNStageIntLLROutputS0xD(207)(1);
  VNStageIntLLRInputS0xD(148)(3) <= CNStageIntLLROutputS0xD(207)(2);
  VNStageIntLLRInputS0xD(245)(3) <= CNStageIntLLROutputS0xD(207)(3);
  VNStageIntLLRInputS0xD(263)(3) <= CNStageIntLLROutputS0xD(207)(4);
  VNStageIntLLRInputS0xD(361)(3) <= CNStageIntLLROutputS0xD(207)(5);
  VNStageIntLLRInputS0xD(17)(3) <= CNStageIntLLROutputS0xD(208)(0);
  VNStageIntLLRInputS0xD(83)(3) <= CNStageIntLLROutputS0xD(208)(1);
  VNStageIntLLRInputS0xD(180)(1) <= CNStageIntLLROutputS0xD(208)(2);
  VNStageIntLLRInputS0xD(198)(3) <= CNStageIntLLROutputS0xD(208)(3);
  VNStageIntLLRInputS0xD(296)(3) <= CNStageIntLLROutputS0xD(208)(4);
  VNStageIntLLRInputS0xD(370)(2) <= CNStageIntLLROutputS0xD(208)(5);
  VNStageIntLLRInputS0xD(16)(2) <= CNStageIntLLROutputS0xD(209)(0);
  VNStageIntLLRInputS0xD(115)(3) <= CNStageIntLLROutputS0xD(209)(1);
  VNStageIntLLRInputS0xD(133)(1) <= CNStageIntLLROutputS0xD(209)(2);
  VNStageIntLLRInputS0xD(231)(2) <= CNStageIntLLROutputS0xD(209)(3);
  VNStageIntLLRInputS0xD(305)(3) <= CNStageIntLLROutputS0xD(209)(4);
  VNStageIntLLRInputS0xD(383)(3) <= CNStageIntLLROutputS0xD(209)(5);
  VNStageIntLLRInputS0xD(15)(3) <= CNStageIntLLROutputS0xD(210)(0);
  VNStageIntLLRInputS0xD(68)(2) <= CNStageIntLLROutputS0xD(210)(1);
  VNStageIntLLRInputS0xD(166)(3) <= CNStageIntLLROutputS0xD(210)(2);
  VNStageIntLLRInputS0xD(240)(3) <= CNStageIntLLROutputS0xD(210)(3);
  VNStageIntLLRInputS0xD(318)(1) <= CNStageIntLLROutputS0xD(210)(4);
  VNStageIntLLRInputS0xD(362)(3) <= CNStageIntLLROutputS0xD(210)(5);
  VNStageIntLLRInputS0xD(14)(3) <= CNStageIntLLROutputS0xD(211)(0);
  VNStageIntLLRInputS0xD(101)(3) <= CNStageIntLLROutputS0xD(211)(1);
  VNStageIntLLRInputS0xD(175)(3) <= CNStageIntLLROutputS0xD(211)(2);
  VNStageIntLLRInputS0xD(253)(2) <= CNStageIntLLROutputS0xD(211)(3);
  VNStageIntLLRInputS0xD(297)(3) <= CNStageIntLLROutputS0xD(211)(4);
  VNStageIntLLRInputS0xD(327)(3) <= CNStageIntLLROutputS0xD(211)(5);
  VNStageIntLLRInputS0xD(13)(2) <= CNStageIntLLROutputS0xD(212)(0);
  VNStageIntLLRInputS0xD(110)(3) <= CNStageIntLLROutputS0xD(212)(1);
  VNStageIntLLRInputS0xD(188)(1) <= CNStageIntLLROutputS0xD(212)(2);
  VNStageIntLLRInputS0xD(232)(2) <= CNStageIntLLROutputS0xD(212)(3);
  VNStageIntLLRInputS0xD(262)(3) <= CNStageIntLLROutputS0xD(212)(4);
  VNStageIntLLRInputS0xD(329)(3) <= CNStageIntLLROutputS0xD(212)(5);
  VNStageIntLLRInputS0xD(12)(3) <= CNStageIntLLROutputS0xD(213)(0);
  VNStageIntLLRInputS0xD(123)(2) <= CNStageIntLLROutputS0xD(213)(1);
  VNStageIntLLRInputS0xD(167)(3) <= CNStageIntLLROutputS0xD(213)(2);
  VNStageIntLLRInputS0xD(197)(3) <= CNStageIntLLROutputS0xD(213)(3);
  VNStageIntLLRInputS0xD(264)(3) <= CNStageIntLLROutputS0xD(213)(4);
  VNStageIntLLRInputS0xD(374)(3) <= CNStageIntLLROutputS0xD(213)(5);
  VNStageIntLLRInputS0xD(11)(3) <= CNStageIntLLROutputS0xD(214)(0);
  VNStageIntLLRInputS0xD(102)(3) <= CNStageIntLLROutputS0xD(214)(1);
  VNStageIntLLRInputS0xD(132)(2) <= CNStageIntLLROutputS0xD(214)(2);
  VNStageIntLLRInputS0xD(199)(3) <= CNStageIntLLROutputS0xD(214)(3);
  VNStageIntLLRInputS0xD(309)(3) <= CNStageIntLLROutputS0xD(214)(4);
  VNStageIntLLRInputS0xD(381)(2) <= CNStageIntLLROutputS0xD(214)(5);
  VNStageIntLLRInputS0xD(9)(3) <= CNStageIntLLROutputS0xD(215)(0);
  VNStageIntLLRInputS0xD(69)(3) <= CNStageIntLLROutputS0xD(215)(1);
  VNStageIntLLRInputS0xD(179)(3) <= CNStageIntLLROutputS0xD(215)(2);
  VNStageIntLLRInputS0xD(251)(2) <= CNStageIntLLROutputS0xD(215)(3);
  VNStageIntLLRInputS0xD(280)(3) <= CNStageIntLLROutputS0xD(215)(4);
  VNStageIntLLRInputS0xD(333)(2) <= CNStageIntLLROutputS0xD(215)(5);
  VNStageIntLLRInputS0xD(8)(2) <= CNStageIntLLROutputS0xD(216)(0);
  VNStageIntLLRInputS0xD(114)(3) <= CNStageIntLLROutputS0xD(216)(1);
  VNStageIntLLRInputS0xD(186)(2) <= CNStageIntLLROutputS0xD(216)(2);
  VNStageIntLLRInputS0xD(215)(3) <= CNStageIntLLROutputS0xD(216)(3);
  VNStageIntLLRInputS0xD(268)(3) <= CNStageIntLLROutputS0xD(216)(4);
  VNStageIntLLRInputS0xD(339)(3) <= CNStageIntLLROutputS0xD(216)(5);
  VNStageIntLLRInputS0xD(7)(3) <= CNStageIntLLROutputS0xD(217)(0);
  VNStageIntLLRInputS0xD(121)(2) <= CNStageIntLLROutputS0xD(217)(1);
  VNStageIntLLRInputS0xD(150)(3) <= CNStageIntLLROutputS0xD(217)(2);
  VNStageIntLLRInputS0xD(203)(3) <= CNStageIntLLROutputS0xD(217)(3);
  VNStageIntLLRInputS0xD(274)(2) <= CNStageIntLLROutputS0xD(217)(4);
  VNStageIntLLRInputS0xD(334)(2) <= CNStageIntLLROutputS0xD(217)(5);
  VNStageIntLLRInputS0xD(6)(3) <= CNStageIntLLROutputS0xD(218)(0);
  VNStageIntLLRInputS0xD(85)(2) <= CNStageIntLLROutputS0xD(218)(1);
  VNStageIntLLRInputS0xD(138)(3) <= CNStageIntLLROutputS0xD(218)(2);
  VNStageIntLLRInputS0xD(209)(3) <= CNStageIntLLROutputS0xD(218)(3);
  VNStageIntLLRInputS0xD(269)(2) <= CNStageIntLLROutputS0xD(218)(4);
  VNStageIntLLRInputS0xD(344)(3) <= CNStageIntLLROutputS0xD(218)(5);
  VNStageIntLLRInputS0xD(5)(3) <= CNStageIntLLROutputS0xD(219)(0);
  VNStageIntLLRInputS0xD(73)(3) <= CNStageIntLLROutputS0xD(219)(1);
  VNStageIntLLRInputS0xD(144)(3) <= CNStageIntLLROutputS0xD(219)(2);
  VNStageIntLLRInputS0xD(204)(3) <= CNStageIntLLROutputS0xD(219)(3);
  VNStageIntLLRInputS0xD(279)(3) <= CNStageIntLLROutputS0xD(219)(4);
  VNStageIntLLRInputS0xD(366)(3) <= CNStageIntLLROutputS0xD(219)(5);
  VNStageIntLLRInputS0xD(4)(2) <= CNStageIntLLROutputS0xD(220)(0);
  VNStageIntLLRInputS0xD(79)(3) <= CNStageIntLLROutputS0xD(220)(1);
  VNStageIntLLRInputS0xD(139)(3) <= CNStageIntLLROutputS0xD(220)(2);
  VNStageIntLLRInputS0xD(214)(3) <= CNStageIntLLROutputS0xD(220)(3);
  VNStageIntLLRInputS0xD(301)(3) <= CNStageIntLLROutputS0xD(220)(4);
  VNStageIntLLRInputS0xD(321)(3) <= CNStageIntLLROutputS0xD(220)(5);
  VNStageIntLLRInputS0xD(3)(2) <= CNStageIntLLROutputS0xD(221)(0);
  VNStageIntLLRInputS0xD(74)(3) <= CNStageIntLLROutputS0xD(221)(1);
  VNStageIntLLRInputS0xD(149)(3) <= CNStageIntLLROutputS0xD(221)(2);
  VNStageIntLLRInputS0xD(236)(3) <= CNStageIntLLROutputS0xD(221)(3);
  VNStageIntLLRInputS0xD(319)(3) <= CNStageIntLLROutputS0xD(221)(4);
  VNStageIntLLRInputS0xD(369)(2) <= CNStageIntLLROutputS0xD(221)(5);
  VNStageIntLLRInputS0xD(2)(3) <= CNStageIntLLROutputS0xD(222)(0);
  VNStageIntLLRInputS0xD(84)(3) <= CNStageIntLLROutputS0xD(222)(1);
  VNStageIntLLRInputS0xD(171)(2) <= CNStageIntLLROutputS0xD(222)(2);
  VNStageIntLLRInputS0xD(254)(1) <= CNStageIntLLROutputS0xD(222)(3);
  VNStageIntLLRInputS0xD(304)(3) <= CNStageIntLLROutputS0xD(222)(4);
  VNStageIntLLRInputS0xD(356)(3) <= CNStageIntLLROutputS0xD(222)(5);
  VNStageIntLLRInputS0xD(1)(2) <= CNStageIntLLROutputS0xD(223)(0);
  VNStageIntLLRInputS0xD(106)(2) <= CNStageIntLLROutputS0xD(223)(1);
  VNStageIntLLRInputS0xD(189)(2) <= CNStageIntLLROutputS0xD(223)(2);
  VNStageIntLLRInputS0xD(239)(3) <= CNStageIntLLROutputS0xD(223)(3);
  VNStageIntLLRInputS0xD(291)(3) <= CNStageIntLLROutputS0xD(223)(4);
  VNStageIntLLRInputS0xD(324)(3) <= CNStageIntLLROutputS0xD(223)(5);
  VNStageIntLLRInputS0xD(0)(3) <= CNStageIntLLROutputS0xD(224)(0);
  VNStageIntLLRInputS0xD(93)(3) <= CNStageIntLLROutputS0xD(224)(1);
  VNStageIntLLRInputS0xD(158)(3) <= CNStageIntLLROutputS0xD(224)(2);
  VNStageIntLLRInputS0xD(223)(3) <= CNStageIntLLROutputS0xD(224)(3);
  VNStageIntLLRInputS0xD(288)(3) <= CNStageIntLLROutputS0xD(224)(4);
  VNStageIntLLRInputS0xD(353)(3) <= CNStageIntLLROutputS0xD(224)(5);
  VNStageIntLLRInputS0xD(18)(4) <= CNStageIntLLROutputS0xD(225)(0);
  VNStageIntLLRInputS0xD(110)(4) <= CNStageIntLLROutputS0xD(225)(1);
  VNStageIntLLRInputS0xD(167)(4) <= CNStageIntLLROutputS0xD(225)(2);
  VNStageIntLLRInputS0xD(249)(2) <= CNStageIntLLROutputS0xD(225)(3);
  VNStageIntLLRInputS0xD(311)(3) <= CNStageIntLLROutputS0xD(225)(4);
  VNStageIntLLRInputS0xD(347)(4) <= CNStageIntLLROutputS0xD(225)(5);
  VNStageIntLLRInputS0xD(17)(4) <= CNStageIntLLROutputS0xD(226)(0);
  VNStageIntLLRInputS0xD(102)(4) <= CNStageIntLLROutputS0xD(226)(1);
  VNStageIntLLRInputS0xD(184)(4) <= CNStageIntLLROutputS0xD(226)(2);
  VNStageIntLLRInputS0xD(246)(4) <= CNStageIntLLROutputS0xD(226)(3);
  VNStageIntLLRInputS0xD(282)(4) <= CNStageIntLLROutputS0xD(226)(4);
  VNStageIntLLRInputS0xD(367)(4) <= CNStageIntLLROutputS0xD(226)(5);
  VNStageIntLLRInputS0xD(16)(3) <= CNStageIntLLROutputS0xD(227)(0);
  VNStageIntLLRInputS0xD(119)(3) <= CNStageIntLLROutputS0xD(227)(1);
  VNStageIntLLRInputS0xD(181)(4) <= CNStageIntLLROutputS0xD(227)(2);
  VNStageIntLLRInputS0xD(217)(4) <= CNStageIntLLROutputS0xD(227)(3);
  VNStageIntLLRInputS0xD(302)(4) <= CNStageIntLLROutputS0xD(227)(4);
  VNStageIntLLRInputS0xD(353)(4) <= CNStageIntLLROutputS0xD(227)(5);
  VNStageIntLLRInputS0xD(15)(4) <= CNStageIntLLROutputS0xD(228)(0);
  VNStageIntLLRInputS0xD(116)(3) <= CNStageIntLLROutputS0xD(228)(1);
  VNStageIntLLRInputS0xD(152)(4) <= CNStageIntLLROutputS0xD(228)(2);
  VNStageIntLLRInputS0xD(237)(3) <= CNStageIntLLROutputS0xD(228)(3);
  VNStageIntLLRInputS0xD(288)(4) <= CNStageIntLLROutputS0xD(228)(4);
  VNStageIntLLRInputS0xD(343)(4) <= CNStageIntLLROutputS0xD(228)(5);
  VNStageIntLLRInputS0xD(14)(4) <= CNStageIntLLROutputS0xD(229)(0);
  VNStageIntLLRInputS0xD(87)(4) <= CNStageIntLLROutputS0xD(229)(1);
  VNStageIntLLRInputS0xD(172)(3) <= CNStageIntLLROutputS0xD(229)(2);
  VNStageIntLLRInputS0xD(223)(4) <= CNStageIntLLROutputS0xD(229)(3);
  VNStageIntLLRInputS0xD(278)(3) <= CNStageIntLLROutputS0xD(229)(4);
  VNStageIntLLRInputS0xD(372)(3) <= CNStageIntLLROutputS0xD(229)(5);
  VNStageIntLLRInputS0xD(13)(3) <= CNStageIntLLROutputS0xD(230)(0);
  VNStageIntLLRInputS0xD(107)(3) <= CNStageIntLLROutputS0xD(230)(1);
  VNStageIntLLRInputS0xD(158)(4) <= CNStageIntLLROutputS0xD(230)(2);
  VNStageIntLLRInputS0xD(213)(3) <= CNStageIntLLROutputS0xD(230)(3);
  VNStageIntLLRInputS0xD(307)(4) <= CNStageIntLLROutputS0xD(230)(4);
  VNStageIntLLRInputS0xD(355)(4) <= CNStageIntLLROutputS0xD(230)(5);
  VNStageIntLLRInputS0xD(12)(4) <= CNStageIntLLROutputS0xD(231)(0);
  VNStageIntLLRInputS0xD(93)(4) <= CNStageIntLLROutputS0xD(231)(1);
  VNStageIntLLRInputS0xD(148)(4) <= CNStageIntLLROutputS0xD(231)(2);
  VNStageIntLLRInputS0xD(242)(4) <= CNStageIntLLROutputS0xD(231)(3);
  VNStageIntLLRInputS0xD(290)(4) <= CNStageIntLLROutputS0xD(231)(4);
  VNStageIntLLRInputS0xD(322)(3) <= CNStageIntLLROutputS0xD(231)(5);
  VNStageIntLLRInputS0xD(11)(4) <= CNStageIntLLROutputS0xD(232)(0);
  VNStageIntLLRInputS0xD(83)(4) <= CNStageIntLLROutputS0xD(232)(1);
  VNStageIntLLRInputS0xD(177)(4) <= CNStageIntLLROutputS0xD(232)(2);
  VNStageIntLLRInputS0xD(225)(4) <= CNStageIntLLROutputS0xD(232)(3);
  VNStageIntLLRInputS0xD(257)(4) <= CNStageIntLLROutputS0xD(232)(4);
  VNStageIntLLRInputS0xD(345)(3) <= CNStageIntLLROutputS0xD(232)(5);
  VNStageIntLLRInputS0xD(10)(3) <= CNStageIntLLROutputS0xD(233)(0);
  VNStageIntLLRInputS0xD(112)(4) <= CNStageIntLLROutputS0xD(233)(1);
  VNStageIntLLRInputS0xD(160)(4) <= CNStageIntLLROutputS0xD(233)(2);
  VNStageIntLLRInputS0xD(255)(4) <= CNStageIntLLROutputS0xD(233)(3);
  VNStageIntLLRInputS0xD(280)(4) <= CNStageIntLLROutputS0xD(233)(4);
  VNStageIntLLRInputS0xD(381)(3) <= CNStageIntLLROutputS0xD(233)(5);
  VNStageIntLLRInputS0xD(9)(4) <= CNStageIntLLROutputS0xD(234)(0);
  VNStageIntLLRInputS0xD(95)(4) <= CNStageIntLLROutputS0xD(234)(1);
  VNStageIntLLRInputS0xD(190)(2) <= CNStageIntLLROutputS0xD(234)(2);
  VNStageIntLLRInputS0xD(215)(4) <= CNStageIntLLROutputS0xD(234)(3);
  VNStageIntLLRInputS0xD(316)(2) <= CNStageIntLLROutputS0xD(234)(4);
  VNStageIntLLRInputS0xD(365)(4) <= CNStageIntLLROutputS0xD(234)(5);
  VNStageIntLLRInputS0xD(7)(4) <= CNStageIntLLROutputS0xD(235)(0);
  VNStageIntLLRInputS0xD(85)(3) <= CNStageIntLLROutputS0xD(235)(1);
  VNStageIntLLRInputS0xD(186)(3) <= CNStageIntLLROutputS0xD(235)(2);
  VNStageIntLLRInputS0xD(235)(3) <= CNStageIntLLROutputS0xD(235)(3);
  VNStageIntLLRInputS0xD(303)(4) <= CNStageIntLLROutputS0xD(235)(4);
  VNStageIntLLRInputS0xD(346)(4) <= CNStageIntLLROutputS0xD(235)(5);
  VNStageIntLLRInputS0xD(6)(4) <= CNStageIntLLROutputS0xD(236)(0);
  VNStageIntLLRInputS0xD(121)(3) <= CNStageIntLLROutputS0xD(236)(1);
  VNStageIntLLRInputS0xD(170)(3) <= CNStageIntLLROutputS0xD(236)(2);
  VNStageIntLLRInputS0xD(238)(4) <= CNStageIntLLROutputS0xD(236)(3);
  VNStageIntLLRInputS0xD(281)(4) <= CNStageIntLLROutputS0xD(236)(4);
  VNStageIntLLRInputS0xD(321)(4) <= CNStageIntLLROutputS0xD(236)(5);
  VNStageIntLLRInputS0xD(5)(4) <= CNStageIntLLROutputS0xD(237)(0);
  VNStageIntLLRInputS0xD(105)(3) <= CNStageIntLLROutputS0xD(237)(1);
  VNStageIntLLRInputS0xD(173)(4) <= CNStageIntLLROutputS0xD(237)(2);
  VNStageIntLLRInputS0xD(216)(4) <= CNStageIntLLROutputS0xD(237)(3);
  VNStageIntLLRInputS0xD(319)(4) <= CNStageIntLLROutputS0xD(237)(4);
  VNStageIntLLRInputS0xD(382)(3) <= CNStageIntLLROutputS0xD(237)(5);
  VNStageIntLLRInputS0xD(4)(3) <= CNStageIntLLROutputS0xD(238)(0);
  VNStageIntLLRInputS0xD(108)(4) <= CNStageIntLLROutputS0xD(238)(1);
  VNStageIntLLRInputS0xD(151)(4) <= CNStageIntLLROutputS0xD(238)(2);
  VNStageIntLLRInputS0xD(254)(2) <= CNStageIntLLROutputS0xD(238)(3);
  VNStageIntLLRInputS0xD(317)(1) <= CNStageIntLLROutputS0xD(238)(4);
  VNStageIntLLRInputS0xD(344)(4) <= CNStageIntLLROutputS0xD(238)(5);
  VNStageIntLLRInputS0xD(3)(3) <= CNStageIntLLROutputS0xD(239)(0);
  VNStageIntLLRInputS0xD(86)(2) <= CNStageIntLLROutputS0xD(239)(1);
  VNStageIntLLRInputS0xD(189)(3) <= CNStageIntLLROutputS0xD(239)(2);
  VNStageIntLLRInputS0xD(252)(3) <= CNStageIntLLROutputS0xD(239)(3);
  VNStageIntLLRInputS0xD(279)(4) <= CNStageIntLLROutputS0xD(239)(4);
  VNStageIntLLRInputS0xD(352)(4) <= CNStageIntLLROutputS0xD(239)(5);
  VNStageIntLLRInputS0xD(2)(4) <= CNStageIntLLROutputS0xD(240)(0);
  VNStageIntLLRInputS0xD(124)(2) <= CNStageIntLLROutputS0xD(240)(1);
  VNStageIntLLRInputS0xD(187)(3) <= CNStageIntLLROutputS0xD(240)(2);
  VNStageIntLLRInputS0xD(214)(4) <= CNStageIntLLROutputS0xD(240)(3);
  VNStageIntLLRInputS0xD(287)(4) <= CNStageIntLLROutputS0xD(240)(4);
  VNStageIntLLRInputS0xD(332)(4) <= CNStageIntLLROutputS0xD(240)(5);
  VNStageIntLLRInputS0xD(1)(3) <= CNStageIntLLROutputS0xD(241)(0);
  VNStageIntLLRInputS0xD(122)(3) <= CNStageIntLLROutputS0xD(241)(1);
  VNStageIntLLRInputS0xD(149)(4) <= CNStageIntLLROutputS0xD(241)(2);
  VNStageIntLLRInputS0xD(222)(2) <= CNStageIntLLROutputS0xD(241)(3);
  VNStageIntLLRInputS0xD(267)(4) <= CNStageIntLLROutputS0xD(241)(4);
  VNStageIntLLRInputS0xD(326)(3) <= CNStageIntLLROutputS0xD(241)(5);
  VNStageIntLLRInputS0xD(62)(3) <= CNStageIntLLROutputS0xD(242)(0);
  VNStageIntLLRInputS0xD(92)(4) <= CNStageIntLLROutputS0xD(242)(1);
  VNStageIntLLRInputS0xD(137)(4) <= CNStageIntLLROutputS0xD(242)(2);
  VNStageIntLLRInputS0xD(196)(4) <= CNStageIntLLROutputS0xD(242)(3);
  VNStageIntLLRInputS0xD(256)(3) <= CNStageIntLLROutputS0xD(242)(4);
  VNStageIntLLRInputS0xD(325)(4) <= CNStageIntLLROutputS0xD(242)(5);
  VNStageIntLLRInputS0xD(61)(3) <= CNStageIntLLROutputS0xD(243)(0);
  VNStageIntLLRInputS0xD(72)(4) <= CNStageIntLLROutputS0xD(243)(1);
  VNStageIntLLRInputS0xD(131)(3) <= CNStageIntLLROutputS0xD(243)(2);
  VNStageIntLLRInputS0xD(192)(4) <= CNStageIntLLROutputS0xD(243)(3);
  VNStageIntLLRInputS0xD(260)(4) <= CNStageIntLLROutputS0xD(243)(4);
  VNStageIntLLRInputS0xD(330)(4) <= CNStageIntLLROutputS0xD(243)(5);
  VNStageIntLLRInputS0xD(60)(3) <= CNStageIntLLROutputS0xD(244)(0);
  VNStageIntLLRInputS0xD(66)(3) <= CNStageIntLLROutputS0xD(244)(1);
  VNStageIntLLRInputS0xD(128)(4) <= CNStageIntLLROutputS0xD(244)(2);
  VNStageIntLLRInputS0xD(195)(3) <= CNStageIntLLROutputS0xD(244)(3);
  VNStageIntLLRInputS0xD(265)(3) <= CNStageIntLLROutputS0xD(244)(4);
  VNStageIntLLRInputS0xD(349)(3) <= CNStageIntLLROutputS0xD(244)(5);
  VNStageIntLLRInputS0xD(59)(2) <= CNStageIntLLROutputS0xD(245)(0);
  VNStageIntLLRInputS0xD(64)(3) <= CNStageIntLLROutputS0xD(245)(1);
  VNStageIntLLRInputS0xD(130)(4) <= CNStageIntLLROutputS0xD(245)(2);
  VNStageIntLLRInputS0xD(200)(4) <= CNStageIntLLROutputS0xD(245)(3);
  VNStageIntLLRInputS0xD(284)(4) <= CNStageIntLLROutputS0xD(245)(4);
  VNStageIntLLRInputS0xD(340)(4) <= CNStageIntLLROutputS0xD(245)(5);
  VNStageIntLLRInputS0xD(57)(3) <= CNStageIntLLROutputS0xD(246)(0);
  VNStageIntLLRInputS0xD(70)(4) <= CNStageIntLLROutputS0xD(246)(1);
  VNStageIntLLRInputS0xD(154)(3) <= CNStageIntLLROutputS0xD(246)(2);
  VNStageIntLLRInputS0xD(210)(4) <= CNStageIntLLROutputS0xD(246)(3);
  VNStageIntLLRInputS0xD(312)(3) <= CNStageIntLLROutputS0xD(246)(4);
  VNStageIntLLRInputS0xD(378)(3) <= CNStageIntLLROutputS0xD(246)(5);
  VNStageIntLLRInputS0xD(56)(4) <= CNStageIntLLROutputS0xD(247)(0);
  VNStageIntLLRInputS0xD(89)(4) <= CNStageIntLLROutputS0xD(247)(1);
  VNStageIntLLRInputS0xD(145)(4) <= CNStageIntLLROutputS0xD(247)(2);
  VNStageIntLLRInputS0xD(247)(4) <= CNStageIntLLROutputS0xD(247)(3);
  VNStageIntLLRInputS0xD(313)(2) <= CNStageIntLLROutputS0xD(247)(4);
  VNStageIntLLRInputS0xD(339)(4) <= CNStageIntLLROutputS0xD(247)(5);
  VNStageIntLLRInputS0xD(55)(4) <= CNStageIntLLROutputS0xD(248)(0);
  VNStageIntLLRInputS0xD(80)(4) <= CNStageIntLLROutputS0xD(248)(1);
  VNStageIntLLRInputS0xD(182)(4) <= CNStageIntLLROutputS0xD(248)(2);
  VNStageIntLLRInputS0xD(248)(4) <= CNStageIntLLROutputS0xD(248)(3);
  VNStageIntLLRInputS0xD(274)(3) <= CNStageIntLLROutputS0xD(248)(4);
  VNStageIntLLRInputS0xD(360)(4) <= CNStageIntLLROutputS0xD(248)(5);
  VNStageIntLLRInputS0xD(53)(3) <= CNStageIntLLROutputS0xD(249)(0);
  VNStageIntLLRInputS0xD(118)(3) <= CNStageIntLLROutputS0xD(249)(1);
  VNStageIntLLRInputS0xD(144)(4) <= CNStageIntLLROutputS0xD(249)(2);
  VNStageIntLLRInputS0xD(230)(3) <= CNStageIntLLROutputS0xD(249)(3);
  VNStageIntLLRInputS0xD(291)(4) <= CNStageIntLLROutputS0xD(249)(4);
  VNStageIntLLRInputS0xD(371)(3) <= CNStageIntLLROutputS0xD(249)(5);
  VNStageIntLLRInputS0xD(51)(3) <= CNStageIntLLROutputS0xD(250)(0);
  VNStageIntLLRInputS0xD(100)(4) <= CNStageIntLLROutputS0xD(250)(1);
  VNStageIntLLRInputS0xD(161)(4) <= CNStageIntLLROutputS0xD(250)(2);
  VNStageIntLLRInputS0xD(241)(3) <= CNStageIntLLROutputS0xD(250)(3);
  VNStageIntLLRInputS0xD(269)(3) <= CNStageIntLLROutputS0xD(250)(4);
  VNStageIntLLRInputS0xD(373)(2) <= CNStageIntLLROutputS0xD(250)(5);
  VNStageIntLLRInputS0xD(50)(4) <= CNStageIntLLROutputS0xD(251)(0);
  VNStageIntLLRInputS0xD(96)(4) <= CNStageIntLLROutputS0xD(251)(1);
  VNStageIntLLRInputS0xD(176)(4) <= CNStageIntLLROutputS0xD(251)(2);
  VNStageIntLLRInputS0xD(204)(4) <= CNStageIntLLROutputS0xD(251)(3);
  VNStageIntLLRInputS0xD(308)(2) <= CNStageIntLLROutputS0xD(251)(4);
  VNStageIntLLRInputS0xD(342)(3) <= CNStageIntLLROutputS0xD(251)(5);
  VNStageIntLLRInputS0xD(49)(4) <= CNStageIntLLROutputS0xD(252)(0);
  VNStageIntLLRInputS0xD(111)(4) <= CNStageIntLLROutputS0xD(252)(1);
  VNStageIntLLRInputS0xD(139)(4) <= CNStageIntLLROutputS0xD(252)(2);
  VNStageIntLLRInputS0xD(243)(4) <= CNStageIntLLROutputS0xD(252)(3);
  VNStageIntLLRInputS0xD(277)(4) <= CNStageIntLLROutputS0xD(252)(4);
  VNStageIntLLRInputS0xD(358)(3) <= CNStageIntLLROutputS0xD(252)(5);
  VNStageIntLLRInputS0xD(47)(2) <= CNStageIntLLROutputS0xD(253)(0);
  VNStageIntLLRInputS0xD(113)(4) <= CNStageIntLLROutputS0xD(253)(1);
  VNStageIntLLRInputS0xD(147)(4) <= CNStageIntLLROutputS0xD(253)(2);
  VNStageIntLLRInputS0xD(228)(4) <= CNStageIntLLROutputS0xD(253)(3);
  VNStageIntLLRInputS0xD(263)(4) <= CNStageIntLLROutputS0xD(253)(4);
  VNStageIntLLRInputS0xD(337)(4) <= CNStageIntLLROutputS0xD(253)(5);
  VNStageIntLLRInputS0xD(46)(4) <= CNStageIntLLROutputS0xD(254)(0);
  VNStageIntLLRInputS0xD(82)(4) <= CNStageIntLLROutputS0xD(254)(1);
  VNStageIntLLRInputS0xD(163)(3) <= CNStageIntLLROutputS0xD(254)(2);
  VNStageIntLLRInputS0xD(198)(4) <= CNStageIntLLROutputS0xD(254)(3);
  VNStageIntLLRInputS0xD(272)(4) <= CNStageIntLLROutputS0xD(254)(4);
  VNStageIntLLRInputS0xD(350)(4) <= CNStageIntLLROutputS0xD(254)(5);
  VNStageIntLLRInputS0xD(45)(4) <= CNStageIntLLROutputS0xD(255)(0);
  VNStageIntLLRInputS0xD(98)(3) <= CNStageIntLLROutputS0xD(255)(1);
  VNStageIntLLRInputS0xD(133)(2) <= CNStageIntLLROutputS0xD(255)(2);
  VNStageIntLLRInputS0xD(207)(3) <= CNStageIntLLROutputS0xD(255)(3);
  VNStageIntLLRInputS0xD(285)(4) <= CNStageIntLLROutputS0xD(255)(4);
  VNStageIntLLRInputS0xD(329)(4) <= CNStageIntLLROutputS0xD(255)(5);
  VNStageIntLLRInputS0xD(44)(4) <= CNStageIntLLROutputS0xD(256)(0);
  VNStageIntLLRInputS0xD(68)(3) <= CNStageIntLLROutputS0xD(256)(1);
  VNStageIntLLRInputS0xD(142)(3) <= CNStageIntLLROutputS0xD(256)(2);
  VNStageIntLLRInputS0xD(220)(4) <= CNStageIntLLROutputS0xD(256)(3);
  VNStageIntLLRInputS0xD(264)(4) <= CNStageIntLLROutputS0xD(256)(4);
  VNStageIntLLRInputS0xD(357)(4) <= CNStageIntLLROutputS0xD(256)(5);
  VNStageIntLLRInputS0xD(43)(3) <= CNStageIntLLROutputS0xD(257)(0);
  VNStageIntLLRInputS0xD(77)(2) <= CNStageIntLLROutputS0xD(257)(1);
  VNStageIntLLRInputS0xD(155)(4) <= CNStageIntLLROutputS0xD(257)(2);
  VNStageIntLLRInputS0xD(199)(4) <= CNStageIntLLROutputS0xD(257)(3);
  VNStageIntLLRInputS0xD(292)(4) <= CNStageIntLLROutputS0xD(257)(4);
  VNStageIntLLRInputS0xD(359)(4) <= CNStageIntLLROutputS0xD(257)(5);
  VNStageIntLLRInputS0xD(42)(4) <= CNStageIntLLROutputS0xD(258)(0);
  VNStageIntLLRInputS0xD(90)(4) <= CNStageIntLLROutputS0xD(258)(1);
  VNStageIntLLRInputS0xD(134)(3) <= CNStageIntLLROutputS0xD(258)(2);
  VNStageIntLLRInputS0xD(227)(4) <= CNStageIntLLROutputS0xD(258)(3);
  VNStageIntLLRInputS0xD(294)(4) <= CNStageIntLLROutputS0xD(258)(4);
  VNStageIntLLRInputS0xD(341)(4) <= CNStageIntLLROutputS0xD(258)(5);
  VNStageIntLLRInputS0xD(41)(4) <= CNStageIntLLROutputS0xD(259)(0);
  VNStageIntLLRInputS0xD(69)(4) <= CNStageIntLLROutputS0xD(259)(1);
  VNStageIntLLRInputS0xD(162)(4) <= CNStageIntLLROutputS0xD(259)(2);
  VNStageIntLLRInputS0xD(229)(3) <= CNStageIntLLROutputS0xD(259)(3);
  VNStageIntLLRInputS0xD(276)(4) <= CNStageIntLLROutputS0xD(259)(4);
  VNStageIntLLRInputS0xD(348)(4) <= CNStageIntLLROutputS0xD(259)(5);
  VNStageIntLLRInputS0xD(40)(3) <= CNStageIntLLROutputS0xD(260)(0);
  VNStageIntLLRInputS0xD(97)(4) <= CNStageIntLLROutputS0xD(260)(1);
  VNStageIntLLRInputS0xD(164)(4) <= CNStageIntLLROutputS0xD(260)(2);
  VNStageIntLLRInputS0xD(211)(4) <= CNStageIntLLROutputS0xD(260)(3);
  VNStageIntLLRInputS0xD(283)(4) <= CNStageIntLLROutputS0xD(260)(4);
  VNStageIntLLRInputS0xD(375)(3) <= CNStageIntLLROutputS0xD(260)(5);
  VNStageIntLLRInputS0xD(39)(4) <= CNStageIntLLROutputS0xD(261)(0);
  VNStageIntLLRInputS0xD(99)(4) <= CNStageIntLLROutputS0xD(261)(1);
  VNStageIntLLRInputS0xD(146)(3) <= CNStageIntLLROutputS0xD(261)(2);
  VNStageIntLLRInputS0xD(218)(4) <= CNStageIntLLROutputS0xD(261)(3);
  VNStageIntLLRInputS0xD(310)(3) <= CNStageIntLLROutputS0xD(261)(4);
  VNStageIntLLRInputS0xD(363)(3) <= CNStageIntLLROutputS0xD(261)(5);
  VNStageIntLLRInputS0xD(38)(4) <= CNStageIntLLROutputS0xD(262)(0);
  VNStageIntLLRInputS0xD(81)(3) <= CNStageIntLLROutputS0xD(262)(1);
  VNStageIntLLRInputS0xD(153)(4) <= CNStageIntLLROutputS0xD(262)(2);
  VNStageIntLLRInputS0xD(245)(4) <= CNStageIntLLROutputS0xD(262)(3);
  VNStageIntLLRInputS0xD(298)(4) <= CNStageIntLLROutputS0xD(262)(4);
  VNStageIntLLRInputS0xD(369)(3) <= CNStageIntLLROutputS0xD(262)(5);
  VNStageIntLLRInputS0xD(37)(4) <= CNStageIntLLROutputS0xD(263)(0);
  VNStageIntLLRInputS0xD(88)(4) <= CNStageIntLLROutputS0xD(263)(1);
  VNStageIntLLRInputS0xD(180)(2) <= CNStageIntLLROutputS0xD(263)(2);
  VNStageIntLLRInputS0xD(233)(3) <= CNStageIntLLROutputS0xD(263)(3);
  VNStageIntLLRInputS0xD(304)(4) <= CNStageIntLLROutputS0xD(263)(4);
  VNStageIntLLRInputS0xD(364)(4) <= CNStageIntLLROutputS0xD(263)(5);
  VNStageIntLLRInputS0xD(36)(3) <= CNStageIntLLROutputS0xD(264)(0);
  VNStageIntLLRInputS0xD(115)(4) <= CNStageIntLLROutputS0xD(264)(1);
  VNStageIntLLRInputS0xD(168)(3) <= CNStageIntLLROutputS0xD(264)(2);
  VNStageIntLLRInputS0xD(239)(4) <= CNStageIntLLROutputS0xD(264)(3);
  VNStageIntLLRInputS0xD(299)(3) <= CNStageIntLLROutputS0xD(264)(4);
  VNStageIntLLRInputS0xD(374)(4) <= CNStageIntLLROutputS0xD(264)(5);
  VNStageIntLLRInputS0xD(35)(4) <= CNStageIntLLROutputS0xD(265)(0);
  VNStageIntLLRInputS0xD(103)(4) <= CNStageIntLLROutputS0xD(265)(1);
  VNStageIntLLRInputS0xD(174)(3) <= CNStageIntLLROutputS0xD(265)(2);
  VNStageIntLLRInputS0xD(234)(4) <= CNStageIntLLROutputS0xD(265)(3);
  VNStageIntLLRInputS0xD(309)(4) <= CNStageIntLLROutputS0xD(265)(4);
  VNStageIntLLRInputS0xD(333)(3) <= CNStageIntLLROutputS0xD(265)(5);
  VNStageIntLLRInputS0xD(34)(4) <= CNStageIntLLROutputS0xD(266)(0);
  VNStageIntLLRInputS0xD(109)(4) <= CNStageIntLLROutputS0xD(266)(1);
  VNStageIntLLRInputS0xD(169)(4) <= CNStageIntLLROutputS0xD(266)(2);
  VNStageIntLLRInputS0xD(244)(1) <= CNStageIntLLROutputS0xD(266)(3);
  VNStageIntLLRInputS0xD(268)(4) <= CNStageIntLLROutputS0xD(266)(4);
  VNStageIntLLRInputS0xD(351)(3) <= CNStageIntLLROutputS0xD(266)(5);
  VNStageIntLLRInputS0xD(33)(4) <= CNStageIntLLROutputS0xD(267)(0);
  VNStageIntLLRInputS0xD(104)(4) <= CNStageIntLLROutputS0xD(267)(1);
  VNStageIntLLRInputS0xD(179)(4) <= CNStageIntLLROutputS0xD(267)(2);
  VNStageIntLLRInputS0xD(203)(4) <= CNStageIntLLROutputS0xD(267)(3);
  VNStageIntLLRInputS0xD(286)(4) <= CNStageIntLLROutputS0xD(267)(4);
  VNStageIntLLRInputS0xD(336)(3) <= CNStageIntLLROutputS0xD(267)(5);
  VNStageIntLLRInputS0xD(32)(3) <= CNStageIntLLROutputS0xD(268)(0);
  VNStageIntLLRInputS0xD(114)(4) <= CNStageIntLLROutputS0xD(268)(1);
  VNStageIntLLRInputS0xD(138)(4) <= CNStageIntLLROutputS0xD(268)(2);
  VNStageIntLLRInputS0xD(221)(4) <= CNStageIntLLROutputS0xD(268)(3);
  VNStageIntLLRInputS0xD(271)(3) <= CNStageIntLLROutputS0xD(268)(4);
  VNStageIntLLRInputS0xD(323)(3) <= CNStageIntLLROutputS0xD(268)(5);
  VNStageIntLLRInputS0xD(30)(4) <= CNStageIntLLROutputS0xD(269)(0);
  VNStageIntLLRInputS0xD(91)(4) <= CNStageIntLLROutputS0xD(269)(1);
  VNStageIntLLRInputS0xD(141)(2) <= CNStageIntLLROutputS0xD(269)(2);
  VNStageIntLLRInputS0xD(193)(3) <= CNStageIntLLROutputS0xD(269)(3);
  VNStageIntLLRInputS0xD(289)(4) <= CNStageIntLLROutputS0xD(269)(4);
  VNStageIntLLRInputS0xD(366)(4) <= CNStageIntLLROutputS0xD(269)(5);
  VNStageIntLLRInputS0xD(29)(3) <= CNStageIntLLROutputS0xD(270)(0);
  VNStageIntLLRInputS0xD(76)(4) <= CNStageIntLLROutputS0xD(270)(1);
  VNStageIntLLRInputS0xD(191)(4) <= CNStageIntLLROutputS0xD(270)(2);
  VNStageIntLLRInputS0xD(224)(4) <= CNStageIntLLROutputS0xD(270)(3);
  VNStageIntLLRInputS0xD(301)(4) <= CNStageIntLLROutputS0xD(270)(4);
  VNStageIntLLRInputS0xD(380)(3) <= CNStageIntLLROutputS0xD(270)(5);
  VNStageIntLLRInputS0xD(28)(4) <= CNStageIntLLROutputS0xD(271)(0);
  VNStageIntLLRInputS0xD(126)(3) <= CNStageIntLLROutputS0xD(271)(1);
  VNStageIntLLRInputS0xD(159)(3) <= CNStageIntLLROutputS0xD(271)(2);
  VNStageIntLLRInputS0xD(236)(4) <= CNStageIntLLROutputS0xD(271)(3);
  VNStageIntLLRInputS0xD(315)(3) <= CNStageIntLLROutputS0xD(271)(4);
  VNStageIntLLRInputS0xD(361)(4) <= CNStageIntLLROutputS0xD(271)(5);
  VNStageIntLLRInputS0xD(26)(4) <= CNStageIntLLROutputS0xD(272)(0);
  VNStageIntLLRInputS0xD(106)(3) <= CNStageIntLLROutputS0xD(272)(1);
  VNStageIntLLRInputS0xD(185)(1) <= CNStageIntLLROutputS0xD(272)(2);
  VNStageIntLLRInputS0xD(231)(3) <= CNStageIntLLROutputS0xD(272)(3);
  VNStageIntLLRInputS0xD(273)(3) <= CNStageIntLLROutputS0xD(272)(4);
  VNStageIntLLRInputS0xD(327)(4) <= CNStageIntLLROutputS0xD(272)(5);
  VNStageIntLLRInputS0xD(24)(4) <= CNStageIntLLROutputS0xD(273)(0);
  VNStageIntLLRInputS0xD(101)(4) <= CNStageIntLLROutputS0xD(273)(1);
  VNStageIntLLRInputS0xD(143)(4) <= CNStageIntLLROutputS0xD(273)(2);
  VNStageIntLLRInputS0xD(197)(4) <= CNStageIntLLROutputS0xD(273)(3);
  VNStageIntLLRInputS0xD(266)(3) <= CNStageIntLLROutputS0xD(273)(4);
  VNStageIntLLRInputS0xD(324)(4) <= CNStageIntLLROutputS0xD(273)(5);
  VNStageIntLLRInputS0xD(23)(4) <= CNStageIntLLROutputS0xD(274)(0);
  VNStageIntLLRInputS0xD(78)(4) <= CNStageIntLLROutputS0xD(274)(1);
  VNStageIntLLRInputS0xD(132)(3) <= CNStageIntLLROutputS0xD(274)(2);
  VNStageIntLLRInputS0xD(201)(4) <= CNStageIntLLROutputS0xD(274)(3);
  VNStageIntLLRInputS0xD(259)(2) <= CNStageIntLLROutputS0xD(274)(4);
  VNStageIntLLRInputS0xD(335)(4) <= CNStageIntLLROutputS0xD(274)(5);
  VNStageIntLLRInputS0xD(22)(4) <= CNStageIntLLROutputS0xD(275)(0);
  VNStageIntLLRInputS0xD(67)(1) <= CNStageIntLLROutputS0xD(275)(1);
  VNStageIntLLRInputS0xD(136)(4) <= CNStageIntLLROutputS0xD(275)(2);
  VNStageIntLLRInputS0xD(194)(4) <= CNStageIntLLROutputS0xD(275)(3);
  VNStageIntLLRInputS0xD(270)(4) <= CNStageIntLLROutputS0xD(275)(4);
  VNStageIntLLRInputS0xD(370)(3) <= CNStageIntLLROutputS0xD(275)(5);
  VNStageIntLLRInputS0xD(21)(4) <= CNStageIntLLROutputS0xD(276)(0);
  VNStageIntLLRInputS0xD(71)(3) <= CNStageIntLLROutputS0xD(276)(1);
  VNStageIntLLRInputS0xD(129)(4) <= CNStageIntLLROutputS0xD(276)(2);
  VNStageIntLLRInputS0xD(205)(1) <= CNStageIntLLROutputS0xD(276)(3);
  VNStageIntLLRInputS0xD(305)(4) <= CNStageIntLLROutputS0xD(276)(4);
  VNStageIntLLRInputS0xD(362)(4) <= CNStageIntLLROutputS0xD(276)(5);
  VNStageIntLLRInputS0xD(20)(2) <= CNStageIntLLROutputS0xD(277)(0);
  VNStageIntLLRInputS0xD(127)(4) <= CNStageIntLLROutputS0xD(277)(1);
  VNStageIntLLRInputS0xD(140)(4) <= CNStageIntLLROutputS0xD(277)(2);
  VNStageIntLLRInputS0xD(240)(4) <= CNStageIntLLROutputS0xD(277)(3);
  VNStageIntLLRInputS0xD(297)(4) <= CNStageIntLLROutputS0xD(277)(4);
  VNStageIntLLRInputS0xD(379)(2) <= CNStageIntLLROutputS0xD(277)(5);
  VNStageIntLLRInputS0xD(19)(3) <= CNStageIntLLROutputS0xD(278)(0);
  VNStageIntLLRInputS0xD(75)(4) <= CNStageIntLLROutputS0xD(278)(1);
  VNStageIntLLRInputS0xD(175)(4) <= CNStageIntLLROutputS0xD(278)(2);
  VNStageIntLLRInputS0xD(232)(3) <= CNStageIntLLROutputS0xD(278)(3);
  VNStageIntLLRInputS0xD(314)(1) <= CNStageIntLLROutputS0xD(278)(4);
  VNStageIntLLRInputS0xD(376)(3) <= CNStageIntLLROutputS0xD(278)(5);
  VNStageIntLLRInputS0xD(0)(4) <= CNStageIntLLROutputS0xD(279)(0);
  VNStageIntLLRInputS0xD(123)(3) <= CNStageIntLLROutputS0xD(279)(1);
  VNStageIntLLRInputS0xD(188)(2) <= CNStageIntLLROutputS0xD(279)(2);
  VNStageIntLLRInputS0xD(253)(3) <= CNStageIntLLROutputS0xD(279)(3);
  VNStageIntLLRInputS0xD(318)(2) <= CNStageIntLLROutputS0xD(279)(4);
  VNStageIntLLRInputS0xD(383)(4) <= CNStageIntLLROutputS0xD(279)(5);
  VNStageIntLLRInputS0xD(35)(5) <= CNStageIntLLROutputS0xD(280)(0);
  VNStageIntLLRInputS0xD(91)(5) <= CNStageIntLLROutputS0xD(280)(1);
  VNStageIntLLRInputS0xD(191)(5) <= CNStageIntLLROutputS0xD(280)(2);
  VNStageIntLLRInputS0xD(248)(5) <= CNStageIntLLROutputS0xD(280)(3);
  VNStageIntLLRInputS0xD(267)(5) <= CNStageIntLLROutputS0xD(280)(4);
  VNStageIntLLRInputS0xD(329)(5) <= CNStageIntLLROutputS0xD(280)(5);
  VNStageIntLLRInputS0xD(34)(5) <= CNStageIntLLROutputS0xD(281)(0);
  VNStageIntLLRInputS0xD(126)(4) <= CNStageIntLLROutputS0xD(281)(1);
  VNStageIntLLRInputS0xD(183)(3) <= CNStageIntLLROutputS0xD(281)(2);
  VNStageIntLLRInputS0xD(202)(4) <= CNStageIntLLROutputS0xD(281)(3);
  VNStageIntLLRInputS0xD(264)(5) <= CNStageIntLLROutputS0xD(281)(4);
  VNStageIntLLRInputS0xD(363)(4) <= CNStageIntLLROutputS0xD(281)(5);
  VNStageIntLLRInputS0xD(33)(5) <= CNStageIntLLROutputS0xD(282)(0);
  VNStageIntLLRInputS0xD(118)(4) <= CNStageIntLLROutputS0xD(282)(1);
  VNStageIntLLRInputS0xD(137)(5) <= CNStageIntLLROutputS0xD(282)(2);
  VNStageIntLLRInputS0xD(199)(5) <= CNStageIntLLROutputS0xD(282)(3);
  VNStageIntLLRInputS0xD(298)(5) <= CNStageIntLLROutputS0xD(282)(4);
  VNStageIntLLRInputS0xD(383)(5) <= CNStageIntLLROutputS0xD(282)(5);
  VNStageIntLLRInputS0xD(31)(3) <= CNStageIntLLROutputS0xD(283)(0);
  VNStageIntLLRInputS0xD(69)(5) <= CNStageIntLLROutputS0xD(283)(1);
  VNStageIntLLRInputS0xD(168)(4) <= CNStageIntLLROutputS0xD(283)(2);
  VNStageIntLLRInputS0xD(253)(4) <= CNStageIntLLROutputS0xD(283)(3);
  VNStageIntLLRInputS0xD(304)(5) <= CNStageIntLLROutputS0xD(283)(4);
  VNStageIntLLRInputS0xD(359)(5) <= CNStageIntLLROutputS0xD(283)(5);
  VNStageIntLLRInputS0xD(30)(5) <= CNStageIntLLROutputS0xD(284)(0);
  VNStageIntLLRInputS0xD(103)(5) <= CNStageIntLLROutputS0xD(284)(1);
  VNStageIntLLRInputS0xD(188)(3) <= CNStageIntLLROutputS0xD(284)(2);
  VNStageIntLLRInputS0xD(239)(5) <= CNStageIntLLROutputS0xD(284)(3);
  VNStageIntLLRInputS0xD(294)(5) <= CNStageIntLLROutputS0xD(284)(4);
  VNStageIntLLRInputS0xD(325)(5) <= CNStageIntLLROutputS0xD(284)(5);
  VNStageIntLLRInputS0xD(27)(4) <= CNStageIntLLROutputS0xD(285)(0);
  VNStageIntLLRInputS0xD(99)(5) <= CNStageIntLLROutputS0xD(285)(1);
  VNStageIntLLRInputS0xD(130)(5) <= CNStageIntLLROutputS0xD(285)(2);
  VNStageIntLLRInputS0xD(241)(4) <= CNStageIntLLROutputS0xD(285)(3);
  VNStageIntLLRInputS0xD(273)(4) <= CNStageIntLLROutputS0xD(285)(4);
  VNStageIntLLRInputS0xD(361)(5) <= CNStageIntLLROutputS0xD(285)(5);
  VNStageIntLLRInputS0xD(26)(5) <= CNStageIntLLROutputS0xD(286)(0);
  VNStageIntLLRInputS0xD(65)(4) <= CNStageIntLLROutputS0xD(286)(1);
  VNStageIntLLRInputS0xD(176)(5) <= CNStageIntLLROutputS0xD(286)(2);
  VNStageIntLLRInputS0xD(208)(4) <= CNStageIntLLROutputS0xD(286)(3);
  VNStageIntLLRInputS0xD(296)(4) <= CNStageIntLLROutputS0xD(286)(4);
  VNStageIntLLRInputS0xD(334)(3) <= CNStageIntLLROutputS0xD(286)(5);
  VNStageIntLLRInputS0xD(25)(4) <= CNStageIntLLROutputS0xD(287)(0);
  VNStageIntLLRInputS0xD(111)(5) <= CNStageIntLLROutputS0xD(287)(1);
  VNStageIntLLRInputS0xD(143)(5) <= CNStageIntLLROutputS0xD(287)(2);
  VNStageIntLLRInputS0xD(231)(4) <= CNStageIntLLROutputS0xD(287)(3);
  VNStageIntLLRInputS0xD(269)(4) <= CNStageIntLLROutputS0xD(287)(4);
  VNStageIntLLRInputS0xD(381)(4) <= CNStageIntLLROutputS0xD(287)(5);
  VNStageIntLLRInputS0xD(24)(5) <= CNStageIntLLROutputS0xD(288)(0);
  VNStageIntLLRInputS0xD(78)(5) <= CNStageIntLLROutputS0xD(288)(1);
  VNStageIntLLRInputS0xD(166)(4) <= CNStageIntLLROutputS0xD(288)(2);
  VNStageIntLLRInputS0xD(204)(5) <= CNStageIntLLROutputS0xD(288)(3);
  VNStageIntLLRInputS0xD(316)(3) <= CNStageIntLLROutputS0xD(288)(4);
  VNStageIntLLRInputS0xD(321)(5) <= CNStageIntLLROutputS0xD(288)(5);
  VNStageIntLLRInputS0xD(23)(5) <= CNStageIntLLROutputS0xD(289)(0);
  VNStageIntLLRInputS0xD(101)(5) <= CNStageIntLLROutputS0xD(289)(1);
  VNStageIntLLRInputS0xD(139)(5) <= CNStageIntLLROutputS0xD(289)(2);
  VNStageIntLLRInputS0xD(251)(3) <= CNStageIntLLROutputS0xD(289)(3);
  VNStageIntLLRInputS0xD(319)(5) <= CNStageIntLLROutputS0xD(289)(4);
  VNStageIntLLRInputS0xD(362)(5) <= CNStageIntLLROutputS0xD(289)(5);
  VNStageIntLLRInputS0xD(22)(5) <= CNStageIntLLROutputS0xD(290)(0);
  VNStageIntLLRInputS0xD(74)(4) <= CNStageIntLLROutputS0xD(290)(1);
  VNStageIntLLRInputS0xD(186)(4) <= CNStageIntLLROutputS0xD(290)(2);
  VNStageIntLLRInputS0xD(254)(3) <= CNStageIntLLROutputS0xD(290)(3);
  VNStageIntLLRInputS0xD(297)(5) <= CNStageIntLLROutputS0xD(290)(4);
  VNStageIntLLRInputS0xD(337)(5) <= CNStageIntLLROutputS0xD(290)(5);
  VNStageIntLLRInputS0xD(21)(5) <= CNStageIntLLROutputS0xD(291)(0);
  VNStageIntLLRInputS0xD(121)(4) <= CNStageIntLLROutputS0xD(291)(1);
  VNStageIntLLRInputS0xD(189)(4) <= CNStageIntLLROutputS0xD(291)(2);
  VNStageIntLLRInputS0xD(232)(4) <= CNStageIntLLROutputS0xD(291)(3);
  VNStageIntLLRInputS0xD(272)(5) <= CNStageIntLLROutputS0xD(291)(4);
  VNStageIntLLRInputS0xD(335)(5) <= CNStageIntLLROutputS0xD(291)(5);
  VNStageIntLLRInputS0xD(20)(3) <= CNStageIntLLROutputS0xD(292)(0);
  VNStageIntLLRInputS0xD(124)(3) <= CNStageIntLLROutputS0xD(292)(1);
  VNStageIntLLRInputS0xD(167)(5) <= CNStageIntLLROutputS0xD(292)(2);
  VNStageIntLLRInputS0xD(207)(4) <= CNStageIntLLROutputS0xD(292)(3);
  VNStageIntLLRInputS0xD(270)(5) <= CNStageIntLLROutputS0xD(292)(4);
  VNStageIntLLRInputS0xD(360)(5) <= CNStageIntLLROutputS0xD(292)(5);
  VNStageIntLLRInputS0xD(18)(5) <= CNStageIntLLROutputS0xD(293)(0);
  VNStageIntLLRInputS0xD(77)(3) <= CNStageIntLLROutputS0xD(293)(1);
  VNStageIntLLRInputS0xD(140)(5) <= CNStageIntLLROutputS0xD(293)(2);
  VNStageIntLLRInputS0xD(230)(4) <= CNStageIntLLROutputS0xD(293)(3);
  VNStageIntLLRInputS0xD(303)(5) <= CNStageIntLLROutputS0xD(293)(4);
  VNStageIntLLRInputS0xD(348)(5) <= CNStageIntLLROutputS0xD(293)(5);
  VNStageIntLLRInputS0xD(17)(5) <= CNStageIntLLROutputS0xD(294)(0);
  VNStageIntLLRInputS0xD(75)(5) <= CNStageIntLLROutputS0xD(294)(1);
  VNStageIntLLRInputS0xD(165)(4) <= CNStageIntLLROutputS0xD(294)(2);
  VNStageIntLLRInputS0xD(238)(5) <= CNStageIntLLROutputS0xD(294)(3);
  VNStageIntLLRInputS0xD(283)(5) <= CNStageIntLLROutputS0xD(294)(4);
  VNStageIntLLRInputS0xD(342)(4) <= CNStageIntLLROutputS0xD(294)(5);
  VNStageIntLLRInputS0xD(16)(4) <= CNStageIntLLROutputS0xD(295)(0);
  VNStageIntLLRInputS0xD(100)(5) <= CNStageIntLLROutputS0xD(295)(1);
  VNStageIntLLRInputS0xD(173)(5) <= CNStageIntLLROutputS0xD(295)(2);
  VNStageIntLLRInputS0xD(218)(5) <= CNStageIntLLROutputS0xD(295)(3);
  VNStageIntLLRInputS0xD(277)(5) <= CNStageIntLLROutputS0xD(295)(4);
  VNStageIntLLRInputS0xD(320)(3) <= CNStageIntLLROutputS0xD(295)(5);
  VNStageIntLLRInputS0xD(15)(5) <= CNStageIntLLROutputS0xD(296)(0);
  VNStageIntLLRInputS0xD(108)(5) <= CNStageIntLLROutputS0xD(296)(1);
  VNStageIntLLRInputS0xD(153)(5) <= CNStageIntLLROutputS0xD(296)(2);
  VNStageIntLLRInputS0xD(212)(4) <= CNStageIntLLROutputS0xD(296)(3);
  VNStageIntLLRInputS0xD(256)(4) <= CNStageIntLLROutputS0xD(296)(4);
  VNStageIntLLRInputS0xD(341)(5) <= CNStageIntLLROutputS0xD(296)(5);
  VNStageIntLLRInputS0xD(14)(5) <= CNStageIntLLROutputS0xD(297)(0);
  VNStageIntLLRInputS0xD(88)(5) <= CNStageIntLLROutputS0xD(297)(1);
  VNStageIntLLRInputS0xD(147)(5) <= CNStageIntLLROutputS0xD(297)(2);
  VNStageIntLLRInputS0xD(192)(5) <= CNStageIntLLROutputS0xD(297)(3);
  VNStageIntLLRInputS0xD(276)(5) <= CNStageIntLLROutputS0xD(297)(4);
  VNStageIntLLRInputS0xD(346)(5) <= CNStageIntLLROutputS0xD(297)(5);
  VNStageIntLLRInputS0xD(13)(4) <= CNStageIntLLROutputS0xD(298)(0);
  VNStageIntLLRInputS0xD(82)(5) <= CNStageIntLLROutputS0xD(298)(1);
  VNStageIntLLRInputS0xD(128)(5) <= CNStageIntLLROutputS0xD(298)(2);
  VNStageIntLLRInputS0xD(211)(5) <= CNStageIntLLROutputS0xD(298)(3);
  VNStageIntLLRInputS0xD(281)(5) <= CNStageIntLLROutputS0xD(298)(4);
  VNStageIntLLRInputS0xD(365)(5) <= CNStageIntLLROutputS0xD(298)(5);
  VNStageIntLLRInputS0xD(12)(5) <= CNStageIntLLROutputS0xD(299)(0);
  VNStageIntLLRInputS0xD(64)(4) <= CNStageIntLLROutputS0xD(299)(1);
  VNStageIntLLRInputS0xD(146)(4) <= CNStageIntLLROutputS0xD(299)(2);
  VNStageIntLLRInputS0xD(216)(5) <= CNStageIntLLROutputS0xD(299)(3);
  VNStageIntLLRInputS0xD(300)(4) <= CNStageIntLLROutputS0xD(299)(4);
  VNStageIntLLRInputS0xD(356)(4) <= CNStageIntLLROutputS0xD(299)(5);
  VNStageIntLLRInputS0xD(9)(5) <= CNStageIntLLROutputS0xD(300)(0);
  VNStageIntLLRInputS0xD(105)(4) <= CNStageIntLLROutputS0xD(300)(1);
  VNStageIntLLRInputS0xD(161)(5) <= CNStageIntLLROutputS0xD(300)(2);
  VNStageIntLLRInputS0xD(200)(5) <= CNStageIntLLROutputS0xD(300)(3);
  VNStageIntLLRInputS0xD(266)(4) <= CNStageIntLLROutputS0xD(300)(4);
  VNStageIntLLRInputS0xD(355)(5) <= CNStageIntLLROutputS0xD(300)(5);
  VNStageIntLLRInputS0xD(7)(5) <= CNStageIntLLROutputS0xD(301)(0);
  VNStageIntLLRInputS0xD(70)(5) <= CNStageIntLLROutputS0xD(301)(1);
  VNStageIntLLRInputS0xD(136)(5) <= CNStageIntLLROutputS0xD(301)(2);
  VNStageIntLLRInputS0xD(225)(5) <= CNStageIntLLROutputS0xD(301)(3);
  VNStageIntLLRInputS0xD(311)(4) <= CNStageIntLLROutputS0xD(301)(4);
  VNStageIntLLRInputS0xD(372)(4) <= CNStageIntLLROutputS0xD(301)(5);
  VNStageIntLLRInputS0xD(6)(5) <= CNStageIntLLROutputS0xD(302)(0);
  VNStageIntLLRInputS0xD(71)(4) <= CNStageIntLLROutputS0xD(302)(1);
  VNStageIntLLRInputS0xD(160)(5) <= CNStageIntLLROutputS0xD(302)(2);
  VNStageIntLLRInputS0xD(246)(5) <= CNStageIntLLROutputS0xD(302)(3);
  VNStageIntLLRInputS0xD(307)(5) <= CNStageIntLLROutputS0xD(302)(4);
  VNStageIntLLRInputS0xD(324)(5) <= CNStageIntLLROutputS0xD(302)(5);
  VNStageIntLLRInputS0xD(5)(5) <= CNStageIntLLROutputS0xD(303)(0);
  VNStageIntLLRInputS0xD(95)(5) <= CNStageIntLLROutputS0xD(303)(1);
  VNStageIntLLRInputS0xD(181)(5) <= CNStageIntLLROutputS0xD(303)(2);
  VNStageIntLLRInputS0xD(242)(5) <= CNStageIntLLROutputS0xD(303)(3);
  VNStageIntLLRInputS0xD(259)(3) <= CNStageIntLLROutputS0xD(303)(4);
  VNStageIntLLRInputS0xD(350)(5) <= CNStageIntLLROutputS0xD(303)(5);
  VNStageIntLLRInputS0xD(4)(4) <= CNStageIntLLROutputS0xD(304)(0);
  VNStageIntLLRInputS0xD(116)(4) <= CNStageIntLLROutputS0xD(304)(1);
  VNStageIntLLRInputS0xD(177)(5) <= CNStageIntLLROutputS0xD(304)(2);
  VNStageIntLLRInputS0xD(194)(5) <= CNStageIntLLROutputS0xD(304)(3);
  VNStageIntLLRInputS0xD(285)(5) <= CNStageIntLLROutputS0xD(304)(4);
  VNStageIntLLRInputS0xD(326)(4) <= CNStageIntLLROutputS0xD(304)(5);
  VNStageIntLLRInputS0xD(3)(4) <= CNStageIntLLROutputS0xD(305)(0);
  VNStageIntLLRInputS0xD(112)(5) <= CNStageIntLLROutputS0xD(305)(1);
  VNStageIntLLRInputS0xD(129)(5) <= CNStageIntLLROutputS0xD(305)(2);
  VNStageIntLLRInputS0xD(220)(5) <= CNStageIntLLROutputS0xD(305)(3);
  VNStageIntLLRInputS0xD(261)(4) <= CNStageIntLLROutputS0xD(305)(4);
  VNStageIntLLRInputS0xD(358)(4) <= CNStageIntLLROutputS0xD(305)(5);
  VNStageIntLLRInputS0xD(2)(5) <= CNStageIntLLROutputS0xD(306)(0);
  VNStageIntLLRInputS0xD(127)(5) <= CNStageIntLLROutputS0xD(306)(1);
  VNStageIntLLRInputS0xD(155)(5) <= CNStageIntLLROutputS0xD(306)(2);
  VNStageIntLLRInputS0xD(196)(5) <= CNStageIntLLROutputS0xD(306)(3);
  VNStageIntLLRInputS0xD(293)(4) <= CNStageIntLLROutputS0xD(306)(4);
  VNStageIntLLRInputS0xD(374)(5) <= CNStageIntLLROutputS0xD(306)(5);
  VNStageIntLLRInputS0xD(1)(4) <= CNStageIntLLROutputS0xD(307)(0);
  VNStageIntLLRInputS0xD(90)(5) <= CNStageIntLLROutputS0xD(307)(1);
  VNStageIntLLRInputS0xD(131)(4) <= CNStageIntLLROutputS0xD(307)(2);
  VNStageIntLLRInputS0xD(228)(5) <= CNStageIntLLROutputS0xD(307)(3);
  VNStageIntLLRInputS0xD(309)(5) <= CNStageIntLLROutputS0xD(307)(4);
  VNStageIntLLRInputS0xD(344)(5) <= CNStageIntLLROutputS0xD(307)(5);
  VNStageIntLLRInputS0xD(62)(4) <= CNStageIntLLROutputS0xD(308)(0);
  VNStageIntLLRInputS0xD(98)(4) <= CNStageIntLLROutputS0xD(308)(1);
  VNStageIntLLRInputS0xD(179)(5) <= CNStageIntLLROutputS0xD(308)(2);
  VNStageIntLLRInputS0xD(214)(5) <= CNStageIntLLROutputS0xD(308)(3);
  VNStageIntLLRInputS0xD(288)(5) <= CNStageIntLLROutputS0xD(308)(4);
  VNStageIntLLRInputS0xD(366)(5) <= CNStageIntLLROutputS0xD(308)(5);
  VNStageIntLLRInputS0xD(61)(4) <= CNStageIntLLROutputS0xD(309)(0);
  VNStageIntLLRInputS0xD(114)(5) <= CNStageIntLLROutputS0xD(309)(1);
  VNStageIntLLRInputS0xD(149)(5) <= CNStageIntLLROutputS0xD(309)(2);
  VNStageIntLLRInputS0xD(223)(5) <= CNStageIntLLROutputS0xD(309)(3);
  VNStageIntLLRInputS0xD(301)(5) <= CNStageIntLLROutputS0xD(309)(4);
  VNStageIntLLRInputS0xD(345)(4) <= CNStageIntLLROutputS0xD(309)(5);
  VNStageIntLLRInputS0xD(60)(4) <= CNStageIntLLROutputS0xD(310)(0);
  VNStageIntLLRInputS0xD(84)(4) <= CNStageIntLLROutputS0xD(310)(1);
  VNStageIntLLRInputS0xD(158)(5) <= CNStageIntLLROutputS0xD(310)(2);
  VNStageIntLLRInputS0xD(236)(5) <= CNStageIntLLROutputS0xD(310)(3);
  VNStageIntLLRInputS0xD(280)(5) <= CNStageIntLLROutputS0xD(310)(4);
  VNStageIntLLRInputS0xD(373)(3) <= CNStageIntLLROutputS0xD(310)(5);
  VNStageIntLLRInputS0xD(59)(3) <= CNStageIntLLROutputS0xD(311)(0);
  VNStageIntLLRInputS0xD(93)(5) <= CNStageIntLLROutputS0xD(311)(1);
  VNStageIntLLRInputS0xD(171)(3) <= CNStageIntLLROutputS0xD(311)(2);
  VNStageIntLLRInputS0xD(215)(5) <= CNStageIntLLROutputS0xD(311)(3);
  VNStageIntLLRInputS0xD(308)(3) <= CNStageIntLLROutputS0xD(311)(4);
  VNStageIntLLRInputS0xD(375)(4) <= CNStageIntLLROutputS0xD(311)(5);
  VNStageIntLLRInputS0xD(58)(3) <= CNStageIntLLROutputS0xD(312)(0);
  VNStageIntLLRInputS0xD(106)(4) <= CNStageIntLLROutputS0xD(312)(1);
  VNStageIntLLRInputS0xD(150)(4) <= CNStageIntLLROutputS0xD(312)(2);
  VNStageIntLLRInputS0xD(243)(5) <= CNStageIntLLROutputS0xD(312)(3);
  VNStageIntLLRInputS0xD(310)(4) <= CNStageIntLLROutputS0xD(312)(4);
  VNStageIntLLRInputS0xD(357)(5) <= CNStageIntLLROutputS0xD(312)(5);
  VNStageIntLLRInputS0xD(57)(4) <= CNStageIntLLROutputS0xD(313)(0);
  VNStageIntLLRInputS0xD(85)(4) <= CNStageIntLLROutputS0xD(313)(1);
  VNStageIntLLRInputS0xD(178)(4) <= CNStageIntLLROutputS0xD(313)(2);
  VNStageIntLLRInputS0xD(245)(5) <= CNStageIntLLROutputS0xD(313)(3);
  VNStageIntLLRInputS0xD(292)(5) <= CNStageIntLLROutputS0xD(313)(4);
  VNStageIntLLRInputS0xD(364)(5) <= CNStageIntLLROutputS0xD(313)(5);
  VNStageIntLLRInputS0xD(56)(5) <= CNStageIntLLROutputS0xD(314)(0);
  VNStageIntLLRInputS0xD(113)(5) <= CNStageIntLLROutputS0xD(314)(1);
  VNStageIntLLRInputS0xD(180)(3) <= CNStageIntLLROutputS0xD(314)(2);
  VNStageIntLLRInputS0xD(227)(5) <= CNStageIntLLROutputS0xD(314)(3);
  VNStageIntLLRInputS0xD(299)(4) <= CNStageIntLLROutputS0xD(314)(4);
  VNStageIntLLRInputS0xD(328)(3) <= CNStageIntLLROutputS0xD(314)(5);
  VNStageIntLLRInputS0xD(55)(5) <= CNStageIntLLROutputS0xD(315)(0);
  VNStageIntLLRInputS0xD(115)(5) <= CNStageIntLLROutputS0xD(315)(1);
  VNStageIntLLRInputS0xD(162)(5) <= CNStageIntLLROutputS0xD(315)(2);
  VNStageIntLLRInputS0xD(234)(5) <= CNStageIntLLROutputS0xD(315)(3);
  VNStageIntLLRInputS0xD(263)(5) <= CNStageIntLLROutputS0xD(315)(4);
  VNStageIntLLRInputS0xD(379)(3) <= CNStageIntLLROutputS0xD(315)(5);
  VNStageIntLLRInputS0xD(54)(4) <= CNStageIntLLROutputS0xD(316)(0);
  VNStageIntLLRInputS0xD(97)(5) <= CNStageIntLLROutputS0xD(316)(1);
  VNStageIntLLRInputS0xD(169)(5) <= CNStageIntLLROutputS0xD(316)(2);
  VNStageIntLLRInputS0xD(198)(5) <= CNStageIntLLROutputS0xD(316)(3);
  VNStageIntLLRInputS0xD(314)(2) <= CNStageIntLLROutputS0xD(316)(4);
  VNStageIntLLRInputS0xD(322)(4) <= CNStageIntLLROutputS0xD(316)(5);
  VNStageIntLLRInputS0xD(53)(4) <= CNStageIntLLROutputS0xD(317)(0);
  VNStageIntLLRInputS0xD(104)(5) <= CNStageIntLLROutputS0xD(317)(1);
  VNStageIntLLRInputS0xD(133)(3) <= CNStageIntLLROutputS0xD(317)(2);
  VNStageIntLLRInputS0xD(249)(3) <= CNStageIntLLROutputS0xD(317)(3);
  VNStageIntLLRInputS0xD(257)(5) <= CNStageIntLLROutputS0xD(317)(4);
  VNStageIntLLRInputS0xD(380)(4) <= CNStageIntLLROutputS0xD(317)(5);
  VNStageIntLLRInputS0xD(52)(3) <= CNStageIntLLROutputS0xD(318)(0);
  VNStageIntLLRInputS0xD(68)(4) <= CNStageIntLLROutputS0xD(318)(1);
  VNStageIntLLRInputS0xD(184)(5) <= CNStageIntLLROutputS0xD(318)(2);
  VNStageIntLLRInputS0xD(255)(5) <= CNStageIntLLROutputS0xD(318)(3);
  VNStageIntLLRInputS0xD(315)(4) <= CNStageIntLLROutputS0xD(318)(4);
  VNStageIntLLRInputS0xD(327)(5) <= CNStageIntLLROutputS0xD(318)(5);
  VNStageIntLLRInputS0xD(51)(4) <= CNStageIntLLROutputS0xD(319)(0);
  VNStageIntLLRInputS0xD(119)(4) <= CNStageIntLLROutputS0xD(319)(1);
  VNStageIntLLRInputS0xD(190)(3) <= CNStageIntLLROutputS0xD(319)(2);
  VNStageIntLLRInputS0xD(250)(3) <= CNStageIntLLROutputS0xD(319)(3);
  VNStageIntLLRInputS0xD(262)(4) <= CNStageIntLLROutputS0xD(319)(4);
  VNStageIntLLRInputS0xD(349)(4) <= CNStageIntLLROutputS0xD(319)(5);
  VNStageIntLLRInputS0xD(50)(5) <= CNStageIntLLROutputS0xD(320)(0);
  VNStageIntLLRInputS0xD(125)(2) <= CNStageIntLLROutputS0xD(320)(1);
  VNStageIntLLRInputS0xD(185)(2) <= CNStageIntLLROutputS0xD(320)(2);
  VNStageIntLLRInputS0xD(197)(5) <= CNStageIntLLROutputS0xD(320)(3);
  VNStageIntLLRInputS0xD(284)(5) <= CNStageIntLLROutputS0xD(320)(4);
  VNStageIntLLRInputS0xD(367)(5) <= CNStageIntLLROutputS0xD(320)(5);
  VNStageIntLLRInputS0xD(49)(5) <= CNStageIntLLROutputS0xD(321)(0);
  VNStageIntLLRInputS0xD(120)(2) <= CNStageIntLLROutputS0xD(321)(1);
  VNStageIntLLRInputS0xD(132)(4) <= CNStageIntLLROutputS0xD(321)(2);
  VNStageIntLLRInputS0xD(219)(4) <= CNStageIntLLROutputS0xD(321)(3);
  VNStageIntLLRInputS0xD(302)(5) <= CNStageIntLLROutputS0xD(321)(4);
  VNStageIntLLRInputS0xD(352)(5) <= CNStageIntLLROutputS0xD(321)(5);
  VNStageIntLLRInputS0xD(48)(2) <= CNStageIntLLROutputS0xD(322)(0);
  VNStageIntLLRInputS0xD(67)(2) <= CNStageIntLLROutputS0xD(322)(1);
  VNStageIntLLRInputS0xD(154)(4) <= CNStageIntLLROutputS0xD(322)(2);
  VNStageIntLLRInputS0xD(237)(4) <= CNStageIntLLROutputS0xD(322)(3);
  VNStageIntLLRInputS0xD(287)(5) <= CNStageIntLLROutputS0xD(322)(4);
  VNStageIntLLRInputS0xD(339)(5) <= CNStageIntLLROutputS0xD(322)(5);
  VNStageIntLLRInputS0xD(46)(5) <= CNStageIntLLROutputS0xD(323)(0);
  VNStageIntLLRInputS0xD(107)(4) <= CNStageIntLLROutputS0xD(323)(1);
  VNStageIntLLRInputS0xD(157)(4) <= CNStageIntLLROutputS0xD(323)(2);
  VNStageIntLLRInputS0xD(209)(4) <= CNStageIntLLROutputS0xD(323)(3);
  VNStageIntLLRInputS0xD(305)(5) <= CNStageIntLLROutputS0xD(323)(4);
  VNStageIntLLRInputS0xD(382)(4) <= CNStageIntLLROutputS0xD(323)(5);
  VNStageIntLLRInputS0xD(45)(5) <= CNStageIntLLROutputS0xD(324)(0);
  VNStageIntLLRInputS0xD(92)(5) <= CNStageIntLLROutputS0xD(324)(1);
  VNStageIntLLRInputS0xD(144)(5) <= CNStageIntLLROutputS0xD(324)(2);
  VNStageIntLLRInputS0xD(240)(5) <= CNStageIntLLROutputS0xD(324)(3);
  VNStageIntLLRInputS0xD(317)(2) <= CNStageIntLLROutputS0xD(324)(4);
  VNStageIntLLRInputS0xD(333)(4) <= CNStageIntLLROutputS0xD(324)(5);
  VNStageIntLLRInputS0xD(44)(5) <= CNStageIntLLROutputS0xD(325)(0);
  VNStageIntLLRInputS0xD(79)(4) <= CNStageIntLLROutputS0xD(325)(1);
  VNStageIntLLRInputS0xD(175)(5) <= CNStageIntLLROutputS0xD(325)(2);
  VNStageIntLLRInputS0xD(252)(4) <= CNStageIntLLROutputS0xD(325)(3);
  VNStageIntLLRInputS0xD(268)(5) <= CNStageIntLLROutputS0xD(325)(4);
  VNStageIntLLRInputS0xD(377)(3) <= CNStageIntLLROutputS0xD(325)(5);
  VNStageIntLLRInputS0xD(43)(4) <= CNStageIntLLROutputS0xD(326)(0);
  VNStageIntLLRInputS0xD(110)(5) <= CNStageIntLLROutputS0xD(326)(1);
  VNStageIntLLRInputS0xD(187)(4) <= CNStageIntLLROutputS0xD(326)(2);
  VNStageIntLLRInputS0xD(203)(5) <= CNStageIntLLROutputS0xD(326)(3);
  VNStageIntLLRInputS0xD(312)(4) <= CNStageIntLLROutputS0xD(326)(4);
  VNStageIntLLRInputS0xD(354)(4) <= CNStageIntLLROutputS0xD(326)(5);
  VNStageIntLLRInputS0xD(42)(5) <= CNStageIntLLROutputS0xD(327)(0);
  VNStageIntLLRInputS0xD(122)(4) <= CNStageIntLLROutputS0xD(327)(1);
  VNStageIntLLRInputS0xD(138)(5) <= CNStageIntLLROutputS0xD(327)(2);
  VNStageIntLLRInputS0xD(247)(5) <= CNStageIntLLROutputS0xD(327)(3);
  VNStageIntLLRInputS0xD(289)(5) <= CNStageIntLLROutputS0xD(327)(4);
  VNStageIntLLRInputS0xD(343)(5) <= CNStageIntLLROutputS0xD(327)(5);
  VNStageIntLLRInputS0xD(41)(5) <= CNStageIntLLROutputS0xD(328)(0);
  VNStageIntLLRInputS0xD(73)(4) <= CNStageIntLLROutputS0xD(328)(1);
  VNStageIntLLRInputS0xD(182)(5) <= CNStageIntLLROutputS0xD(328)(2);
  VNStageIntLLRInputS0xD(224)(5) <= CNStageIntLLROutputS0xD(328)(3);
  VNStageIntLLRInputS0xD(278)(4) <= CNStageIntLLROutputS0xD(328)(4);
  VNStageIntLLRInputS0xD(347)(5) <= CNStageIntLLROutputS0xD(328)(5);
  VNStageIntLLRInputS0xD(39)(5) <= CNStageIntLLROutputS0xD(329)(0);
  VNStageIntLLRInputS0xD(94)(3) <= CNStageIntLLROutputS0xD(329)(1);
  VNStageIntLLRInputS0xD(148)(5) <= CNStageIntLLROutputS0xD(329)(2);
  VNStageIntLLRInputS0xD(217)(5) <= CNStageIntLLROutputS0xD(329)(3);
  VNStageIntLLRInputS0xD(275)(4) <= CNStageIntLLROutputS0xD(329)(4);
  VNStageIntLLRInputS0xD(351)(4) <= CNStageIntLLROutputS0xD(329)(5);
  VNStageIntLLRInputS0xD(38)(5) <= CNStageIntLLROutputS0xD(330)(0);
  VNStageIntLLRInputS0xD(83)(5) <= CNStageIntLLROutputS0xD(330)(1);
  VNStageIntLLRInputS0xD(152)(5) <= CNStageIntLLROutputS0xD(330)(2);
  VNStageIntLLRInputS0xD(210)(5) <= CNStageIntLLROutputS0xD(330)(3);
  VNStageIntLLRInputS0xD(286)(5) <= CNStageIntLLROutputS0xD(330)(4);
  VNStageIntLLRInputS0xD(323)(4) <= CNStageIntLLROutputS0xD(330)(5);
  VNStageIntLLRInputS0xD(37)(5) <= CNStageIntLLROutputS0xD(331)(0);
  VNStageIntLLRInputS0xD(87)(5) <= CNStageIntLLROutputS0xD(331)(1);
  VNStageIntLLRInputS0xD(145)(5) <= CNStageIntLLROutputS0xD(331)(2);
  VNStageIntLLRInputS0xD(221)(5) <= CNStageIntLLROutputS0xD(331)(3);
  VNStageIntLLRInputS0xD(258)(2) <= CNStageIntLLROutputS0xD(331)(4);
  VNStageIntLLRInputS0xD(378)(4) <= CNStageIntLLROutputS0xD(331)(5);
  VNStageIntLLRInputS0xD(0)(5) <= CNStageIntLLROutputS0xD(332)(0);
  VNStageIntLLRInputS0xD(76)(5) <= CNStageIntLLROutputS0xD(332)(1);
  VNStageIntLLRInputS0xD(141)(3) <= CNStageIntLLROutputS0xD(332)(2);
  VNStageIntLLRInputS0xD(206)(3) <= CNStageIntLLROutputS0xD(332)(3);
  VNStageIntLLRInputS0xD(271)(4) <= CNStageIntLLROutputS0xD(332)(4);
  VNStageIntLLRInputS0xD(336)(4) <= CNStageIntLLROutputS0xD(332)(5);
  VNStageIntLLRInputS0xD(28)(5) <= CNStageIntLLROutputS0xD(333)(0);
  VNStageIntLLRInputS0xD(106)(5) <= CNStageIntLLROutputS0xD(333)(1);
  VNStageIntLLRInputS0xD(144)(6) <= CNStageIntLLROutputS0xD(333)(2);
  VNStageIntLLRInputS0xD(193)(4) <= CNStageIntLLROutputS0xD(333)(3);
  VNStageIntLLRInputS0xD(261)(5) <= CNStageIntLLROutputS0xD(333)(4);
  VNStageIntLLRInputS0xD(367)(6) <= CNStageIntLLROutputS0xD(333)(5);
  VNStageIntLLRInputS0xD(26)(6) <= CNStageIntLLROutputS0xD(334)(0);
  VNStageIntLLRInputS0xD(126)(5) <= CNStageIntLLROutputS0xD(334)(1);
  VNStageIntLLRInputS0xD(131)(5) <= CNStageIntLLROutputS0xD(334)(2);
  VNStageIntLLRInputS0xD(237)(5) <= CNStageIntLLROutputS0xD(334)(3);
  VNStageIntLLRInputS0xD(277)(6) <= CNStageIntLLROutputS0xD(334)(4);
  VNStageIntLLRInputS0xD(340)(5) <= CNStageIntLLROutputS0xD(334)(5);
  VNStageIntLLRInputS0xD(24)(6) <= CNStageIntLLROutputS0xD(335)(0);
  VNStageIntLLRInputS0xD(107)(5) <= CNStageIntLLROutputS0xD(335)(1);
  VNStageIntLLRInputS0xD(147)(6) <= CNStageIntLLROutputS0xD(335)(2);
  VNStageIntLLRInputS0xD(210)(6) <= CNStageIntLLROutputS0xD(335)(3);
  VNStageIntLLRInputS0xD(300)(5) <= CNStageIntLLROutputS0xD(335)(4);
  VNStageIntLLRInputS0xD(373)(4) <= CNStageIntLLROutputS0xD(335)(5);
  VNStageIntLLRInputS0xD(23)(6) <= CNStageIntLLROutputS0xD(336)(0);
  VNStageIntLLRInputS0xD(82)(6) <= CNStageIntLLROutputS0xD(336)(1);
  VNStageIntLLRInputS0xD(145)(6) <= CNStageIntLLROutputS0xD(336)(2);
  VNStageIntLLRInputS0xD(235)(4) <= CNStageIntLLROutputS0xD(336)(3);
  VNStageIntLLRInputS0xD(308)(4) <= CNStageIntLLROutputS0xD(336)(4);
  VNStageIntLLRInputS0xD(353)(5) <= CNStageIntLLROutputS0xD(336)(5);
  VNStageIntLLRInputS0xD(22)(6) <= CNStageIntLLROutputS0xD(337)(0);
  VNStageIntLLRInputS0xD(80)(5) <= CNStageIntLLROutputS0xD(337)(1);
  VNStageIntLLRInputS0xD(170)(4) <= CNStageIntLLROutputS0xD(337)(2);
  VNStageIntLLRInputS0xD(243)(6) <= CNStageIntLLROutputS0xD(337)(3);
  VNStageIntLLRInputS0xD(288)(6) <= CNStageIntLLROutputS0xD(337)(4);
  VNStageIntLLRInputS0xD(347)(6) <= CNStageIntLLROutputS0xD(337)(5);
  VNStageIntLLRInputS0xD(21)(6) <= CNStageIntLLROutputS0xD(338)(0);
  VNStageIntLLRInputS0xD(105)(5) <= CNStageIntLLROutputS0xD(338)(1);
  VNStageIntLLRInputS0xD(178)(5) <= CNStageIntLLROutputS0xD(338)(2);
  VNStageIntLLRInputS0xD(223)(6) <= CNStageIntLLROutputS0xD(338)(3);
  VNStageIntLLRInputS0xD(282)(5) <= CNStageIntLLROutputS0xD(338)(4);
  VNStageIntLLRInputS0xD(320)(4) <= CNStageIntLLROutputS0xD(338)(5);
  VNStageIntLLRInputS0xD(20)(4) <= CNStageIntLLROutputS0xD(339)(0);
  VNStageIntLLRInputS0xD(113)(6) <= CNStageIntLLROutputS0xD(339)(1);
  VNStageIntLLRInputS0xD(158)(6) <= CNStageIntLLROutputS0xD(339)(2);
  VNStageIntLLRInputS0xD(217)(6) <= CNStageIntLLROutputS0xD(339)(3);
  VNStageIntLLRInputS0xD(256)(5) <= CNStageIntLLROutputS0xD(339)(4);
  VNStageIntLLRInputS0xD(346)(6) <= CNStageIntLLROutputS0xD(339)(5);
  VNStageIntLLRInputS0xD(19)(4) <= CNStageIntLLROutputS0xD(340)(0);
  VNStageIntLLRInputS0xD(93)(6) <= CNStageIntLLROutputS0xD(340)(1);
  VNStageIntLLRInputS0xD(152)(6) <= CNStageIntLLROutputS0xD(340)(2);
  VNStageIntLLRInputS0xD(192)(6) <= CNStageIntLLROutputS0xD(340)(3);
  VNStageIntLLRInputS0xD(281)(6) <= CNStageIntLLROutputS0xD(340)(4);
  VNStageIntLLRInputS0xD(351)(5) <= CNStageIntLLROutputS0xD(340)(5);
  VNStageIntLLRInputS0xD(18)(6) <= CNStageIntLLROutputS0xD(341)(0);
  VNStageIntLLRInputS0xD(87)(6) <= CNStageIntLLROutputS0xD(341)(1);
  VNStageIntLLRInputS0xD(128)(6) <= CNStageIntLLROutputS0xD(341)(2);
  VNStageIntLLRInputS0xD(216)(6) <= CNStageIntLLROutputS0xD(341)(3);
  VNStageIntLLRInputS0xD(286)(6) <= CNStageIntLLROutputS0xD(341)(4);
  VNStageIntLLRInputS0xD(370)(4) <= CNStageIntLLROutputS0xD(341)(5);
  VNStageIntLLRInputS0xD(17)(6) <= CNStageIntLLROutputS0xD(342)(0);
  VNStageIntLLRInputS0xD(64)(5) <= CNStageIntLLROutputS0xD(342)(1);
  VNStageIntLLRInputS0xD(151)(5) <= CNStageIntLLROutputS0xD(342)(2);
  VNStageIntLLRInputS0xD(221)(6) <= CNStageIntLLROutputS0xD(342)(3);
  VNStageIntLLRInputS0xD(305)(6) <= CNStageIntLLROutputS0xD(342)(4);
  VNStageIntLLRInputS0xD(361)(6) <= CNStageIntLLROutputS0xD(342)(5);
  VNStageIntLLRInputS0xD(16)(5) <= CNStageIntLLROutputS0xD(343)(0);
  VNStageIntLLRInputS0xD(86)(3) <= CNStageIntLLROutputS0xD(343)(1);
  VNStageIntLLRInputS0xD(156)(3) <= CNStageIntLLROutputS0xD(343)(2);
  VNStageIntLLRInputS0xD(240)(6) <= CNStageIntLLROutputS0xD(343)(3);
  VNStageIntLLRInputS0xD(296)(5) <= CNStageIntLLROutputS0xD(343)(4);
  VNStageIntLLRInputS0xD(335)(6) <= CNStageIntLLROutputS0xD(343)(5);
  VNStageIntLLRInputS0xD(15)(6) <= CNStageIntLLROutputS0xD(344)(0);
  VNStageIntLLRInputS0xD(91)(6) <= CNStageIntLLROutputS0xD(344)(1);
  VNStageIntLLRInputS0xD(175)(6) <= CNStageIntLLROutputS0xD(344)(2);
  VNStageIntLLRInputS0xD(231)(5) <= CNStageIntLLROutputS0xD(344)(3);
  VNStageIntLLRInputS0xD(270)(6) <= CNStageIntLLROutputS0xD(344)(4);
  VNStageIntLLRInputS0xD(336)(5) <= CNStageIntLLROutputS0xD(344)(5);
  VNStageIntLLRInputS0xD(14)(6) <= CNStageIntLLROutputS0xD(345)(0);
  VNStageIntLLRInputS0xD(110)(6) <= CNStageIntLLROutputS0xD(345)(1);
  VNStageIntLLRInputS0xD(166)(5) <= CNStageIntLLROutputS0xD(345)(2);
  VNStageIntLLRInputS0xD(205)(2) <= CNStageIntLLROutputS0xD(345)(3);
  VNStageIntLLRInputS0xD(271)(5) <= CNStageIntLLROutputS0xD(345)(4);
  VNStageIntLLRInputS0xD(360)(6) <= CNStageIntLLROutputS0xD(345)(5);
  VNStageIntLLRInputS0xD(13)(5) <= CNStageIntLLROutputS0xD(346)(0);
  VNStageIntLLRInputS0xD(101)(6) <= CNStageIntLLROutputS0xD(346)(1);
  VNStageIntLLRInputS0xD(140)(6) <= CNStageIntLLROutputS0xD(346)(2);
  VNStageIntLLRInputS0xD(206)(4) <= CNStageIntLLROutputS0xD(346)(3);
  VNStageIntLLRInputS0xD(295)(4) <= CNStageIntLLROutputS0xD(346)(4);
  VNStageIntLLRInputS0xD(381)(5) <= CNStageIntLLROutputS0xD(346)(5);
  VNStageIntLLRInputS0xD(12)(6) <= CNStageIntLLROutputS0xD(347)(0);
  VNStageIntLLRInputS0xD(75)(6) <= CNStageIntLLROutputS0xD(347)(1);
  VNStageIntLLRInputS0xD(141)(4) <= CNStageIntLLROutputS0xD(347)(2);
  VNStageIntLLRInputS0xD(230)(5) <= CNStageIntLLROutputS0xD(347)(3);
  VNStageIntLLRInputS0xD(316)(4) <= CNStageIntLLROutputS0xD(347)(4);
  VNStageIntLLRInputS0xD(377)(4) <= CNStageIntLLROutputS0xD(347)(5);
  VNStageIntLLRInputS0xD(11)(5) <= CNStageIntLLROutputS0xD(348)(0);
  VNStageIntLLRInputS0xD(76)(6) <= CNStageIntLLROutputS0xD(348)(1);
  VNStageIntLLRInputS0xD(165)(5) <= CNStageIntLLROutputS0xD(348)(2);
  VNStageIntLLRInputS0xD(251)(4) <= CNStageIntLLROutputS0xD(348)(3);
  VNStageIntLLRInputS0xD(312)(5) <= CNStageIntLLROutputS0xD(348)(4);
  VNStageIntLLRInputS0xD(329)(6) <= CNStageIntLLROutputS0xD(348)(5);
  VNStageIntLLRInputS0xD(10)(4) <= CNStageIntLLROutputS0xD(349)(0);
  VNStageIntLLRInputS0xD(100)(6) <= CNStageIntLLROutputS0xD(349)(1);
  VNStageIntLLRInputS0xD(186)(5) <= CNStageIntLLROutputS0xD(349)(2);
  VNStageIntLLRInputS0xD(247)(6) <= CNStageIntLLROutputS0xD(349)(3);
  VNStageIntLLRInputS0xD(264)(6) <= CNStageIntLLROutputS0xD(349)(4);
  VNStageIntLLRInputS0xD(355)(6) <= CNStageIntLLROutputS0xD(349)(5);
  VNStageIntLLRInputS0xD(9)(6) <= CNStageIntLLROutputS0xD(350)(0);
  VNStageIntLLRInputS0xD(121)(5) <= CNStageIntLLROutputS0xD(350)(1);
  VNStageIntLLRInputS0xD(182)(6) <= CNStageIntLLROutputS0xD(350)(2);
  VNStageIntLLRInputS0xD(199)(6) <= CNStageIntLLROutputS0xD(350)(3);
  VNStageIntLLRInputS0xD(290)(5) <= CNStageIntLLROutputS0xD(350)(4);
  VNStageIntLLRInputS0xD(331)(4) <= CNStageIntLLROutputS0xD(350)(5);
  VNStageIntLLRInputS0xD(7)(6) <= CNStageIntLLROutputS0xD(351)(0);
  VNStageIntLLRInputS0xD(69)(6) <= CNStageIntLLROutputS0xD(351)(1);
  VNStageIntLLRInputS0xD(160)(6) <= CNStageIntLLROutputS0xD(351)(2);
  VNStageIntLLRInputS0xD(201)(5) <= CNStageIntLLROutputS0xD(351)(3);
  VNStageIntLLRInputS0xD(298)(6) <= CNStageIntLLROutputS0xD(351)(4);
  VNStageIntLLRInputS0xD(379)(4) <= CNStageIntLLROutputS0xD(351)(5);
  VNStageIntLLRInputS0xD(6)(6) <= CNStageIntLLROutputS0xD(352)(0);
  VNStageIntLLRInputS0xD(95)(6) <= CNStageIntLLROutputS0xD(352)(1);
  VNStageIntLLRInputS0xD(136)(6) <= CNStageIntLLROutputS0xD(352)(2);
  VNStageIntLLRInputS0xD(233)(4) <= CNStageIntLLROutputS0xD(352)(3);
  VNStageIntLLRInputS0xD(314)(3) <= CNStageIntLLROutputS0xD(352)(4);
  VNStageIntLLRInputS0xD(349)(5) <= CNStageIntLLROutputS0xD(352)(5);
  VNStageIntLLRInputS0xD(5)(6) <= CNStageIntLLROutputS0xD(353)(0);
  VNStageIntLLRInputS0xD(71)(5) <= CNStageIntLLROutputS0xD(353)(1);
  VNStageIntLLRInputS0xD(168)(5) <= CNStageIntLLROutputS0xD(353)(2);
  VNStageIntLLRInputS0xD(249)(4) <= CNStageIntLLROutputS0xD(353)(3);
  VNStageIntLLRInputS0xD(284)(6) <= CNStageIntLLROutputS0xD(353)(4);
  VNStageIntLLRInputS0xD(358)(5) <= CNStageIntLLROutputS0xD(353)(5);
  VNStageIntLLRInputS0xD(4)(5) <= CNStageIntLLROutputS0xD(354)(0);
  VNStageIntLLRInputS0xD(103)(6) <= CNStageIntLLROutputS0xD(354)(1);
  VNStageIntLLRInputS0xD(184)(6) <= CNStageIntLLROutputS0xD(354)(2);
  VNStageIntLLRInputS0xD(219)(5) <= CNStageIntLLROutputS0xD(354)(3);
  VNStageIntLLRInputS0xD(293)(5) <= CNStageIntLLROutputS0xD(354)(4);
  VNStageIntLLRInputS0xD(371)(4) <= CNStageIntLLROutputS0xD(354)(5);
  VNStageIntLLRInputS0xD(2)(6) <= CNStageIntLLROutputS0xD(355)(0);
  VNStageIntLLRInputS0xD(89)(5) <= CNStageIntLLROutputS0xD(355)(1);
  VNStageIntLLRInputS0xD(163)(4) <= CNStageIntLLROutputS0xD(355)(2);
  VNStageIntLLRInputS0xD(241)(5) <= CNStageIntLLROutputS0xD(355)(3);
  VNStageIntLLRInputS0xD(285)(6) <= CNStageIntLLROutputS0xD(355)(4);
  VNStageIntLLRInputS0xD(378)(5) <= CNStageIntLLROutputS0xD(355)(5);
  VNStageIntLLRInputS0xD(1)(5) <= CNStageIntLLROutputS0xD(356)(0);
  VNStageIntLLRInputS0xD(98)(5) <= CNStageIntLLROutputS0xD(356)(1);
  VNStageIntLLRInputS0xD(176)(6) <= CNStageIntLLROutputS0xD(356)(2);
  VNStageIntLLRInputS0xD(220)(6) <= CNStageIntLLROutputS0xD(356)(3);
  VNStageIntLLRInputS0xD(313)(3) <= CNStageIntLLROutputS0xD(356)(4);
  VNStageIntLLRInputS0xD(380)(5) <= CNStageIntLLROutputS0xD(356)(5);
  VNStageIntLLRInputS0xD(63)(3) <= CNStageIntLLROutputS0xD(357)(0);
  VNStageIntLLRInputS0xD(111)(6) <= CNStageIntLLROutputS0xD(357)(1);
  VNStageIntLLRInputS0xD(155)(6) <= CNStageIntLLROutputS0xD(357)(2);
  VNStageIntLLRInputS0xD(248)(6) <= CNStageIntLLROutputS0xD(357)(3);
  VNStageIntLLRInputS0xD(315)(5) <= CNStageIntLLROutputS0xD(357)(4);
  VNStageIntLLRInputS0xD(362)(6) <= CNStageIntLLROutputS0xD(357)(5);
  VNStageIntLLRInputS0xD(62)(5) <= CNStageIntLLROutputS0xD(358)(0);
  VNStageIntLLRInputS0xD(90)(6) <= CNStageIntLLROutputS0xD(358)(1);
  VNStageIntLLRInputS0xD(183)(4) <= CNStageIntLLROutputS0xD(358)(2);
  VNStageIntLLRInputS0xD(250)(4) <= CNStageIntLLROutputS0xD(358)(3);
  VNStageIntLLRInputS0xD(297)(6) <= CNStageIntLLROutputS0xD(358)(4);
  VNStageIntLLRInputS0xD(369)(4) <= CNStageIntLLROutputS0xD(358)(5);
  VNStageIntLLRInputS0xD(61)(5) <= CNStageIntLLROutputS0xD(359)(0);
  VNStageIntLLRInputS0xD(118)(5) <= CNStageIntLLROutputS0xD(359)(1);
  VNStageIntLLRInputS0xD(185)(3) <= CNStageIntLLROutputS0xD(359)(2);
  VNStageIntLLRInputS0xD(232)(5) <= CNStageIntLLROutputS0xD(359)(3);
  VNStageIntLLRInputS0xD(304)(6) <= CNStageIntLLROutputS0xD(359)(4);
  VNStageIntLLRInputS0xD(333)(5) <= CNStageIntLLROutputS0xD(359)(5);
  VNStageIntLLRInputS0xD(60)(5) <= CNStageIntLLROutputS0xD(360)(0);
  VNStageIntLLRInputS0xD(120)(3) <= CNStageIntLLROutputS0xD(360)(1);
  VNStageIntLLRInputS0xD(167)(6) <= CNStageIntLLROutputS0xD(360)(2);
  VNStageIntLLRInputS0xD(239)(6) <= CNStageIntLLROutputS0xD(360)(3);
  VNStageIntLLRInputS0xD(268)(6) <= CNStageIntLLROutputS0xD(360)(4);
  VNStageIntLLRInputS0xD(321)(6) <= CNStageIntLLROutputS0xD(360)(5);
  VNStageIntLLRInputS0xD(59)(4) <= CNStageIntLLROutputS0xD(361)(0);
  VNStageIntLLRInputS0xD(102)(5) <= CNStageIntLLROutputS0xD(361)(1);
  VNStageIntLLRInputS0xD(174)(4) <= CNStageIntLLROutputS0xD(361)(2);
  VNStageIntLLRInputS0xD(203)(6) <= CNStageIntLLROutputS0xD(361)(3);
  VNStageIntLLRInputS0xD(319)(6) <= CNStageIntLLROutputS0xD(361)(4);
  VNStageIntLLRInputS0xD(327)(6) <= CNStageIntLLROutputS0xD(361)(5);
  VNStageIntLLRInputS0xD(58)(4) <= CNStageIntLLROutputS0xD(362)(0);
  VNStageIntLLRInputS0xD(109)(5) <= CNStageIntLLROutputS0xD(362)(1);
  VNStageIntLLRInputS0xD(138)(6) <= CNStageIntLLROutputS0xD(362)(2);
  VNStageIntLLRInputS0xD(254)(4) <= CNStageIntLLROutputS0xD(362)(3);
  VNStageIntLLRInputS0xD(262)(5) <= CNStageIntLLROutputS0xD(362)(4);
  VNStageIntLLRInputS0xD(322)(5) <= CNStageIntLLROutputS0xD(362)(5);
  VNStageIntLLRInputS0xD(57)(5) <= CNStageIntLLROutputS0xD(363)(0);
  VNStageIntLLRInputS0xD(73)(5) <= CNStageIntLLROutputS0xD(363)(1);
  VNStageIntLLRInputS0xD(189)(5) <= CNStageIntLLROutputS0xD(363)(2);
  VNStageIntLLRInputS0xD(197)(6) <= CNStageIntLLROutputS0xD(363)(3);
  VNStageIntLLRInputS0xD(257)(6) <= CNStageIntLLROutputS0xD(363)(4);
  VNStageIntLLRInputS0xD(332)(5) <= CNStageIntLLROutputS0xD(363)(5);
  VNStageIntLLRInputS0xD(56)(6) <= CNStageIntLLROutputS0xD(364)(0);
  VNStageIntLLRInputS0xD(124)(4) <= CNStageIntLLROutputS0xD(364)(1);
  VNStageIntLLRInputS0xD(132)(5) <= CNStageIntLLROutputS0xD(364)(2);
  VNStageIntLLRInputS0xD(255)(6) <= CNStageIntLLROutputS0xD(364)(3);
  VNStageIntLLRInputS0xD(267)(6) <= CNStageIntLLROutputS0xD(364)(4);
  VNStageIntLLRInputS0xD(354)(5) <= CNStageIntLLROutputS0xD(364)(5);
  VNStageIntLLRInputS0xD(55)(6) <= CNStageIntLLROutputS0xD(365)(0);
  VNStageIntLLRInputS0xD(67)(3) <= CNStageIntLLROutputS0xD(365)(1);
  VNStageIntLLRInputS0xD(190)(4) <= CNStageIntLLROutputS0xD(365)(2);
  VNStageIntLLRInputS0xD(202)(5) <= CNStageIntLLROutputS0xD(365)(3);
  VNStageIntLLRInputS0xD(289)(6) <= CNStageIntLLROutputS0xD(365)(4);
  VNStageIntLLRInputS0xD(372)(5) <= CNStageIntLLROutputS0xD(365)(5);
  VNStageIntLLRInputS0xD(54)(5) <= CNStageIntLLROutputS0xD(366)(0);
  VNStageIntLLRInputS0xD(125)(3) <= CNStageIntLLROutputS0xD(366)(1);
  VNStageIntLLRInputS0xD(137)(6) <= CNStageIntLLROutputS0xD(366)(2);
  VNStageIntLLRInputS0xD(224)(6) <= CNStageIntLLROutputS0xD(366)(3);
  VNStageIntLLRInputS0xD(307)(6) <= CNStageIntLLROutputS0xD(366)(4);
  VNStageIntLLRInputS0xD(357)(6) <= CNStageIntLLROutputS0xD(366)(5);
  VNStageIntLLRInputS0xD(53)(5) <= CNStageIntLLROutputS0xD(367)(0);
  VNStageIntLLRInputS0xD(72)(5) <= CNStageIntLLROutputS0xD(367)(1);
  VNStageIntLLRInputS0xD(159)(4) <= CNStageIntLLROutputS0xD(367)(2);
  VNStageIntLLRInputS0xD(242)(6) <= CNStageIntLLROutputS0xD(367)(3);
  VNStageIntLLRInputS0xD(292)(6) <= CNStageIntLLROutputS0xD(367)(4);
  VNStageIntLLRInputS0xD(344)(6) <= CNStageIntLLROutputS0xD(367)(5);
  VNStageIntLLRInputS0xD(52)(4) <= CNStageIntLLROutputS0xD(368)(0);
  VNStageIntLLRInputS0xD(94)(4) <= CNStageIntLLROutputS0xD(368)(1);
  VNStageIntLLRInputS0xD(177)(6) <= CNStageIntLLROutputS0xD(368)(2);
  VNStageIntLLRInputS0xD(227)(6) <= CNStageIntLLROutputS0xD(368)(3);
  VNStageIntLLRInputS0xD(279)(5) <= CNStageIntLLROutputS0xD(368)(4);
  VNStageIntLLRInputS0xD(375)(5) <= CNStageIntLLROutputS0xD(368)(5);
  VNStageIntLLRInputS0xD(51)(5) <= CNStageIntLLROutputS0xD(369)(0);
  VNStageIntLLRInputS0xD(112)(6) <= CNStageIntLLROutputS0xD(369)(1);
  VNStageIntLLRInputS0xD(162)(6) <= CNStageIntLLROutputS0xD(369)(2);
  VNStageIntLLRInputS0xD(214)(6) <= CNStageIntLLROutputS0xD(369)(3);
  VNStageIntLLRInputS0xD(310)(5) <= CNStageIntLLROutputS0xD(369)(4);
  VNStageIntLLRInputS0xD(324)(6) <= CNStageIntLLROutputS0xD(369)(5);
  VNStageIntLLRInputS0xD(50)(6) <= CNStageIntLLROutputS0xD(370)(0);
  VNStageIntLLRInputS0xD(97)(6) <= CNStageIntLLROutputS0xD(370)(1);
  VNStageIntLLRInputS0xD(149)(6) <= CNStageIntLLROutputS0xD(370)(2);
  VNStageIntLLRInputS0xD(245)(6) <= CNStageIntLLROutputS0xD(370)(3);
  VNStageIntLLRInputS0xD(259)(4) <= CNStageIntLLROutputS0xD(370)(4);
  VNStageIntLLRInputS0xD(338)(4) <= CNStageIntLLROutputS0xD(370)(5);
  VNStageIntLLRInputS0xD(49)(6) <= CNStageIntLLROutputS0xD(371)(0);
  VNStageIntLLRInputS0xD(84)(5) <= CNStageIntLLROutputS0xD(371)(1);
  VNStageIntLLRInputS0xD(180)(4) <= CNStageIntLLROutputS0xD(371)(2);
  VNStageIntLLRInputS0xD(194)(6) <= CNStageIntLLROutputS0xD(371)(3);
  VNStageIntLLRInputS0xD(273)(5) <= CNStageIntLLROutputS0xD(371)(4);
  VNStageIntLLRInputS0xD(382)(5) <= CNStageIntLLROutputS0xD(371)(5);
  VNStageIntLLRInputS0xD(48)(3) <= CNStageIntLLROutputS0xD(372)(0);
  VNStageIntLLRInputS0xD(115)(6) <= CNStageIntLLROutputS0xD(372)(1);
  VNStageIntLLRInputS0xD(129)(6) <= CNStageIntLLROutputS0xD(372)(2);
  VNStageIntLLRInputS0xD(208)(5) <= CNStageIntLLROutputS0xD(372)(3);
  VNStageIntLLRInputS0xD(317)(3) <= CNStageIntLLROutputS0xD(372)(4);
  VNStageIntLLRInputS0xD(359)(6) <= CNStageIntLLROutputS0xD(372)(5);
  VNStageIntLLRInputS0xD(47)(3) <= CNStageIntLLROutputS0xD(373)(0);
  VNStageIntLLRInputS0xD(127)(6) <= CNStageIntLLROutputS0xD(373)(1);
  VNStageIntLLRInputS0xD(143)(6) <= CNStageIntLLROutputS0xD(373)(2);
  VNStageIntLLRInputS0xD(252)(5) <= CNStageIntLLROutputS0xD(373)(3);
  VNStageIntLLRInputS0xD(294)(6) <= CNStageIntLLROutputS0xD(373)(4);
  VNStageIntLLRInputS0xD(348)(6) <= CNStageIntLLROutputS0xD(373)(5);
  VNStageIntLLRInputS0xD(46)(6) <= CNStageIntLLROutputS0xD(374)(0);
  VNStageIntLLRInputS0xD(78)(6) <= CNStageIntLLROutputS0xD(374)(1);
  VNStageIntLLRInputS0xD(187)(5) <= CNStageIntLLROutputS0xD(374)(2);
  VNStageIntLLRInputS0xD(229)(4) <= CNStageIntLLROutputS0xD(374)(3);
  VNStageIntLLRInputS0xD(283)(6) <= CNStageIntLLROutputS0xD(374)(4);
  VNStageIntLLRInputS0xD(352)(6) <= CNStageIntLLROutputS0xD(374)(5);
  VNStageIntLLRInputS0xD(45)(6) <= CNStageIntLLROutputS0xD(375)(0);
  VNStageIntLLRInputS0xD(122)(5) <= CNStageIntLLROutputS0xD(375)(1);
  VNStageIntLLRInputS0xD(164)(5) <= CNStageIntLLROutputS0xD(375)(2);
  VNStageIntLLRInputS0xD(218)(6) <= CNStageIntLLROutputS0xD(375)(3);
  VNStageIntLLRInputS0xD(287)(6) <= CNStageIntLLROutputS0xD(375)(4);
  VNStageIntLLRInputS0xD(345)(5) <= CNStageIntLLROutputS0xD(375)(5);
  VNStageIntLLRInputS0xD(44)(6) <= CNStageIntLLROutputS0xD(376)(0);
  VNStageIntLLRInputS0xD(99)(6) <= CNStageIntLLROutputS0xD(376)(1);
  VNStageIntLLRInputS0xD(153)(6) <= CNStageIntLLROutputS0xD(376)(2);
  VNStageIntLLRInputS0xD(222)(3) <= CNStageIntLLROutputS0xD(376)(3);
  VNStageIntLLRInputS0xD(280)(6) <= CNStageIntLLROutputS0xD(376)(4);
  VNStageIntLLRInputS0xD(356)(5) <= CNStageIntLLROutputS0xD(376)(5);
  VNStageIntLLRInputS0xD(43)(5) <= CNStageIntLLROutputS0xD(377)(0);
  VNStageIntLLRInputS0xD(88)(6) <= CNStageIntLLROutputS0xD(377)(1);
  VNStageIntLLRInputS0xD(157)(5) <= CNStageIntLLROutputS0xD(377)(2);
  VNStageIntLLRInputS0xD(215)(6) <= CNStageIntLLROutputS0xD(377)(3);
  VNStageIntLLRInputS0xD(291)(5) <= CNStageIntLLROutputS0xD(377)(4);
  VNStageIntLLRInputS0xD(328)(4) <= CNStageIntLLROutputS0xD(377)(5);
  VNStageIntLLRInputS0xD(42)(6) <= CNStageIntLLROutputS0xD(378)(0);
  VNStageIntLLRInputS0xD(92)(6) <= CNStageIntLLROutputS0xD(378)(1);
  VNStageIntLLRInputS0xD(150)(5) <= CNStageIntLLROutputS0xD(378)(2);
  VNStageIntLLRInputS0xD(226)(2) <= CNStageIntLLROutputS0xD(378)(3);
  VNStageIntLLRInputS0xD(263)(6) <= CNStageIntLLROutputS0xD(378)(4);
  VNStageIntLLRInputS0xD(383)(6) <= CNStageIntLLROutputS0xD(378)(5);
  VNStageIntLLRInputS0xD(41)(6) <= CNStageIntLLROutputS0xD(379)(0);
  VNStageIntLLRInputS0xD(85)(5) <= CNStageIntLLROutputS0xD(379)(1);
  VNStageIntLLRInputS0xD(161)(6) <= CNStageIntLLROutputS0xD(379)(2);
  VNStageIntLLRInputS0xD(198)(6) <= CNStageIntLLROutputS0xD(379)(3);
  VNStageIntLLRInputS0xD(318)(3) <= CNStageIntLLROutputS0xD(379)(4);
  VNStageIntLLRInputS0xD(337)(6) <= CNStageIntLLROutputS0xD(379)(5);
  VNStageIntLLRInputS0xD(40)(4) <= CNStageIntLLROutputS0xD(380)(0);
  VNStageIntLLRInputS0xD(96)(5) <= CNStageIntLLROutputS0xD(380)(1);
  VNStageIntLLRInputS0xD(133)(4) <= CNStageIntLLROutputS0xD(380)(2);
  VNStageIntLLRInputS0xD(253)(5) <= CNStageIntLLROutputS0xD(380)(3);
  VNStageIntLLRInputS0xD(272)(6) <= CNStageIntLLROutputS0xD(380)(4);
  VNStageIntLLRInputS0xD(334)(4) <= CNStageIntLLROutputS0xD(380)(5);
  VNStageIntLLRInputS0xD(39)(6) <= CNStageIntLLROutputS0xD(381)(0);
  VNStageIntLLRInputS0xD(68)(5) <= CNStageIntLLROutputS0xD(381)(1);
  VNStageIntLLRInputS0xD(188)(4) <= CNStageIntLLROutputS0xD(381)(2);
  VNStageIntLLRInputS0xD(207)(5) <= CNStageIntLLROutputS0xD(381)(3);
  VNStageIntLLRInputS0xD(269)(5) <= CNStageIntLLROutputS0xD(381)(4);
  VNStageIntLLRInputS0xD(368)(2) <= CNStageIntLLROutputS0xD(381)(5);
  VNStageIntLLRInputS0xD(38)(6) <= CNStageIntLLROutputS0xD(382)(0);
  VNStageIntLLRInputS0xD(123)(4) <= CNStageIntLLROutputS0xD(382)(1);
  VNStageIntLLRInputS0xD(142)(4) <= CNStageIntLLROutputS0xD(382)(2);
  VNStageIntLLRInputS0xD(204)(6) <= CNStageIntLLROutputS0xD(382)(3);
  VNStageIntLLRInputS0xD(303)(6) <= CNStageIntLLROutputS0xD(382)(4);
  VNStageIntLLRInputS0xD(325)(6) <= CNStageIntLLROutputS0xD(382)(5);
  VNStageIntLLRInputS0xD(37)(6) <= CNStageIntLLROutputS0xD(383)(0);
  VNStageIntLLRInputS0xD(77)(4) <= CNStageIntLLROutputS0xD(383)(1);
  VNStageIntLLRInputS0xD(139)(6) <= CNStageIntLLROutputS0xD(383)(2);
  VNStageIntLLRInputS0xD(238)(6) <= CNStageIntLLROutputS0xD(383)(3);
  VNStageIntLLRInputS0xD(260)(5) <= CNStageIntLLROutputS0xD(383)(4);
  VNStageIntLLRInputS0xD(374)(6) <= CNStageIntLLROutputS0xD(383)(5);

  -- Check Nodes (Iteration 1)
  CNStageIntLLRInputS1xD(53)(0) <= VNStageIntLLROutputS0xD(0)(0);
  CNStageIntLLRInputS1xD(110)(0) <= VNStageIntLLROutputS0xD(0)(1);
  CNStageIntLLRInputS1xD(170)(0) <= VNStageIntLLROutputS0xD(0)(2);
  CNStageIntLLRInputS1xD(224)(0) <= VNStageIntLLROutputS0xD(0)(3);
  CNStageIntLLRInputS1xD(279)(0) <= VNStageIntLLROutputS0xD(0)(4);
  CNStageIntLLRInputS1xD(332)(0) <= VNStageIntLLROutputS0xD(0)(5);
  CNStageIntLLRInputS1xD(51)(0) <= VNStageIntLLROutputS0xD(1)(0);
  CNStageIntLLRInputS1xD(139)(0) <= VNStageIntLLROutputS0xD(1)(1);
  CNStageIntLLRInputS1xD(223)(0) <= VNStageIntLLROutputS0xD(1)(2);
  CNStageIntLLRInputS1xD(241)(0) <= VNStageIntLLROutputS0xD(1)(3);
  CNStageIntLLRInputS1xD(307)(0) <= VNStageIntLLROutputS0xD(1)(4);
  CNStageIntLLRInputS1xD(356)(0) <= VNStageIntLLROutputS0xD(1)(5);
  CNStageIntLLRInputS1xD(50)(0) <= VNStageIntLLROutputS0xD(2)(0);
  CNStageIntLLRInputS1xD(92)(0) <= VNStageIntLLROutputS0xD(2)(1);
  CNStageIntLLRInputS1xD(138)(0) <= VNStageIntLLROutputS0xD(2)(2);
  CNStageIntLLRInputS1xD(222)(0) <= VNStageIntLLROutputS0xD(2)(3);
  CNStageIntLLRInputS1xD(240)(0) <= VNStageIntLLROutputS0xD(2)(4);
  CNStageIntLLRInputS1xD(306)(0) <= VNStageIntLLROutputS0xD(2)(5);
  CNStageIntLLRInputS1xD(355)(0) <= VNStageIntLLROutputS0xD(2)(6);
  CNStageIntLLRInputS1xD(91)(0) <= VNStageIntLLROutputS0xD(3)(0);
  CNStageIntLLRInputS1xD(137)(0) <= VNStageIntLLROutputS0xD(3)(1);
  CNStageIntLLRInputS1xD(221)(0) <= VNStageIntLLROutputS0xD(3)(2);
  CNStageIntLLRInputS1xD(239)(0) <= VNStageIntLLROutputS0xD(3)(3);
  CNStageIntLLRInputS1xD(305)(0) <= VNStageIntLLROutputS0xD(3)(4);
  CNStageIntLLRInputS1xD(49)(0) <= VNStageIntLLROutputS0xD(4)(0);
  CNStageIntLLRInputS1xD(90)(0) <= VNStageIntLLROutputS0xD(4)(1);
  CNStageIntLLRInputS1xD(220)(0) <= VNStageIntLLROutputS0xD(4)(2);
  CNStageIntLLRInputS1xD(238)(0) <= VNStageIntLLROutputS0xD(4)(3);
  CNStageIntLLRInputS1xD(304)(0) <= VNStageIntLLROutputS0xD(4)(4);
  CNStageIntLLRInputS1xD(354)(0) <= VNStageIntLLROutputS0xD(4)(5);
  CNStageIntLLRInputS1xD(48)(0) <= VNStageIntLLROutputS0xD(5)(0);
  CNStageIntLLRInputS1xD(89)(0) <= VNStageIntLLROutputS0xD(5)(1);
  CNStageIntLLRInputS1xD(136)(0) <= VNStageIntLLROutputS0xD(5)(2);
  CNStageIntLLRInputS1xD(219)(0) <= VNStageIntLLROutputS0xD(5)(3);
  CNStageIntLLRInputS1xD(237)(0) <= VNStageIntLLROutputS0xD(5)(4);
  CNStageIntLLRInputS1xD(303)(0) <= VNStageIntLLROutputS0xD(5)(5);
  CNStageIntLLRInputS1xD(353)(0) <= VNStageIntLLROutputS0xD(5)(6);
  CNStageIntLLRInputS1xD(47)(0) <= VNStageIntLLROutputS0xD(6)(0);
  CNStageIntLLRInputS1xD(88)(0) <= VNStageIntLLROutputS0xD(6)(1);
  CNStageIntLLRInputS1xD(135)(0) <= VNStageIntLLROutputS0xD(6)(2);
  CNStageIntLLRInputS1xD(218)(0) <= VNStageIntLLROutputS0xD(6)(3);
  CNStageIntLLRInputS1xD(236)(0) <= VNStageIntLLROutputS0xD(6)(4);
  CNStageIntLLRInputS1xD(302)(0) <= VNStageIntLLROutputS0xD(6)(5);
  CNStageIntLLRInputS1xD(352)(0) <= VNStageIntLLROutputS0xD(6)(6);
  CNStageIntLLRInputS1xD(46)(0) <= VNStageIntLLROutputS0xD(7)(0);
  CNStageIntLLRInputS1xD(87)(0) <= VNStageIntLLROutputS0xD(7)(1);
  CNStageIntLLRInputS1xD(134)(0) <= VNStageIntLLROutputS0xD(7)(2);
  CNStageIntLLRInputS1xD(217)(0) <= VNStageIntLLROutputS0xD(7)(3);
  CNStageIntLLRInputS1xD(235)(0) <= VNStageIntLLROutputS0xD(7)(4);
  CNStageIntLLRInputS1xD(301)(0) <= VNStageIntLLROutputS0xD(7)(5);
  CNStageIntLLRInputS1xD(351)(0) <= VNStageIntLLROutputS0xD(7)(6);
  CNStageIntLLRInputS1xD(45)(0) <= VNStageIntLLROutputS0xD(8)(0);
  CNStageIntLLRInputS1xD(133)(0) <= VNStageIntLLROutputS0xD(8)(1);
  CNStageIntLLRInputS1xD(216)(0) <= VNStageIntLLROutputS0xD(8)(2);
  CNStageIntLLRInputS1xD(44)(0) <= VNStageIntLLROutputS0xD(9)(0);
  CNStageIntLLRInputS1xD(86)(0) <= VNStageIntLLROutputS0xD(9)(1);
  CNStageIntLLRInputS1xD(132)(0) <= VNStageIntLLROutputS0xD(9)(2);
  CNStageIntLLRInputS1xD(215)(0) <= VNStageIntLLROutputS0xD(9)(3);
  CNStageIntLLRInputS1xD(234)(0) <= VNStageIntLLROutputS0xD(9)(4);
  CNStageIntLLRInputS1xD(300)(0) <= VNStageIntLLROutputS0xD(9)(5);
  CNStageIntLLRInputS1xD(350)(0) <= VNStageIntLLROutputS0xD(9)(6);
  CNStageIntLLRInputS1xD(43)(0) <= VNStageIntLLROutputS0xD(10)(0);
  CNStageIntLLRInputS1xD(85)(0) <= VNStageIntLLROutputS0xD(10)(1);
  CNStageIntLLRInputS1xD(131)(0) <= VNStageIntLLROutputS0xD(10)(2);
  CNStageIntLLRInputS1xD(233)(0) <= VNStageIntLLROutputS0xD(10)(3);
  CNStageIntLLRInputS1xD(349)(0) <= VNStageIntLLROutputS0xD(10)(4);
  CNStageIntLLRInputS1xD(42)(0) <= VNStageIntLLROutputS0xD(11)(0);
  CNStageIntLLRInputS1xD(84)(0) <= VNStageIntLLROutputS0xD(11)(1);
  CNStageIntLLRInputS1xD(130)(0) <= VNStageIntLLROutputS0xD(11)(2);
  CNStageIntLLRInputS1xD(214)(0) <= VNStageIntLLROutputS0xD(11)(3);
  CNStageIntLLRInputS1xD(232)(0) <= VNStageIntLLROutputS0xD(11)(4);
  CNStageIntLLRInputS1xD(348)(0) <= VNStageIntLLROutputS0xD(11)(5);
  CNStageIntLLRInputS1xD(41)(0) <= VNStageIntLLROutputS0xD(12)(0);
  CNStageIntLLRInputS1xD(83)(0) <= VNStageIntLLROutputS0xD(12)(1);
  CNStageIntLLRInputS1xD(129)(0) <= VNStageIntLLROutputS0xD(12)(2);
  CNStageIntLLRInputS1xD(213)(0) <= VNStageIntLLROutputS0xD(12)(3);
  CNStageIntLLRInputS1xD(231)(0) <= VNStageIntLLROutputS0xD(12)(4);
  CNStageIntLLRInputS1xD(299)(0) <= VNStageIntLLROutputS0xD(12)(5);
  CNStageIntLLRInputS1xD(347)(0) <= VNStageIntLLROutputS0xD(12)(6);
  CNStageIntLLRInputS1xD(82)(0) <= VNStageIntLLROutputS0xD(13)(0);
  CNStageIntLLRInputS1xD(128)(0) <= VNStageIntLLROutputS0xD(13)(1);
  CNStageIntLLRInputS1xD(212)(0) <= VNStageIntLLROutputS0xD(13)(2);
  CNStageIntLLRInputS1xD(230)(0) <= VNStageIntLLROutputS0xD(13)(3);
  CNStageIntLLRInputS1xD(298)(0) <= VNStageIntLLROutputS0xD(13)(4);
  CNStageIntLLRInputS1xD(346)(0) <= VNStageIntLLROutputS0xD(13)(5);
  CNStageIntLLRInputS1xD(40)(0) <= VNStageIntLLROutputS0xD(14)(0);
  CNStageIntLLRInputS1xD(81)(0) <= VNStageIntLLROutputS0xD(14)(1);
  CNStageIntLLRInputS1xD(127)(0) <= VNStageIntLLROutputS0xD(14)(2);
  CNStageIntLLRInputS1xD(211)(0) <= VNStageIntLLROutputS0xD(14)(3);
  CNStageIntLLRInputS1xD(229)(0) <= VNStageIntLLROutputS0xD(14)(4);
  CNStageIntLLRInputS1xD(297)(0) <= VNStageIntLLROutputS0xD(14)(5);
  CNStageIntLLRInputS1xD(345)(0) <= VNStageIntLLROutputS0xD(14)(6);
  CNStageIntLLRInputS1xD(39)(0) <= VNStageIntLLROutputS0xD(15)(0);
  CNStageIntLLRInputS1xD(80)(0) <= VNStageIntLLROutputS0xD(15)(1);
  CNStageIntLLRInputS1xD(126)(0) <= VNStageIntLLROutputS0xD(15)(2);
  CNStageIntLLRInputS1xD(210)(0) <= VNStageIntLLROutputS0xD(15)(3);
  CNStageIntLLRInputS1xD(228)(0) <= VNStageIntLLROutputS0xD(15)(4);
  CNStageIntLLRInputS1xD(296)(0) <= VNStageIntLLROutputS0xD(15)(5);
  CNStageIntLLRInputS1xD(344)(0) <= VNStageIntLLROutputS0xD(15)(6);
  CNStageIntLLRInputS1xD(38)(0) <= VNStageIntLLROutputS0xD(16)(0);
  CNStageIntLLRInputS1xD(125)(0) <= VNStageIntLLROutputS0xD(16)(1);
  CNStageIntLLRInputS1xD(209)(0) <= VNStageIntLLROutputS0xD(16)(2);
  CNStageIntLLRInputS1xD(227)(0) <= VNStageIntLLROutputS0xD(16)(3);
  CNStageIntLLRInputS1xD(295)(0) <= VNStageIntLLROutputS0xD(16)(4);
  CNStageIntLLRInputS1xD(343)(0) <= VNStageIntLLROutputS0xD(16)(5);
  CNStageIntLLRInputS1xD(37)(0) <= VNStageIntLLROutputS0xD(17)(0);
  CNStageIntLLRInputS1xD(79)(0) <= VNStageIntLLROutputS0xD(17)(1);
  CNStageIntLLRInputS1xD(124)(0) <= VNStageIntLLROutputS0xD(17)(2);
  CNStageIntLLRInputS1xD(208)(0) <= VNStageIntLLROutputS0xD(17)(3);
  CNStageIntLLRInputS1xD(226)(0) <= VNStageIntLLROutputS0xD(17)(4);
  CNStageIntLLRInputS1xD(294)(0) <= VNStageIntLLROutputS0xD(17)(5);
  CNStageIntLLRInputS1xD(342)(0) <= VNStageIntLLROutputS0xD(17)(6);
  CNStageIntLLRInputS1xD(36)(0) <= VNStageIntLLROutputS0xD(18)(0);
  CNStageIntLLRInputS1xD(78)(0) <= VNStageIntLLROutputS0xD(18)(1);
  CNStageIntLLRInputS1xD(123)(0) <= VNStageIntLLROutputS0xD(18)(2);
  CNStageIntLLRInputS1xD(207)(0) <= VNStageIntLLROutputS0xD(18)(3);
  CNStageIntLLRInputS1xD(225)(0) <= VNStageIntLLROutputS0xD(18)(4);
  CNStageIntLLRInputS1xD(293)(0) <= VNStageIntLLROutputS0xD(18)(5);
  CNStageIntLLRInputS1xD(341)(0) <= VNStageIntLLROutputS0xD(18)(6);
  CNStageIntLLRInputS1xD(35)(0) <= VNStageIntLLROutputS0xD(19)(0);
  CNStageIntLLRInputS1xD(77)(0) <= VNStageIntLLROutputS0xD(19)(1);
  CNStageIntLLRInputS1xD(122)(0) <= VNStageIntLLROutputS0xD(19)(2);
  CNStageIntLLRInputS1xD(278)(0) <= VNStageIntLLROutputS0xD(19)(3);
  CNStageIntLLRInputS1xD(340)(0) <= VNStageIntLLROutputS0xD(19)(4);
  CNStageIntLLRInputS1xD(34)(0) <= VNStageIntLLROutputS0xD(20)(0);
  CNStageIntLLRInputS1xD(76)(0) <= VNStageIntLLROutputS0xD(20)(1);
  CNStageIntLLRInputS1xD(277)(0) <= VNStageIntLLROutputS0xD(20)(2);
  CNStageIntLLRInputS1xD(292)(0) <= VNStageIntLLROutputS0xD(20)(3);
  CNStageIntLLRInputS1xD(339)(0) <= VNStageIntLLROutputS0xD(20)(4);
  CNStageIntLLRInputS1xD(33)(0) <= VNStageIntLLROutputS0xD(21)(0);
  CNStageIntLLRInputS1xD(75)(0) <= VNStageIntLLROutputS0xD(21)(1);
  CNStageIntLLRInputS1xD(121)(0) <= VNStageIntLLROutputS0xD(21)(2);
  CNStageIntLLRInputS1xD(206)(0) <= VNStageIntLLROutputS0xD(21)(3);
  CNStageIntLLRInputS1xD(276)(0) <= VNStageIntLLROutputS0xD(21)(4);
  CNStageIntLLRInputS1xD(291)(0) <= VNStageIntLLROutputS0xD(21)(5);
  CNStageIntLLRInputS1xD(338)(0) <= VNStageIntLLROutputS0xD(21)(6);
  CNStageIntLLRInputS1xD(32)(0) <= VNStageIntLLROutputS0xD(22)(0);
  CNStageIntLLRInputS1xD(74)(0) <= VNStageIntLLROutputS0xD(22)(1);
  CNStageIntLLRInputS1xD(120)(0) <= VNStageIntLLROutputS0xD(22)(2);
  CNStageIntLLRInputS1xD(205)(0) <= VNStageIntLLROutputS0xD(22)(3);
  CNStageIntLLRInputS1xD(275)(0) <= VNStageIntLLROutputS0xD(22)(4);
  CNStageIntLLRInputS1xD(290)(0) <= VNStageIntLLROutputS0xD(22)(5);
  CNStageIntLLRInputS1xD(337)(0) <= VNStageIntLLROutputS0xD(22)(6);
  CNStageIntLLRInputS1xD(31)(0) <= VNStageIntLLROutputS0xD(23)(0);
  CNStageIntLLRInputS1xD(73)(0) <= VNStageIntLLROutputS0xD(23)(1);
  CNStageIntLLRInputS1xD(119)(0) <= VNStageIntLLROutputS0xD(23)(2);
  CNStageIntLLRInputS1xD(204)(0) <= VNStageIntLLROutputS0xD(23)(3);
  CNStageIntLLRInputS1xD(274)(0) <= VNStageIntLLROutputS0xD(23)(4);
  CNStageIntLLRInputS1xD(289)(0) <= VNStageIntLLROutputS0xD(23)(5);
  CNStageIntLLRInputS1xD(336)(0) <= VNStageIntLLROutputS0xD(23)(6);
  CNStageIntLLRInputS1xD(30)(0) <= VNStageIntLLROutputS0xD(24)(0);
  CNStageIntLLRInputS1xD(72)(0) <= VNStageIntLLROutputS0xD(24)(1);
  CNStageIntLLRInputS1xD(118)(0) <= VNStageIntLLROutputS0xD(24)(2);
  CNStageIntLLRInputS1xD(203)(0) <= VNStageIntLLROutputS0xD(24)(3);
  CNStageIntLLRInputS1xD(273)(0) <= VNStageIntLLROutputS0xD(24)(4);
  CNStageIntLLRInputS1xD(288)(0) <= VNStageIntLLROutputS0xD(24)(5);
  CNStageIntLLRInputS1xD(335)(0) <= VNStageIntLLROutputS0xD(24)(6);
  CNStageIntLLRInputS1xD(29)(0) <= VNStageIntLLROutputS0xD(25)(0);
  CNStageIntLLRInputS1xD(71)(0) <= VNStageIntLLROutputS0xD(25)(1);
  CNStageIntLLRInputS1xD(117)(0) <= VNStageIntLLROutputS0xD(25)(2);
  CNStageIntLLRInputS1xD(202)(0) <= VNStageIntLLROutputS0xD(25)(3);
  CNStageIntLLRInputS1xD(287)(0) <= VNStageIntLLROutputS0xD(25)(4);
  CNStageIntLLRInputS1xD(28)(0) <= VNStageIntLLROutputS0xD(26)(0);
  CNStageIntLLRInputS1xD(70)(0) <= VNStageIntLLROutputS0xD(26)(1);
  CNStageIntLLRInputS1xD(116)(0) <= VNStageIntLLROutputS0xD(26)(2);
  CNStageIntLLRInputS1xD(201)(0) <= VNStageIntLLROutputS0xD(26)(3);
  CNStageIntLLRInputS1xD(272)(0) <= VNStageIntLLROutputS0xD(26)(4);
  CNStageIntLLRInputS1xD(286)(0) <= VNStageIntLLROutputS0xD(26)(5);
  CNStageIntLLRInputS1xD(334)(0) <= VNStageIntLLROutputS0xD(26)(6);
  CNStageIntLLRInputS1xD(27)(0) <= VNStageIntLLROutputS0xD(27)(0);
  CNStageIntLLRInputS1xD(69)(0) <= VNStageIntLLROutputS0xD(27)(1);
  CNStageIntLLRInputS1xD(115)(0) <= VNStageIntLLROutputS0xD(27)(2);
  CNStageIntLLRInputS1xD(200)(0) <= VNStageIntLLROutputS0xD(27)(3);
  CNStageIntLLRInputS1xD(285)(0) <= VNStageIntLLROutputS0xD(27)(4);
  CNStageIntLLRInputS1xD(26)(0) <= VNStageIntLLROutputS0xD(28)(0);
  CNStageIntLLRInputS1xD(68)(0) <= VNStageIntLLROutputS0xD(28)(1);
  CNStageIntLLRInputS1xD(114)(0) <= VNStageIntLLROutputS0xD(28)(2);
  CNStageIntLLRInputS1xD(199)(0) <= VNStageIntLLROutputS0xD(28)(3);
  CNStageIntLLRInputS1xD(271)(0) <= VNStageIntLLROutputS0xD(28)(4);
  CNStageIntLLRInputS1xD(333)(0) <= VNStageIntLLROutputS0xD(28)(5);
  CNStageIntLLRInputS1xD(25)(0) <= VNStageIntLLROutputS0xD(29)(0);
  CNStageIntLLRInputS1xD(67)(0) <= VNStageIntLLROutputS0xD(29)(1);
  CNStageIntLLRInputS1xD(113)(0) <= VNStageIntLLROutputS0xD(29)(2);
  CNStageIntLLRInputS1xD(270)(0) <= VNStageIntLLROutputS0xD(29)(3);
  CNStageIntLLRInputS1xD(24)(0) <= VNStageIntLLROutputS0xD(30)(0);
  CNStageIntLLRInputS1xD(66)(0) <= VNStageIntLLROutputS0xD(30)(1);
  CNStageIntLLRInputS1xD(112)(0) <= VNStageIntLLROutputS0xD(30)(2);
  CNStageIntLLRInputS1xD(198)(0) <= VNStageIntLLROutputS0xD(30)(3);
  CNStageIntLLRInputS1xD(269)(0) <= VNStageIntLLROutputS0xD(30)(4);
  CNStageIntLLRInputS1xD(284)(0) <= VNStageIntLLROutputS0xD(30)(5);
  CNStageIntLLRInputS1xD(23)(0) <= VNStageIntLLROutputS0xD(31)(0);
  CNStageIntLLRInputS1xD(65)(0) <= VNStageIntLLROutputS0xD(31)(1);
  CNStageIntLLRInputS1xD(197)(0) <= VNStageIntLLROutputS0xD(31)(2);
  CNStageIntLLRInputS1xD(283)(0) <= VNStageIntLLROutputS0xD(31)(3);
  CNStageIntLLRInputS1xD(22)(0) <= VNStageIntLLROutputS0xD(32)(0);
  CNStageIntLLRInputS1xD(64)(0) <= VNStageIntLLROutputS0xD(32)(1);
  CNStageIntLLRInputS1xD(111)(0) <= VNStageIntLLROutputS0xD(32)(2);
  CNStageIntLLRInputS1xD(268)(0) <= VNStageIntLLROutputS0xD(32)(3);
  CNStageIntLLRInputS1xD(21)(0) <= VNStageIntLLROutputS0xD(33)(0);
  CNStageIntLLRInputS1xD(63)(0) <= VNStageIntLLROutputS0xD(33)(1);
  CNStageIntLLRInputS1xD(169)(0) <= VNStageIntLLROutputS0xD(33)(2);
  CNStageIntLLRInputS1xD(196)(0) <= VNStageIntLLROutputS0xD(33)(3);
  CNStageIntLLRInputS1xD(267)(0) <= VNStageIntLLROutputS0xD(33)(4);
  CNStageIntLLRInputS1xD(282)(0) <= VNStageIntLLROutputS0xD(33)(5);
  CNStageIntLLRInputS1xD(20)(0) <= VNStageIntLLROutputS0xD(34)(0);
  CNStageIntLLRInputS1xD(62)(0) <= VNStageIntLLROutputS0xD(34)(1);
  CNStageIntLLRInputS1xD(168)(0) <= VNStageIntLLROutputS0xD(34)(2);
  CNStageIntLLRInputS1xD(195)(0) <= VNStageIntLLROutputS0xD(34)(3);
  CNStageIntLLRInputS1xD(266)(0) <= VNStageIntLLROutputS0xD(34)(4);
  CNStageIntLLRInputS1xD(281)(0) <= VNStageIntLLROutputS0xD(34)(5);
  CNStageIntLLRInputS1xD(19)(0) <= VNStageIntLLROutputS0xD(35)(0);
  CNStageIntLLRInputS1xD(61)(0) <= VNStageIntLLROutputS0xD(35)(1);
  CNStageIntLLRInputS1xD(167)(0) <= VNStageIntLLROutputS0xD(35)(2);
  CNStageIntLLRInputS1xD(194)(0) <= VNStageIntLLROutputS0xD(35)(3);
  CNStageIntLLRInputS1xD(265)(0) <= VNStageIntLLROutputS0xD(35)(4);
  CNStageIntLLRInputS1xD(280)(0) <= VNStageIntLLROutputS0xD(35)(5);
  CNStageIntLLRInputS1xD(18)(0) <= VNStageIntLLROutputS0xD(36)(0);
  CNStageIntLLRInputS1xD(60)(0) <= VNStageIntLLROutputS0xD(36)(1);
  CNStageIntLLRInputS1xD(166)(0) <= VNStageIntLLROutputS0xD(36)(2);
  CNStageIntLLRInputS1xD(264)(0) <= VNStageIntLLROutputS0xD(36)(3);
  CNStageIntLLRInputS1xD(17)(0) <= VNStageIntLLROutputS0xD(37)(0);
  CNStageIntLLRInputS1xD(59)(0) <= VNStageIntLLROutputS0xD(37)(1);
  CNStageIntLLRInputS1xD(165)(0) <= VNStageIntLLROutputS0xD(37)(2);
  CNStageIntLLRInputS1xD(193)(0) <= VNStageIntLLROutputS0xD(37)(3);
  CNStageIntLLRInputS1xD(263)(0) <= VNStageIntLLROutputS0xD(37)(4);
  CNStageIntLLRInputS1xD(331)(0) <= VNStageIntLLROutputS0xD(37)(5);
  CNStageIntLLRInputS1xD(383)(0) <= VNStageIntLLROutputS0xD(37)(6);
  CNStageIntLLRInputS1xD(16)(0) <= VNStageIntLLROutputS0xD(38)(0);
  CNStageIntLLRInputS1xD(58)(0) <= VNStageIntLLROutputS0xD(38)(1);
  CNStageIntLLRInputS1xD(164)(0) <= VNStageIntLLROutputS0xD(38)(2);
  CNStageIntLLRInputS1xD(192)(0) <= VNStageIntLLROutputS0xD(38)(3);
  CNStageIntLLRInputS1xD(262)(0) <= VNStageIntLLROutputS0xD(38)(4);
  CNStageIntLLRInputS1xD(330)(0) <= VNStageIntLLROutputS0xD(38)(5);
  CNStageIntLLRInputS1xD(382)(0) <= VNStageIntLLROutputS0xD(38)(6);
  CNStageIntLLRInputS1xD(15)(0) <= VNStageIntLLROutputS0xD(39)(0);
  CNStageIntLLRInputS1xD(57)(0) <= VNStageIntLLROutputS0xD(39)(1);
  CNStageIntLLRInputS1xD(163)(0) <= VNStageIntLLROutputS0xD(39)(2);
  CNStageIntLLRInputS1xD(191)(0) <= VNStageIntLLROutputS0xD(39)(3);
  CNStageIntLLRInputS1xD(261)(0) <= VNStageIntLLROutputS0xD(39)(4);
  CNStageIntLLRInputS1xD(329)(0) <= VNStageIntLLROutputS0xD(39)(5);
  CNStageIntLLRInputS1xD(381)(0) <= VNStageIntLLROutputS0xD(39)(6);
  CNStageIntLLRInputS1xD(14)(0) <= VNStageIntLLROutputS0xD(40)(0);
  CNStageIntLLRInputS1xD(56)(0) <= VNStageIntLLROutputS0xD(40)(1);
  CNStageIntLLRInputS1xD(162)(0) <= VNStageIntLLROutputS0xD(40)(2);
  CNStageIntLLRInputS1xD(260)(0) <= VNStageIntLLROutputS0xD(40)(3);
  CNStageIntLLRInputS1xD(380)(0) <= VNStageIntLLROutputS0xD(40)(4);
  CNStageIntLLRInputS1xD(13)(0) <= VNStageIntLLROutputS0xD(41)(0);
  CNStageIntLLRInputS1xD(55)(0) <= VNStageIntLLROutputS0xD(41)(1);
  CNStageIntLLRInputS1xD(161)(0) <= VNStageIntLLROutputS0xD(41)(2);
  CNStageIntLLRInputS1xD(190)(0) <= VNStageIntLLROutputS0xD(41)(3);
  CNStageIntLLRInputS1xD(259)(0) <= VNStageIntLLROutputS0xD(41)(4);
  CNStageIntLLRInputS1xD(328)(0) <= VNStageIntLLROutputS0xD(41)(5);
  CNStageIntLLRInputS1xD(379)(0) <= VNStageIntLLROutputS0xD(41)(6);
  CNStageIntLLRInputS1xD(12)(0) <= VNStageIntLLROutputS0xD(42)(0);
  CNStageIntLLRInputS1xD(54)(0) <= VNStageIntLLROutputS0xD(42)(1);
  CNStageIntLLRInputS1xD(160)(0) <= VNStageIntLLROutputS0xD(42)(2);
  CNStageIntLLRInputS1xD(189)(0) <= VNStageIntLLROutputS0xD(42)(3);
  CNStageIntLLRInputS1xD(258)(0) <= VNStageIntLLROutputS0xD(42)(4);
  CNStageIntLLRInputS1xD(327)(0) <= VNStageIntLLROutputS0xD(42)(5);
  CNStageIntLLRInputS1xD(378)(0) <= VNStageIntLLROutputS0xD(42)(6);
  CNStageIntLLRInputS1xD(109)(0) <= VNStageIntLLROutputS0xD(43)(0);
  CNStageIntLLRInputS1xD(159)(0) <= VNStageIntLLROutputS0xD(43)(1);
  CNStageIntLLRInputS1xD(188)(0) <= VNStageIntLLROutputS0xD(43)(2);
  CNStageIntLLRInputS1xD(257)(0) <= VNStageIntLLROutputS0xD(43)(3);
  CNStageIntLLRInputS1xD(326)(0) <= VNStageIntLLROutputS0xD(43)(4);
  CNStageIntLLRInputS1xD(377)(0) <= VNStageIntLLROutputS0xD(43)(5);
  CNStageIntLLRInputS1xD(11)(0) <= VNStageIntLLROutputS0xD(44)(0);
  CNStageIntLLRInputS1xD(108)(0) <= VNStageIntLLROutputS0xD(44)(1);
  CNStageIntLLRInputS1xD(158)(0) <= VNStageIntLLROutputS0xD(44)(2);
  CNStageIntLLRInputS1xD(187)(0) <= VNStageIntLLROutputS0xD(44)(3);
  CNStageIntLLRInputS1xD(256)(0) <= VNStageIntLLROutputS0xD(44)(4);
  CNStageIntLLRInputS1xD(325)(0) <= VNStageIntLLROutputS0xD(44)(5);
  CNStageIntLLRInputS1xD(376)(0) <= VNStageIntLLROutputS0xD(44)(6);
  CNStageIntLLRInputS1xD(10)(0) <= VNStageIntLLROutputS0xD(45)(0);
  CNStageIntLLRInputS1xD(107)(0) <= VNStageIntLLROutputS0xD(45)(1);
  CNStageIntLLRInputS1xD(157)(0) <= VNStageIntLLROutputS0xD(45)(2);
  CNStageIntLLRInputS1xD(186)(0) <= VNStageIntLLROutputS0xD(45)(3);
  CNStageIntLLRInputS1xD(255)(0) <= VNStageIntLLROutputS0xD(45)(4);
  CNStageIntLLRInputS1xD(324)(0) <= VNStageIntLLROutputS0xD(45)(5);
  CNStageIntLLRInputS1xD(375)(0) <= VNStageIntLLROutputS0xD(45)(6);
  CNStageIntLLRInputS1xD(9)(0) <= VNStageIntLLROutputS0xD(46)(0);
  CNStageIntLLRInputS1xD(106)(0) <= VNStageIntLLROutputS0xD(46)(1);
  CNStageIntLLRInputS1xD(156)(0) <= VNStageIntLLROutputS0xD(46)(2);
  CNStageIntLLRInputS1xD(185)(0) <= VNStageIntLLROutputS0xD(46)(3);
  CNStageIntLLRInputS1xD(254)(0) <= VNStageIntLLROutputS0xD(46)(4);
  CNStageIntLLRInputS1xD(323)(0) <= VNStageIntLLROutputS0xD(46)(5);
  CNStageIntLLRInputS1xD(374)(0) <= VNStageIntLLROutputS0xD(46)(6);
  CNStageIntLLRInputS1xD(8)(0) <= VNStageIntLLROutputS0xD(47)(0);
  CNStageIntLLRInputS1xD(155)(0) <= VNStageIntLLROutputS0xD(47)(1);
  CNStageIntLLRInputS1xD(253)(0) <= VNStageIntLLROutputS0xD(47)(2);
  CNStageIntLLRInputS1xD(373)(0) <= VNStageIntLLROutputS0xD(47)(3);
  CNStageIntLLRInputS1xD(7)(0) <= VNStageIntLLROutputS0xD(48)(0);
  CNStageIntLLRInputS1xD(154)(0) <= VNStageIntLLROutputS0xD(48)(1);
  CNStageIntLLRInputS1xD(322)(0) <= VNStageIntLLROutputS0xD(48)(2);
  CNStageIntLLRInputS1xD(372)(0) <= VNStageIntLLROutputS0xD(48)(3);
  CNStageIntLLRInputS1xD(6)(0) <= VNStageIntLLROutputS0xD(49)(0);
  CNStageIntLLRInputS1xD(105)(0) <= VNStageIntLLROutputS0xD(49)(1);
  CNStageIntLLRInputS1xD(153)(0) <= VNStageIntLLROutputS0xD(49)(2);
  CNStageIntLLRInputS1xD(184)(0) <= VNStageIntLLROutputS0xD(49)(3);
  CNStageIntLLRInputS1xD(252)(0) <= VNStageIntLLROutputS0xD(49)(4);
  CNStageIntLLRInputS1xD(321)(0) <= VNStageIntLLROutputS0xD(49)(5);
  CNStageIntLLRInputS1xD(371)(0) <= VNStageIntLLROutputS0xD(49)(6);
  CNStageIntLLRInputS1xD(5)(0) <= VNStageIntLLROutputS0xD(50)(0);
  CNStageIntLLRInputS1xD(104)(0) <= VNStageIntLLROutputS0xD(50)(1);
  CNStageIntLLRInputS1xD(152)(0) <= VNStageIntLLROutputS0xD(50)(2);
  CNStageIntLLRInputS1xD(183)(0) <= VNStageIntLLROutputS0xD(50)(3);
  CNStageIntLLRInputS1xD(251)(0) <= VNStageIntLLROutputS0xD(50)(4);
  CNStageIntLLRInputS1xD(320)(0) <= VNStageIntLLROutputS0xD(50)(5);
  CNStageIntLLRInputS1xD(370)(0) <= VNStageIntLLROutputS0xD(50)(6);
  CNStageIntLLRInputS1xD(4)(0) <= VNStageIntLLROutputS0xD(51)(0);
  CNStageIntLLRInputS1xD(103)(0) <= VNStageIntLLROutputS0xD(51)(1);
  CNStageIntLLRInputS1xD(182)(0) <= VNStageIntLLROutputS0xD(51)(2);
  CNStageIntLLRInputS1xD(250)(0) <= VNStageIntLLROutputS0xD(51)(3);
  CNStageIntLLRInputS1xD(319)(0) <= VNStageIntLLROutputS0xD(51)(4);
  CNStageIntLLRInputS1xD(369)(0) <= VNStageIntLLROutputS0xD(51)(5);
  CNStageIntLLRInputS1xD(102)(0) <= VNStageIntLLROutputS0xD(52)(0);
  CNStageIntLLRInputS1xD(151)(0) <= VNStageIntLLROutputS0xD(52)(1);
  CNStageIntLLRInputS1xD(181)(0) <= VNStageIntLLROutputS0xD(52)(2);
  CNStageIntLLRInputS1xD(318)(0) <= VNStageIntLLROutputS0xD(52)(3);
  CNStageIntLLRInputS1xD(368)(0) <= VNStageIntLLROutputS0xD(52)(4);
  CNStageIntLLRInputS1xD(3)(0) <= VNStageIntLLROutputS0xD(53)(0);
  CNStageIntLLRInputS1xD(150)(0) <= VNStageIntLLROutputS0xD(53)(1);
  CNStageIntLLRInputS1xD(180)(0) <= VNStageIntLLROutputS0xD(53)(2);
  CNStageIntLLRInputS1xD(249)(0) <= VNStageIntLLROutputS0xD(53)(3);
  CNStageIntLLRInputS1xD(317)(0) <= VNStageIntLLROutputS0xD(53)(4);
  CNStageIntLLRInputS1xD(367)(0) <= VNStageIntLLROutputS0xD(53)(5);
  CNStageIntLLRInputS1xD(2)(0) <= VNStageIntLLROutputS0xD(54)(0);
  CNStageIntLLRInputS1xD(101)(0) <= VNStageIntLLROutputS0xD(54)(1);
  CNStageIntLLRInputS1xD(149)(0) <= VNStageIntLLROutputS0xD(54)(2);
  CNStageIntLLRInputS1xD(179)(0) <= VNStageIntLLROutputS0xD(54)(3);
  CNStageIntLLRInputS1xD(316)(0) <= VNStageIntLLROutputS0xD(54)(4);
  CNStageIntLLRInputS1xD(366)(0) <= VNStageIntLLROutputS0xD(54)(5);
  CNStageIntLLRInputS1xD(1)(0) <= VNStageIntLLROutputS0xD(55)(0);
  CNStageIntLLRInputS1xD(100)(0) <= VNStageIntLLROutputS0xD(55)(1);
  CNStageIntLLRInputS1xD(148)(0) <= VNStageIntLLROutputS0xD(55)(2);
  CNStageIntLLRInputS1xD(178)(0) <= VNStageIntLLROutputS0xD(55)(3);
  CNStageIntLLRInputS1xD(248)(0) <= VNStageIntLLROutputS0xD(55)(4);
  CNStageIntLLRInputS1xD(315)(0) <= VNStageIntLLROutputS0xD(55)(5);
  CNStageIntLLRInputS1xD(365)(0) <= VNStageIntLLROutputS0xD(55)(6);
  CNStageIntLLRInputS1xD(0)(0) <= VNStageIntLLROutputS0xD(56)(0);
  CNStageIntLLRInputS1xD(99)(0) <= VNStageIntLLROutputS0xD(56)(1);
  CNStageIntLLRInputS1xD(147)(0) <= VNStageIntLLROutputS0xD(56)(2);
  CNStageIntLLRInputS1xD(177)(0) <= VNStageIntLLROutputS0xD(56)(3);
  CNStageIntLLRInputS1xD(247)(0) <= VNStageIntLLROutputS0xD(56)(4);
  CNStageIntLLRInputS1xD(314)(0) <= VNStageIntLLROutputS0xD(56)(5);
  CNStageIntLLRInputS1xD(364)(0) <= VNStageIntLLROutputS0xD(56)(6);
  CNStageIntLLRInputS1xD(98)(0) <= VNStageIntLLROutputS0xD(57)(0);
  CNStageIntLLRInputS1xD(146)(0) <= VNStageIntLLROutputS0xD(57)(1);
  CNStageIntLLRInputS1xD(176)(0) <= VNStageIntLLROutputS0xD(57)(2);
  CNStageIntLLRInputS1xD(246)(0) <= VNStageIntLLROutputS0xD(57)(3);
  CNStageIntLLRInputS1xD(313)(0) <= VNStageIntLLROutputS0xD(57)(4);
  CNStageIntLLRInputS1xD(363)(0) <= VNStageIntLLROutputS0xD(57)(5);
  CNStageIntLLRInputS1xD(97)(0) <= VNStageIntLLROutputS0xD(58)(0);
  CNStageIntLLRInputS1xD(145)(0) <= VNStageIntLLROutputS0xD(58)(1);
  CNStageIntLLRInputS1xD(175)(0) <= VNStageIntLLROutputS0xD(58)(2);
  CNStageIntLLRInputS1xD(312)(0) <= VNStageIntLLROutputS0xD(58)(3);
  CNStageIntLLRInputS1xD(362)(0) <= VNStageIntLLROutputS0xD(58)(4);
  CNStageIntLLRInputS1xD(144)(0) <= VNStageIntLLROutputS0xD(59)(0);
  CNStageIntLLRInputS1xD(174)(0) <= VNStageIntLLROutputS0xD(59)(1);
  CNStageIntLLRInputS1xD(245)(0) <= VNStageIntLLROutputS0xD(59)(2);
  CNStageIntLLRInputS1xD(311)(0) <= VNStageIntLLROutputS0xD(59)(3);
  CNStageIntLLRInputS1xD(361)(0) <= VNStageIntLLROutputS0xD(59)(4);
  CNStageIntLLRInputS1xD(96)(0) <= VNStageIntLLROutputS0xD(60)(0);
  CNStageIntLLRInputS1xD(143)(0) <= VNStageIntLLROutputS0xD(60)(1);
  CNStageIntLLRInputS1xD(173)(0) <= VNStageIntLLROutputS0xD(60)(2);
  CNStageIntLLRInputS1xD(244)(0) <= VNStageIntLLROutputS0xD(60)(3);
  CNStageIntLLRInputS1xD(310)(0) <= VNStageIntLLROutputS0xD(60)(4);
  CNStageIntLLRInputS1xD(360)(0) <= VNStageIntLLROutputS0xD(60)(5);
  CNStageIntLLRInputS1xD(95)(0) <= VNStageIntLLROutputS0xD(61)(0);
  CNStageIntLLRInputS1xD(142)(0) <= VNStageIntLLROutputS0xD(61)(1);
  CNStageIntLLRInputS1xD(172)(0) <= VNStageIntLLROutputS0xD(61)(2);
  CNStageIntLLRInputS1xD(243)(0) <= VNStageIntLLROutputS0xD(61)(3);
  CNStageIntLLRInputS1xD(309)(0) <= VNStageIntLLROutputS0xD(61)(4);
  CNStageIntLLRInputS1xD(359)(0) <= VNStageIntLLROutputS0xD(61)(5);
  CNStageIntLLRInputS1xD(94)(0) <= VNStageIntLLROutputS0xD(62)(0);
  CNStageIntLLRInputS1xD(141)(0) <= VNStageIntLLROutputS0xD(62)(1);
  CNStageIntLLRInputS1xD(171)(0) <= VNStageIntLLROutputS0xD(62)(2);
  CNStageIntLLRInputS1xD(242)(0) <= VNStageIntLLROutputS0xD(62)(3);
  CNStageIntLLRInputS1xD(308)(0) <= VNStageIntLLROutputS0xD(62)(4);
  CNStageIntLLRInputS1xD(358)(0) <= VNStageIntLLROutputS0xD(62)(5);
  CNStageIntLLRInputS1xD(52)(0) <= VNStageIntLLROutputS0xD(63)(0);
  CNStageIntLLRInputS1xD(93)(0) <= VNStageIntLLROutputS0xD(63)(1);
  CNStageIntLLRInputS1xD(140)(0) <= VNStageIntLLROutputS0xD(63)(2);
  CNStageIntLLRInputS1xD(357)(0) <= VNStageIntLLROutputS0xD(63)(3);
  CNStageIntLLRInputS1xD(53)(1) <= VNStageIntLLROutputS0xD(64)(0);
  CNStageIntLLRInputS1xD(109)(1) <= VNStageIntLLROutputS0xD(64)(1);
  CNStageIntLLRInputS1xD(130)(1) <= VNStageIntLLROutputS0xD(64)(2);
  CNStageIntLLRInputS1xD(245)(1) <= VNStageIntLLROutputS0xD(64)(3);
  CNStageIntLLRInputS1xD(299)(1) <= VNStageIntLLROutputS0xD(64)(4);
  CNStageIntLLRInputS1xD(342)(1) <= VNStageIntLLROutputS0xD(64)(5);
  CNStageIntLLRInputS1xD(51)(1) <= VNStageIntLLROutputS0xD(65)(0);
  CNStageIntLLRInputS1xD(74)(1) <= VNStageIntLLROutputS0xD(65)(1);
  CNStageIntLLRInputS1xD(141)(1) <= VNStageIntLLROutputS0xD(65)(2);
  CNStageIntLLRInputS1xD(189)(1) <= VNStageIntLLROutputS0xD(65)(3);
  CNStageIntLLRInputS1xD(286)(1) <= VNStageIntLLROutputS0xD(65)(4);
  CNStageIntLLRInputS1xD(50)(1) <= VNStageIntLLROutputS0xD(66)(0);
  CNStageIntLLRInputS1xD(66)(1) <= VNStageIntLLROutputS0xD(66)(1);
  CNStageIntLLRInputS1xD(155)(1) <= VNStageIntLLROutputS0xD(66)(2);
  CNStageIntLLRInputS1xD(244)(1) <= VNStageIntLLROutputS0xD(66)(3);
  CNStageIntLLRInputS1xD(97)(1) <= VNStageIntLLROutputS0xD(67)(0);
  CNStageIntLLRInputS1xD(275)(1) <= VNStageIntLLROutputS0xD(67)(1);
  CNStageIntLLRInputS1xD(322)(1) <= VNStageIntLLROutputS0xD(67)(2);
  CNStageIntLLRInputS1xD(365)(1) <= VNStageIntLLROutputS0xD(67)(3);
  CNStageIntLLRInputS1xD(49)(1) <= VNStageIntLLROutputS0xD(68)(0);
  CNStageIntLLRInputS1xD(112)(1) <= VNStageIntLLROutputS0xD(68)(1);
  CNStageIntLLRInputS1xD(210)(1) <= VNStageIntLLROutputS0xD(68)(2);
  CNStageIntLLRInputS1xD(256)(1) <= VNStageIntLLROutputS0xD(68)(3);
  CNStageIntLLRInputS1xD(318)(1) <= VNStageIntLLROutputS0xD(68)(4);
  CNStageIntLLRInputS1xD(381)(1) <= VNStageIntLLROutputS0xD(68)(5);
  CNStageIntLLRInputS1xD(48)(1) <= VNStageIntLLROutputS0xD(69)(0);
  CNStageIntLLRInputS1xD(101)(1) <= VNStageIntLLROutputS0xD(69)(1);
  CNStageIntLLRInputS1xD(135)(1) <= VNStageIntLLROutputS0xD(69)(2);
  CNStageIntLLRInputS1xD(215)(1) <= VNStageIntLLROutputS0xD(69)(3);
  CNStageIntLLRInputS1xD(259)(1) <= VNStageIntLLROutputS0xD(69)(4);
  CNStageIntLLRInputS1xD(283)(1) <= VNStageIntLLROutputS0xD(69)(5);
  CNStageIntLLRInputS1xD(351)(1) <= VNStageIntLLROutputS0xD(69)(6);
  CNStageIntLLRInputS1xD(47)(1) <= VNStageIntLLROutputS0xD(70)(0);
  CNStageIntLLRInputS1xD(104)(1) <= VNStageIntLLROutputS0xD(70)(1);
  CNStageIntLLRInputS1xD(136)(1) <= VNStageIntLLROutputS0xD(70)(2);
  CNStageIntLLRInputS1xD(206)(1) <= VNStageIntLLROutputS0xD(70)(3);
  CNStageIntLLRInputS1xD(246)(1) <= VNStageIntLLROutputS0xD(70)(4);
  CNStageIntLLRInputS1xD(301)(1) <= VNStageIntLLROutputS0xD(70)(5);
  CNStageIntLLRInputS1xD(46)(1) <= VNStageIntLLROutputS0xD(71)(0);
  CNStageIntLLRInputS1xD(95)(1) <= VNStageIntLLROutputS0xD(71)(1);
  CNStageIntLLRInputS1xD(176)(1) <= VNStageIntLLROutputS0xD(71)(2);
  CNStageIntLLRInputS1xD(276)(1) <= VNStageIntLLROutputS0xD(71)(3);
  CNStageIntLLRInputS1xD(302)(1) <= VNStageIntLLROutputS0xD(71)(4);
  CNStageIntLLRInputS1xD(353)(1) <= VNStageIntLLROutputS0xD(71)(5);
  CNStageIntLLRInputS1xD(45)(1) <= VNStageIntLLROutputS0xD(72)(0);
  CNStageIntLLRInputS1xD(75)(1) <= VNStageIntLLROutputS0xD(72)(1);
  CNStageIntLLRInputS1xD(162)(1) <= VNStageIntLLROutputS0xD(72)(2);
  CNStageIntLLRInputS1xD(183)(1) <= VNStageIntLLROutputS0xD(72)(3);
  CNStageIntLLRInputS1xD(243)(1) <= VNStageIntLLROutputS0xD(72)(4);
  CNStageIntLLRInputS1xD(367)(1) <= VNStageIntLLROutputS0xD(72)(5);
  CNStageIntLLRInputS1xD(44)(1) <= VNStageIntLLROutputS0xD(73)(0);
  CNStageIntLLRInputS1xD(56)(1) <= VNStageIntLLROutputS0xD(73)(1);
  CNStageIntLLRInputS1xD(121)(1) <= VNStageIntLLROutputS0xD(73)(2);
  CNStageIntLLRInputS1xD(219)(1) <= VNStageIntLLROutputS0xD(73)(3);
  CNStageIntLLRInputS1xD(328)(1) <= VNStageIntLLROutputS0xD(73)(4);
  CNStageIntLLRInputS1xD(363)(1) <= VNStageIntLLROutputS0xD(73)(5);
  CNStageIntLLRInputS1xD(43)(1) <= VNStageIntLLROutputS0xD(74)(0);
  CNStageIntLLRInputS1xD(70)(1) <= VNStageIntLLROutputS0xD(74)(1);
  CNStageIntLLRInputS1xD(125)(1) <= VNStageIntLLROutputS0xD(74)(2);
  CNStageIntLLRInputS1xD(221)(1) <= VNStageIntLLROutputS0xD(74)(3);
  CNStageIntLLRInputS1xD(290)(1) <= VNStageIntLLROutputS0xD(74)(4);
  CNStageIntLLRInputS1xD(42)(1) <= VNStageIntLLROutputS0xD(75)(0);
  CNStageIntLLRInputS1xD(81)(1) <= VNStageIntLLROutputS0xD(75)(1);
  CNStageIntLLRInputS1xD(170)(1) <= VNStageIntLLROutputS0xD(75)(2);
  CNStageIntLLRInputS1xD(192)(1) <= VNStageIntLLROutputS0xD(75)(3);
  CNStageIntLLRInputS1xD(278)(1) <= VNStageIntLLROutputS0xD(75)(4);
  CNStageIntLLRInputS1xD(294)(1) <= VNStageIntLLROutputS0xD(75)(5);
  CNStageIntLLRInputS1xD(347)(1) <= VNStageIntLLROutputS0xD(75)(6);
  CNStageIntLLRInputS1xD(41)(1) <= VNStageIntLLROutputS0xD(76)(0);
  CNStageIntLLRInputS1xD(106)(1) <= VNStageIntLLROutputS0xD(76)(1);
  CNStageIntLLRInputS1xD(124)(1) <= VNStageIntLLROutputS0xD(76)(2);
  CNStageIntLLRInputS1xD(174)(1) <= VNStageIntLLROutputS0xD(76)(3);
  CNStageIntLLRInputS1xD(270)(1) <= VNStageIntLLROutputS0xD(76)(4);
  CNStageIntLLRInputS1xD(332)(1) <= VNStageIntLLROutputS0xD(76)(5);
  CNStageIntLLRInputS1xD(348)(1) <= VNStageIntLLROutputS0xD(76)(6);
  CNStageIntLLRInputS1xD(119)(1) <= VNStageIntLLROutputS0xD(77)(0);
  CNStageIntLLRInputS1xD(185)(1) <= VNStageIntLLROutputS0xD(77)(1);
  CNStageIntLLRInputS1xD(257)(1) <= VNStageIntLLROutputS0xD(77)(2);
  CNStageIntLLRInputS1xD(293)(1) <= VNStageIntLLROutputS0xD(77)(3);
  CNStageIntLLRInputS1xD(383)(1) <= VNStageIntLLROutputS0xD(77)(4);
  CNStageIntLLRInputS1xD(40)(1) <= VNStageIntLLROutputS0xD(78)(0);
  CNStageIntLLRInputS1xD(84)(1) <= VNStageIntLLROutputS0xD(78)(1);
  CNStageIntLLRInputS1xD(159)(1) <= VNStageIntLLROutputS0xD(78)(2);
  CNStageIntLLRInputS1xD(193)(1) <= VNStageIntLLROutputS0xD(78)(3);
  CNStageIntLLRInputS1xD(274)(1) <= VNStageIntLLROutputS0xD(78)(4);
  CNStageIntLLRInputS1xD(288)(1) <= VNStageIntLLROutputS0xD(78)(5);
  CNStageIntLLRInputS1xD(374)(1) <= VNStageIntLLROutputS0xD(78)(6);
  CNStageIntLLRInputS1xD(39)(1) <= VNStageIntLLROutputS0xD(79)(0);
  CNStageIntLLRInputS1xD(99)(1) <= VNStageIntLLROutputS0xD(79)(1);
  CNStageIntLLRInputS1xD(167)(1) <= VNStageIntLLROutputS0xD(79)(2);
  CNStageIntLLRInputS1xD(220)(1) <= VNStageIntLLROutputS0xD(79)(3);
  CNStageIntLLRInputS1xD(325)(1) <= VNStageIntLLROutputS0xD(79)(4);
  CNStageIntLLRInputS1xD(38)(1) <= VNStageIntLLROutputS0xD(80)(0);
  CNStageIntLLRInputS1xD(62)(1) <= VNStageIntLLROutputS0xD(80)(1);
  CNStageIntLLRInputS1xD(131)(1) <= VNStageIntLLROutputS0xD(80)(2);
  CNStageIntLLRInputS1xD(182)(1) <= VNStageIntLLROutputS0xD(80)(3);
  CNStageIntLLRInputS1xD(248)(1) <= VNStageIntLLROutputS0xD(80)(4);
  CNStageIntLLRInputS1xD(337)(1) <= VNStageIntLLROutputS0xD(80)(5);
  CNStageIntLLRInputS1xD(37)(1) <= VNStageIntLLROutputS0xD(81)(0);
  CNStageIntLLRInputS1xD(72)(1) <= VNStageIntLLROutputS0xD(81)(1);
  CNStageIntLLRInputS1xD(129)(1) <= VNStageIntLLROutputS0xD(81)(2);
  CNStageIntLLRInputS1xD(262)(1) <= VNStageIntLLROutputS0xD(81)(3);
  CNStageIntLLRInputS1xD(36)(1) <= VNStageIntLLROutputS0xD(82)(0);
  CNStageIntLLRInputS1xD(67)(1) <= VNStageIntLLROutputS0xD(82)(1);
  CNStageIntLLRInputS1xD(165)(1) <= VNStageIntLLROutputS0xD(82)(2);
  CNStageIntLLRInputS1xD(188)(1) <= VNStageIntLLROutputS0xD(82)(3);
  CNStageIntLLRInputS1xD(254)(1) <= VNStageIntLLROutputS0xD(82)(4);
  CNStageIntLLRInputS1xD(298)(1) <= VNStageIntLLROutputS0xD(82)(5);
  CNStageIntLLRInputS1xD(336)(1) <= VNStageIntLLROutputS0xD(82)(6);
  CNStageIntLLRInputS1xD(35)(1) <= VNStageIntLLROutputS0xD(83)(0);
  CNStageIntLLRInputS1xD(73)(1) <= VNStageIntLLROutputS0xD(83)(1);
  CNStageIntLLRInputS1xD(144)(1) <= VNStageIntLLROutputS0xD(83)(2);
  CNStageIntLLRInputS1xD(208)(1) <= VNStageIntLLROutputS0xD(83)(3);
  CNStageIntLLRInputS1xD(232)(1) <= VNStageIntLLROutputS0xD(83)(4);
  CNStageIntLLRInputS1xD(330)(1) <= VNStageIntLLROutputS0xD(83)(5);
  CNStageIntLLRInputS1xD(34)(1) <= VNStageIntLLROutputS0xD(84)(0);
  CNStageIntLLRInputS1xD(61)(1) <= VNStageIntLLROutputS0xD(84)(1);
  CNStageIntLLRInputS1xD(147)(1) <= VNStageIntLLROutputS0xD(84)(2);
  CNStageIntLLRInputS1xD(222)(1) <= VNStageIntLLROutputS0xD(84)(3);
  CNStageIntLLRInputS1xD(310)(1) <= VNStageIntLLROutputS0xD(84)(4);
  CNStageIntLLRInputS1xD(371)(1) <= VNStageIntLLROutputS0xD(84)(5);
  CNStageIntLLRInputS1xD(33)(1) <= VNStageIntLLROutputS0xD(85)(0);
  CNStageIntLLRInputS1xD(132)(1) <= VNStageIntLLROutputS0xD(85)(1);
  CNStageIntLLRInputS1xD(218)(1) <= VNStageIntLLROutputS0xD(85)(2);
  CNStageIntLLRInputS1xD(235)(1) <= VNStageIntLLROutputS0xD(85)(3);
  CNStageIntLLRInputS1xD(313)(1) <= VNStageIntLLROutputS0xD(85)(4);
  CNStageIntLLRInputS1xD(379)(1) <= VNStageIntLLROutputS0xD(85)(5);
  CNStageIntLLRInputS1xD(32)(1) <= VNStageIntLLROutputS0xD(86)(0);
  CNStageIntLLRInputS1xD(166)(1) <= VNStageIntLLROutputS0xD(86)(1);
  CNStageIntLLRInputS1xD(239)(1) <= VNStageIntLLROutputS0xD(86)(2);
  CNStageIntLLRInputS1xD(343)(1) <= VNStageIntLLROutputS0xD(86)(3);
  CNStageIntLLRInputS1xD(31)(1) <= VNStageIntLLROutputS0xD(87)(0);
  CNStageIntLLRInputS1xD(77)(1) <= VNStageIntLLROutputS0xD(87)(1);
  CNStageIntLLRInputS1xD(128)(1) <= VNStageIntLLROutputS0xD(87)(2);
  CNStageIntLLRInputS1xD(203)(1) <= VNStageIntLLROutputS0xD(87)(3);
  CNStageIntLLRInputS1xD(229)(1) <= VNStageIntLLROutputS0xD(87)(4);
  CNStageIntLLRInputS1xD(331)(1) <= VNStageIntLLROutputS0xD(87)(5);
  CNStageIntLLRInputS1xD(341)(1) <= VNStageIntLLROutputS0xD(87)(6);
  CNStageIntLLRInputS1xD(30)(1) <= VNStageIntLLROutputS0xD(88)(0);
  CNStageIntLLRInputS1xD(79)(1) <= VNStageIntLLROutputS0xD(88)(1);
  CNStageIntLLRInputS1xD(156)(1) <= VNStageIntLLROutputS0xD(88)(2);
  CNStageIntLLRInputS1xD(204)(1) <= VNStageIntLLROutputS0xD(88)(3);
  CNStageIntLLRInputS1xD(263)(1) <= VNStageIntLLROutputS0xD(88)(4);
  CNStageIntLLRInputS1xD(297)(1) <= VNStageIntLLROutputS0xD(88)(5);
  CNStageIntLLRInputS1xD(377)(1) <= VNStageIntLLROutputS0xD(88)(6);
  CNStageIntLLRInputS1xD(29)(1) <= VNStageIntLLROutputS0xD(89)(0);
  CNStageIntLLRInputS1xD(102)(1) <= VNStageIntLLROutputS0xD(89)(1);
  CNStageIntLLRInputS1xD(140)(1) <= VNStageIntLLROutputS0xD(89)(2);
  CNStageIntLLRInputS1xD(184)(1) <= VNStageIntLLROutputS0xD(89)(3);
  CNStageIntLLRInputS1xD(247)(1) <= VNStageIntLLROutputS0xD(89)(4);
  CNStageIntLLRInputS1xD(355)(1) <= VNStageIntLLROutputS0xD(89)(5);
  CNStageIntLLRInputS1xD(28)(1) <= VNStageIntLLROutputS0xD(90)(0);
  CNStageIntLLRInputS1xD(85)(1) <= VNStageIntLLROutputS0xD(90)(1);
  CNStageIntLLRInputS1xD(168)(1) <= VNStageIntLLROutputS0xD(90)(2);
  CNStageIntLLRInputS1xD(175)(1) <= VNStageIntLLROutputS0xD(90)(3);
  CNStageIntLLRInputS1xD(258)(1) <= VNStageIntLLROutputS0xD(90)(4);
  CNStageIntLLRInputS1xD(307)(1) <= VNStageIntLLROutputS0xD(90)(5);
  CNStageIntLLRInputS1xD(358)(1) <= VNStageIntLLROutputS0xD(90)(6);
  CNStageIntLLRInputS1xD(27)(1) <= VNStageIntLLROutputS0xD(91)(0);
  CNStageIntLLRInputS1xD(96)(1) <= VNStageIntLLROutputS0xD(91)(1);
  CNStageIntLLRInputS1xD(158)(1) <= VNStageIntLLROutputS0xD(91)(2);
  CNStageIntLLRInputS1xD(191)(1) <= VNStageIntLLROutputS0xD(91)(3);
  CNStageIntLLRInputS1xD(269)(1) <= VNStageIntLLROutputS0xD(91)(4);
  CNStageIntLLRInputS1xD(280)(1) <= VNStageIntLLROutputS0xD(91)(5);
  CNStageIntLLRInputS1xD(344)(1) <= VNStageIntLLROutputS0xD(91)(6);
  CNStageIntLLRInputS1xD(26)(1) <= VNStageIntLLROutputS0xD(92)(0);
  CNStageIntLLRInputS1xD(103)(1) <= VNStageIntLLROutputS0xD(92)(1);
  CNStageIntLLRInputS1xD(145)(1) <= VNStageIntLLROutputS0xD(92)(2);
  CNStageIntLLRInputS1xD(195)(1) <= VNStageIntLLROutputS0xD(92)(3);
  CNStageIntLLRInputS1xD(242)(1) <= VNStageIntLLROutputS0xD(92)(4);
  CNStageIntLLRInputS1xD(324)(1) <= VNStageIntLLROutputS0xD(92)(5);
  CNStageIntLLRInputS1xD(378)(1) <= VNStageIntLLROutputS0xD(92)(6);
  CNStageIntLLRInputS1xD(25)(1) <= VNStageIntLLROutputS0xD(93)(0);
  CNStageIntLLRInputS1xD(78)(1) <= VNStageIntLLROutputS0xD(93)(1);
  CNStageIntLLRInputS1xD(164)(1) <= VNStageIntLLROutputS0xD(93)(2);
  CNStageIntLLRInputS1xD(224)(1) <= VNStageIntLLROutputS0xD(93)(3);
  CNStageIntLLRInputS1xD(231)(1) <= VNStageIntLLROutputS0xD(93)(4);
  CNStageIntLLRInputS1xD(311)(1) <= VNStageIntLLROutputS0xD(93)(5);
  CNStageIntLLRInputS1xD(340)(1) <= VNStageIntLLROutputS0xD(93)(6);
  CNStageIntLLRInputS1xD(24)(1) <= VNStageIntLLROutputS0xD(94)(0);
  CNStageIntLLRInputS1xD(92)(1) <= VNStageIntLLROutputS0xD(94)(1);
  CNStageIntLLRInputS1xD(194)(1) <= VNStageIntLLROutputS0xD(94)(2);
  CNStageIntLLRInputS1xD(329)(1) <= VNStageIntLLROutputS0xD(94)(3);
  CNStageIntLLRInputS1xD(368)(1) <= VNStageIntLLROutputS0xD(94)(4);
  CNStageIntLLRInputS1xD(23)(1) <= VNStageIntLLROutputS0xD(95)(0);
  CNStageIntLLRInputS1xD(63)(1) <= VNStageIntLLROutputS0xD(95)(1);
  CNStageIntLLRInputS1xD(134)(1) <= VNStageIntLLROutputS0xD(95)(2);
  CNStageIntLLRInputS1xD(190)(1) <= VNStageIntLLROutputS0xD(95)(3);
  CNStageIntLLRInputS1xD(234)(1) <= VNStageIntLLROutputS0xD(95)(4);
  CNStageIntLLRInputS1xD(303)(1) <= VNStageIntLLROutputS0xD(95)(5);
  CNStageIntLLRInputS1xD(352)(1) <= VNStageIntLLROutputS0xD(95)(6);
  CNStageIntLLRInputS1xD(22)(1) <= VNStageIntLLROutputS0xD(96)(0);
  CNStageIntLLRInputS1xD(98)(1) <= VNStageIntLLROutputS0xD(96)(1);
  CNStageIntLLRInputS1xD(150)(1) <= VNStageIntLLROutputS0xD(96)(2);
  CNStageIntLLRInputS1xD(172)(1) <= VNStageIntLLROutputS0xD(96)(3);
  CNStageIntLLRInputS1xD(251)(1) <= VNStageIntLLROutputS0xD(96)(4);
  CNStageIntLLRInputS1xD(380)(1) <= VNStageIntLLROutputS0xD(96)(5);
  CNStageIntLLRInputS1xD(21)(1) <= VNStageIntLLROutputS0xD(97)(0);
  CNStageIntLLRInputS1xD(65)(1) <= VNStageIntLLROutputS0xD(97)(1);
  CNStageIntLLRInputS1xD(142)(1) <= VNStageIntLLROutputS0xD(97)(2);
  CNStageIntLLRInputS1xD(180)(1) <= VNStageIntLLROutputS0xD(97)(3);
  CNStageIntLLRInputS1xD(260)(1) <= VNStageIntLLROutputS0xD(97)(4);
  CNStageIntLLRInputS1xD(316)(1) <= VNStageIntLLROutputS0xD(97)(5);
  CNStageIntLLRInputS1xD(370)(1) <= VNStageIntLLROutputS0xD(97)(6);
  CNStageIntLLRInputS1xD(20)(1) <= VNStageIntLLROutputS0xD(98)(0);
  CNStageIntLLRInputS1xD(116)(1) <= VNStageIntLLROutputS0xD(98)(1);
  CNStageIntLLRInputS1xD(199)(1) <= VNStageIntLLROutputS0xD(98)(2);
  CNStageIntLLRInputS1xD(255)(1) <= VNStageIntLLROutputS0xD(98)(3);
  CNStageIntLLRInputS1xD(308)(1) <= VNStageIntLLROutputS0xD(98)(4);
  CNStageIntLLRInputS1xD(356)(1) <= VNStageIntLLROutputS0xD(98)(5);
  CNStageIntLLRInputS1xD(19)(1) <= VNStageIntLLROutputS0xD(99)(0);
  CNStageIntLLRInputS1xD(76)(1) <= VNStageIntLLROutputS0xD(99)(1);
  CNStageIntLLRInputS1xD(126)(1) <= VNStageIntLLROutputS0xD(99)(2);
  CNStageIntLLRInputS1xD(198)(1) <= VNStageIntLLROutputS0xD(99)(3);
  CNStageIntLLRInputS1xD(261)(1) <= VNStageIntLLROutputS0xD(99)(4);
  CNStageIntLLRInputS1xD(285)(1) <= VNStageIntLLROutputS0xD(99)(5);
  CNStageIntLLRInputS1xD(376)(1) <= VNStageIntLLROutputS0xD(99)(6);
  CNStageIntLLRInputS1xD(18)(1) <= VNStageIntLLROutputS0xD(100)(0);
  CNStageIntLLRInputS1xD(94)(1) <= VNStageIntLLROutputS0xD(100)(1);
  CNStageIntLLRInputS1xD(120)(1) <= VNStageIntLLROutputS0xD(100)(2);
  CNStageIntLLRInputS1xD(178)(1) <= VNStageIntLLROutputS0xD(100)(3);
  CNStageIntLLRInputS1xD(250)(1) <= VNStageIntLLROutputS0xD(100)(4);
  CNStageIntLLRInputS1xD(295)(1) <= VNStageIntLLROutputS0xD(100)(5);
  CNStageIntLLRInputS1xD(349)(1) <= VNStageIntLLROutputS0xD(100)(6);
  CNStageIntLLRInputS1xD(17)(1) <= VNStageIntLLROutputS0xD(101)(0);
  CNStageIntLLRInputS1xD(58)(1) <= VNStageIntLLROutputS0xD(101)(1);
  CNStageIntLLRInputS1xD(123)(1) <= VNStageIntLLROutputS0xD(101)(2);
  CNStageIntLLRInputS1xD(211)(1) <= VNStageIntLLROutputS0xD(101)(3);
  CNStageIntLLRInputS1xD(273)(1) <= VNStageIntLLROutputS0xD(101)(4);
  CNStageIntLLRInputS1xD(289)(1) <= VNStageIntLLROutputS0xD(101)(5);
  CNStageIntLLRInputS1xD(346)(1) <= VNStageIntLLROutputS0xD(101)(6);
  CNStageIntLLRInputS1xD(16)(1) <= VNStageIntLLROutputS0xD(102)(0);
  CNStageIntLLRInputS1xD(59)(1) <= VNStageIntLLROutputS0xD(102)(1);
  CNStageIntLLRInputS1xD(113)(1) <= VNStageIntLLROutputS0xD(102)(2);
  CNStageIntLLRInputS1xD(214)(1) <= VNStageIntLLROutputS0xD(102)(3);
  CNStageIntLLRInputS1xD(226)(1) <= VNStageIntLLROutputS0xD(102)(4);
  CNStageIntLLRInputS1xD(361)(1) <= VNStageIntLLROutputS0xD(102)(5);
  CNStageIntLLRInputS1xD(15)(1) <= VNStageIntLLROutputS0xD(103)(0);
  CNStageIntLLRInputS1xD(93)(1) <= VNStageIntLLROutputS0xD(103)(1);
  CNStageIntLLRInputS1xD(151)(1) <= VNStageIntLLROutputS0xD(103)(2);
  CNStageIntLLRInputS1xD(200)(1) <= VNStageIntLLROutputS0xD(103)(3);
  CNStageIntLLRInputS1xD(265)(1) <= VNStageIntLLROutputS0xD(103)(4);
  CNStageIntLLRInputS1xD(284)(1) <= VNStageIntLLROutputS0xD(103)(5);
  CNStageIntLLRInputS1xD(354)(1) <= VNStageIntLLROutputS0xD(103)(6);
  CNStageIntLLRInputS1xD(14)(1) <= VNStageIntLLROutputS0xD(104)(0);
  CNStageIntLLRInputS1xD(86)(1) <= VNStageIntLLROutputS0xD(104)(1);
  CNStageIntLLRInputS1xD(133)(1) <= VNStageIntLLROutputS0xD(104)(2);
  CNStageIntLLRInputS1xD(179)(1) <= VNStageIntLLROutputS0xD(104)(3);
  CNStageIntLLRInputS1xD(267)(1) <= VNStageIntLLROutputS0xD(104)(4);
  CNStageIntLLRInputS1xD(317)(1) <= VNStageIntLLROutputS0xD(104)(5);
  CNStageIntLLRInputS1xD(13)(1) <= VNStageIntLLROutputS0xD(105)(0);
  CNStageIntLLRInputS1xD(146)(1) <= VNStageIntLLROutputS0xD(105)(1);
  CNStageIntLLRInputS1xD(197)(1) <= VNStageIntLLROutputS0xD(105)(2);
  CNStageIntLLRInputS1xD(237)(1) <= VNStageIntLLROutputS0xD(105)(3);
  CNStageIntLLRInputS1xD(300)(1) <= VNStageIntLLROutputS0xD(105)(4);
  CNStageIntLLRInputS1xD(338)(1) <= VNStageIntLLROutputS0xD(105)(5);
  CNStageIntLLRInputS1xD(12)(1) <= VNStageIntLLROutputS0xD(106)(0);
  CNStageIntLLRInputS1xD(157)(1) <= VNStageIntLLROutputS0xD(106)(1);
  CNStageIntLLRInputS1xD(223)(1) <= VNStageIntLLROutputS0xD(106)(2);
  CNStageIntLLRInputS1xD(272)(1) <= VNStageIntLLROutputS0xD(106)(3);
  CNStageIntLLRInputS1xD(312)(1) <= VNStageIntLLROutputS0xD(106)(4);
  CNStageIntLLRInputS1xD(333)(1) <= VNStageIntLLROutputS0xD(106)(5);
  CNStageIntLLRInputS1xD(110)(1) <= VNStageIntLLROutputS0xD(107)(0);
  CNStageIntLLRInputS1xD(127)(1) <= VNStageIntLLROutputS0xD(107)(1);
  CNStageIntLLRInputS1xD(207)(1) <= VNStageIntLLROutputS0xD(107)(2);
  CNStageIntLLRInputS1xD(230)(1) <= VNStageIntLLROutputS0xD(107)(3);
  CNStageIntLLRInputS1xD(323)(1) <= VNStageIntLLROutputS0xD(107)(4);
  CNStageIntLLRInputS1xD(335)(1) <= VNStageIntLLROutputS0xD(107)(5);
  CNStageIntLLRInputS1xD(11)(1) <= VNStageIntLLROutputS0xD(108)(0);
  CNStageIntLLRInputS1xD(105)(1) <= VNStageIntLLROutputS0xD(108)(1);
  CNStageIntLLRInputS1xD(115)(1) <= VNStageIntLLROutputS0xD(108)(2);
  CNStageIntLLRInputS1xD(181)(1) <= VNStageIntLLROutputS0xD(108)(3);
  CNStageIntLLRInputS1xD(238)(1) <= VNStageIntLLROutputS0xD(108)(4);
  CNStageIntLLRInputS1xD(296)(1) <= VNStageIntLLROutputS0xD(108)(5);
  CNStageIntLLRInputS1xD(10)(1) <= VNStageIntLLROutputS0xD(109)(0);
  CNStageIntLLRInputS1xD(100)(1) <= VNStageIntLLROutputS0xD(109)(1);
  CNStageIntLLRInputS1xD(160)(1) <= VNStageIntLLROutputS0xD(109)(2);
  CNStageIntLLRInputS1xD(171)(1) <= VNStageIntLLROutputS0xD(109)(3);
  CNStageIntLLRInputS1xD(266)(1) <= VNStageIntLLROutputS0xD(109)(4);
  CNStageIntLLRInputS1xD(362)(1) <= VNStageIntLLROutputS0xD(109)(5);
  CNStageIntLLRInputS1xD(9)(1) <= VNStageIntLLROutputS0xD(110)(0);
  CNStageIntLLRInputS1xD(83)(1) <= VNStageIntLLROutputS0xD(110)(1);
  CNStageIntLLRInputS1xD(118)(1) <= VNStageIntLLROutputS0xD(110)(2);
  CNStageIntLLRInputS1xD(212)(1) <= VNStageIntLLROutputS0xD(110)(3);
  CNStageIntLLRInputS1xD(225)(1) <= VNStageIntLLROutputS0xD(110)(4);
  CNStageIntLLRInputS1xD(326)(1) <= VNStageIntLLROutputS0xD(110)(5);
  CNStageIntLLRInputS1xD(345)(1) <= VNStageIntLLROutputS0xD(110)(6);
  CNStageIntLLRInputS1xD(8)(1) <= VNStageIntLLROutputS0xD(111)(0);
  CNStageIntLLRInputS1xD(90)(1) <= VNStageIntLLROutputS0xD(111)(1);
  CNStageIntLLRInputS1xD(138)(1) <= VNStageIntLLROutputS0xD(111)(2);
  CNStageIntLLRInputS1xD(177)(1) <= VNStageIntLLROutputS0xD(111)(3);
  CNStageIntLLRInputS1xD(252)(1) <= VNStageIntLLROutputS0xD(111)(4);
  CNStageIntLLRInputS1xD(287)(1) <= VNStageIntLLROutputS0xD(111)(5);
  CNStageIntLLRInputS1xD(357)(1) <= VNStageIntLLROutputS0xD(111)(6);
  CNStageIntLLRInputS1xD(7)(1) <= VNStageIntLLROutputS0xD(112)(0);
  CNStageIntLLRInputS1xD(54)(1) <= VNStageIntLLROutputS0xD(112)(1);
  CNStageIntLLRInputS1xD(148)(1) <= VNStageIntLLROutputS0xD(112)(2);
  CNStageIntLLRInputS1xD(205)(1) <= VNStageIntLLROutputS0xD(112)(3);
  CNStageIntLLRInputS1xD(233)(1) <= VNStageIntLLROutputS0xD(112)(4);
  CNStageIntLLRInputS1xD(305)(1) <= VNStageIntLLROutputS0xD(112)(5);
  CNStageIntLLRInputS1xD(369)(1) <= VNStageIntLLROutputS0xD(112)(6);
  CNStageIntLLRInputS1xD(6)(1) <= VNStageIntLLROutputS0xD(113)(0);
  CNStageIntLLRInputS1xD(108)(1) <= VNStageIntLLROutputS0xD(113)(1);
  CNStageIntLLRInputS1xD(143)(1) <= VNStageIntLLROutputS0xD(113)(2);
  CNStageIntLLRInputS1xD(202)(1) <= VNStageIntLLROutputS0xD(113)(3);
  CNStageIntLLRInputS1xD(253)(1) <= VNStageIntLLROutputS0xD(113)(4);
  CNStageIntLLRInputS1xD(314)(1) <= VNStageIntLLROutputS0xD(113)(5);
  CNStageIntLLRInputS1xD(339)(1) <= VNStageIntLLROutputS0xD(113)(6);
  CNStageIntLLRInputS1xD(5)(1) <= VNStageIntLLROutputS0xD(114)(0);
  CNStageIntLLRInputS1xD(88)(1) <= VNStageIntLLROutputS0xD(114)(1);
  CNStageIntLLRInputS1xD(149)(1) <= VNStageIntLLROutputS0xD(114)(2);
  CNStageIntLLRInputS1xD(216)(1) <= VNStageIntLLROutputS0xD(114)(3);
  CNStageIntLLRInputS1xD(268)(1) <= VNStageIntLLROutputS0xD(114)(4);
  CNStageIntLLRInputS1xD(309)(1) <= VNStageIntLLROutputS0xD(114)(5);
  CNStageIntLLRInputS1xD(4)(1) <= VNStageIntLLROutputS0xD(115)(0);
  CNStageIntLLRInputS1xD(68)(1) <= VNStageIntLLROutputS0xD(115)(1);
  CNStageIntLLRInputS1xD(137)(1) <= VNStageIntLLROutputS0xD(115)(2);
  CNStageIntLLRInputS1xD(209)(1) <= VNStageIntLLROutputS0xD(115)(3);
  CNStageIntLLRInputS1xD(264)(1) <= VNStageIntLLROutputS0xD(115)(4);
  CNStageIntLLRInputS1xD(315)(1) <= VNStageIntLLROutputS0xD(115)(5);
  CNStageIntLLRInputS1xD(372)(1) <= VNStageIntLLROutputS0xD(115)(6);
  CNStageIntLLRInputS1xD(71)(1) <= VNStageIntLLROutputS0xD(116)(0);
  CNStageIntLLRInputS1xD(163)(1) <= VNStageIntLLROutputS0xD(116)(1);
  CNStageIntLLRInputS1xD(187)(1) <= VNStageIntLLROutputS0xD(116)(2);
  CNStageIntLLRInputS1xD(228)(1) <= VNStageIntLLROutputS0xD(116)(3);
  CNStageIntLLRInputS1xD(304)(1) <= VNStageIntLLROutputS0xD(116)(4);
  CNStageIntLLRInputS1xD(3)(1) <= VNStageIntLLROutputS0xD(117)(0);
  CNStageIntLLRInputS1xD(55)(1) <= VNStageIntLLROutputS0xD(117)(1);
  CNStageIntLLRInputS1xD(111)(1) <= VNStageIntLLROutputS0xD(117)(2);
  CNStageIntLLRInputS1xD(196)(1) <= VNStageIntLLROutputS0xD(117)(3);
  CNStageIntLLRInputS1xD(2)(1) <= VNStageIntLLROutputS0xD(118)(0);
  CNStageIntLLRInputS1xD(89)(1) <= VNStageIntLLROutputS0xD(118)(1);
  CNStageIntLLRInputS1xD(152)(1) <= VNStageIntLLROutputS0xD(118)(2);
  CNStageIntLLRInputS1xD(249)(1) <= VNStageIntLLROutputS0xD(118)(3);
  CNStageIntLLRInputS1xD(282)(1) <= VNStageIntLLROutputS0xD(118)(4);
  CNStageIntLLRInputS1xD(359)(1) <= VNStageIntLLROutputS0xD(118)(5);
  CNStageIntLLRInputS1xD(1)(1) <= VNStageIntLLROutputS0xD(119)(0);
  CNStageIntLLRInputS1xD(107)(1) <= VNStageIntLLROutputS0xD(119)(1);
  CNStageIntLLRInputS1xD(154)(1) <= VNStageIntLLROutputS0xD(119)(2);
  CNStageIntLLRInputS1xD(227)(1) <= VNStageIntLLROutputS0xD(119)(3);
  CNStageIntLLRInputS1xD(319)(1) <= VNStageIntLLROutputS0xD(119)(4);
  CNStageIntLLRInputS1xD(0)(1) <= VNStageIntLLROutputS0xD(120)(0);
  CNStageIntLLRInputS1xD(80)(1) <= VNStageIntLLROutputS0xD(120)(1);
  CNStageIntLLRInputS1xD(321)(1) <= VNStageIntLLROutputS0xD(120)(2);
  CNStageIntLLRInputS1xD(360)(1) <= VNStageIntLLROutputS0xD(120)(3);
  CNStageIntLLRInputS1xD(64)(1) <= VNStageIntLLROutputS0xD(121)(0);
  CNStageIntLLRInputS1xD(161)(1) <= VNStageIntLLROutputS0xD(121)(1);
  CNStageIntLLRInputS1xD(217)(1) <= VNStageIntLLROutputS0xD(121)(2);
  CNStageIntLLRInputS1xD(236)(1) <= VNStageIntLLROutputS0xD(121)(3);
  CNStageIntLLRInputS1xD(291)(1) <= VNStageIntLLROutputS0xD(121)(4);
  CNStageIntLLRInputS1xD(350)(1) <= VNStageIntLLROutputS0xD(121)(5);
  CNStageIntLLRInputS1xD(91)(1) <= VNStageIntLLROutputS0xD(122)(0);
  CNStageIntLLRInputS1xD(114)(1) <= VNStageIntLLROutputS0xD(122)(1);
  CNStageIntLLRInputS1xD(201)(1) <= VNStageIntLLROutputS0xD(122)(2);
  CNStageIntLLRInputS1xD(241)(1) <= VNStageIntLLROutputS0xD(122)(3);
  CNStageIntLLRInputS1xD(327)(1) <= VNStageIntLLROutputS0xD(122)(4);
  CNStageIntLLRInputS1xD(375)(1) <= VNStageIntLLROutputS0xD(122)(5);
  CNStageIntLLRInputS1xD(82)(1) <= VNStageIntLLROutputS0xD(123)(0);
  CNStageIntLLRInputS1xD(122)(1) <= VNStageIntLLROutputS0xD(123)(1);
  CNStageIntLLRInputS1xD(213)(1) <= VNStageIntLLROutputS0xD(123)(2);
  CNStageIntLLRInputS1xD(279)(1) <= VNStageIntLLROutputS0xD(123)(3);
  CNStageIntLLRInputS1xD(382)(1) <= VNStageIntLLROutputS0xD(123)(4);
  CNStageIntLLRInputS1xD(69)(1) <= VNStageIntLLROutputS0xD(124)(0);
  CNStageIntLLRInputS1xD(153)(1) <= VNStageIntLLROutputS0xD(124)(1);
  CNStageIntLLRInputS1xD(240)(1) <= VNStageIntLLROutputS0xD(124)(2);
  CNStageIntLLRInputS1xD(292)(1) <= VNStageIntLLROutputS0xD(124)(3);
  CNStageIntLLRInputS1xD(364)(1) <= VNStageIntLLROutputS0xD(124)(4);
  CNStageIntLLRInputS1xD(87)(1) <= VNStageIntLLROutputS0xD(125)(0);
  CNStageIntLLRInputS1xD(169)(1) <= VNStageIntLLROutputS0xD(125)(1);
  CNStageIntLLRInputS1xD(320)(1) <= VNStageIntLLROutputS0xD(125)(2);
  CNStageIntLLRInputS1xD(366)(1) <= VNStageIntLLROutputS0xD(125)(3);
  CNStageIntLLRInputS1xD(60)(1) <= VNStageIntLLROutputS0xD(126)(0);
  CNStageIntLLRInputS1xD(139)(1) <= VNStageIntLLROutputS0xD(126)(1);
  CNStageIntLLRInputS1xD(186)(1) <= VNStageIntLLROutputS0xD(126)(2);
  CNStageIntLLRInputS1xD(271)(1) <= VNStageIntLLROutputS0xD(126)(3);
  CNStageIntLLRInputS1xD(281)(1) <= VNStageIntLLROutputS0xD(126)(4);
  CNStageIntLLRInputS1xD(334)(1) <= VNStageIntLLROutputS0xD(126)(5);
  CNStageIntLLRInputS1xD(52)(1) <= VNStageIntLLROutputS0xD(127)(0);
  CNStageIntLLRInputS1xD(57)(1) <= VNStageIntLLROutputS0xD(127)(1);
  CNStageIntLLRInputS1xD(117)(1) <= VNStageIntLLROutputS0xD(127)(2);
  CNStageIntLLRInputS1xD(173)(1) <= VNStageIntLLROutputS0xD(127)(3);
  CNStageIntLLRInputS1xD(277)(1) <= VNStageIntLLROutputS0xD(127)(4);
  CNStageIntLLRInputS1xD(306)(1) <= VNStageIntLLROutputS0xD(127)(5);
  CNStageIntLLRInputS1xD(373)(1) <= VNStageIntLLROutputS0xD(127)(6);
  CNStageIntLLRInputS1xD(53)(2) <= VNStageIntLLROutputS0xD(128)(0);
  CNStageIntLLRInputS1xD(108)(2) <= VNStageIntLLROutputS0xD(128)(1);
  CNStageIntLLRInputS1xD(129)(2) <= VNStageIntLLROutputS0xD(128)(2);
  CNStageIntLLRInputS1xD(198)(2) <= VNStageIntLLROutputS0xD(128)(3);
  CNStageIntLLRInputS1xD(244)(2) <= VNStageIntLLROutputS0xD(128)(4);
  CNStageIntLLRInputS1xD(298)(2) <= VNStageIntLLROutputS0xD(128)(5);
  CNStageIntLLRInputS1xD(341)(2) <= VNStageIntLLROutputS0xD(128)(6);
  CNStageIntLLRInputS1xD(51)(2) <= VNStageIntLLROutputS0xD(129)(0);
  CNStageIntLLRInputS1xD(56)(2) <= VNStageIntLLROutputS0xD(129)(1);
  CNStageIntLLRInputS1xD(116)(2) <= VNStageIntLLROutputS0xD(129)(2);
  CNStageIntLLRInputS1xD(172)(2) <= VNStageIntLLROutputS0xD(129)(3);
  CNStageIntLLRInputS1xD(276)(2) <= VNStageIntLLROutputS0xD(129)(4);
  CNStageIntLLRInputS1xD(305)(2) <= VNStageIntLLROutputS0xD(129)(5);
  CNStageIntLLRInputS1xD(372)(2) <= VNStageIntLLROutputS0xD(129)(6);
  CNStageIntLLRInputS1xD(50)(2) <= VNStageIntLLROutputS0xD(130)(0);
  CNStageIntLLRInputS1xD(73)(2) <= VNStageIntLLROutputS0xD(130)(1);
  CNStageIntLLRInputS1xD(140)(2) <= VNStageIntLLROutputS0xD(130)(2);
  CNStageIntLLRInputS1xD(188)(2) <= VNStageIntLLROutputS0xD(130)(3);
  CNStageIntLLRInputS1xD(245)(2) <= VNStageIntLLROutputS0xD(130)(4);
  CNStageIntLLRInputS1xD(285)(2) <= VNStageIntLLROutputS0xD(130)(5);
  CNStageIntLLRInputS1xD(65)(2) <= VNStageIntLLROutputS0xD(131)(0);
  CNStageIntLLRInputS1xD(154)(2) <= VNStageIntLLROutputS0xD(131)(1);
  CNStageIntLLRInputS1xD(206)(2) <= VNStageIntLLROutputS0xD(131)(2);
  CNStageIntLLRInputS1xD(243)(2) <= VNStageIntLLROutputS0xD(131)(3);
  CNStageIntLLRInputS1xD(307)(2) <= VNStageIntLLROutputS0xD(131)(4);
  CNStageIntLLRInputS1xD(334)(2) <= VNStageIntLLROutputS0xD(131)(5);
  CNStageIntLLRInputS1xD(49)(2) <= VNStageIntLLROutputS0xD(132)(0);
  CNStageIntLLRInputS1xD(151)(2) <= VNStageIntLLROutputS0xD(132)(1);
  CNStageIntLLRInputS1xD(214)(2) <= VNStageIntLLROutputS0xD(132)(2);
  CNStageIntLLRInputS1xD(274)(2) <= VNStageIntLLROutputS0xD(132)(3);
  CNStageIntLLRInputS1xD(321)(2) <= VNStageIntLLROutputS0xD(132)(4);
  CNStageIntLLRInputS1xD(364)(2) <= VNStageIntLLROutputS0xD(132)(5);
  CNStageIntLLRInputS1xD(48)(2) <= VNStageIntLLROutputS0xD(133)(0);
  CNStageIntLLRInputS1xD(209)(2) <= VNStageIntLLROutputS0xD(133)(1);
  CNStageIntLLRInputS1xD(255)(2) <= VNStageIntLLROutputS0xD(133)(2);
  CNStageIntLLRInputS1xD(317)(2) <= VNStageIntLLROutputS0xD(133)(3);
  CNStageIntLLRInputS1xD(380)(2) <= VNStageIntLLROutputS0xD(133)(4);
  CNStageIntLLRInputS1xD(47)(2) <= VNStageIntLLROutputS0xD(134)(0);
  CNStageIntLLRInputS1xD(100)(2) <= VNStageIntLLROutputS0xD(134)(1);
  CNStageIntLLRInputS1xD(134)(2) <= VNStageIntLLROutputS0xD(134)(2);
  CNStageIntLLRInputS1xD(258)(2) <= VNStageIntLLROutputS0xD(134)(3);
  CNStageIntLLRInputS1xD(46)(2) <= VNStageIntLLROutputS0xD(135)(0);
  CNStageIntLLRInputS1xD(103)(2) <= VNStageIntLLROutputS0xD(135)(1);
  CNStageIntLLRInputS1xD(135)(2) <= VNStageIntLLROutputS0xD(135)(2);
  CNStageIntLLRInputS1xD(205)(2) <= VNStageIntLLROutputS0xD(135)(3);
  CNStageIntLLRInputS1xD(45)(2) <= VNStageIntLLROutputS0xD(136)(0);
  CNStageIntLLRInputS1xD(94)(2) <= VNStageIntLLROutputS0xD(136)(1);
  CNStageIntLLRInputS1xD(111)(2) <= VNStageIntLLROutputS0xD(136)(2);
  CNStageIntLLRInputS1xD(175)(2) <= VNStageIntLLROutputS0xD(136)(3);
  CNStageIntLLRInputS1xD(275)(2) <= VNStageIntLLROutputS0xD(136)(4);
  CNStageIntLLRInputS1xD(301)(2) <= VNStageIntLLROutputS0xD(136)(5);
  CNStageIntLLRInputS1xD(352)(2) <= VNStageIntLLROutputS0xD(136)(6);
  CNStageIntLLRInputS1xD(44)(2) <= VNStageIntLLROutputS0xD(137)(0);
  CNStageIntLLRInputS1xD(74)(2) <= VNStageIntLLROutputS0xD(137)(1);
  CNStageIntLLRInputS1xD(161)(2) <= VNStageIntLLROutputS0xD(137)(2);
  CNStageIntLLRInputS1xD(182)(2) <= VNStageIntLLROutputS0xD(137)(3);
  CNStageIntLLRInputS1xD(242)(2) <= VNStageIntLLROutputS0xD(137)(4);
  CNStageIntLLRInputS1xD(282)(2) <= VNStageIntLLROutputS0xD(137)(5);
  CNStageIntLLRInputS1xD(366)(2) <= VNStageIntLLROutputS0xD(137)(6);
  CNStageIntLLRInputS1xD(43)(2) <= VNStageIntLLROutputS0xD(138)(0);
  CNStageIntLLRInputS1xD(55)(2) <= VNStageIntLLROutputS0xD(138)(1);
  CNStageIntLLRInputS1xD(120)(2) <= VNStageIntLLROutputS0xD(138)(2);
  CNStageIntLLRInputS1xD(218)(2) <= VNStageIntLLROutputS0xD(138)(3);
  CNStageIntLLRInputS1xD(268)(2) <= VNStageIntLLROutputS0xD(138)(4);
  CNStageIntLLRInputS1xD(327)(2) <= VNStageIntLLROutputS0xD(138)(5);
  CNStageIntLLRInputS1xD(362)(2) <= VNStageIntLLROutputS0xD(138)(6);
  CNStageIntLLRInputS1xD(42)(2) <= VNStageIntLLROutputS0xD(139)(0);
  CNStageIntLLRInputS1xD(69)(2) <= VNStageIntLLROutputS0xD(139)(1);
  CNStageIntLLRInputS1xD(124)(2) <= VNStageIntLLROutputS0xD(139)(2);
  CNStageIntLLRInputS1xD(220)(2) <= VNStageIntLLROutputS0xD(139)(3);
  CNStageIntLLRInputS1xD(252)(2) <= VNStageIntLLROutputS0xD(139)(4);
  CNStageIntLLRInputS1xD(289)(2) <= VNStageIntLLROutputS0xD(139)(5);
  CNStageIntLLRInputS1xD(383)(2) <= VNStageIntLLROutputS0xD(139)(6);
  CNStageIntLLRInputS1xD(41)(2) <= VNStageIntLLROutputS0xD(140)(0);
  CNStageIntLLRInputS1xD(80)(2) <= VNStageIntLLROutputS0xD(140)(1);
  CNStageIntLLRInputS1xD(170)(2) <= VNStageIntLLROutputS0xD(140)(2);
  CNStageIntLLRInputS1xD(191)(2) <= VNStageIntLLROutputS0xD(140)(3);
  CNStageIntLLRInputS1xD(277)(2) <= VNStageIntLLROutputS0xD(140)(4);
  CNStageIntLLRInputS1xD(293)(2) <= VNStageIntLLROutputS0xD(140)(5);
  CNStageIntLLRInputS1xD(346)(2) <= VNStageIntLLROutputS0xD(140)(6);
  CNStageIntLLRInputS1xD(123)(2) <= VNStageIntLLROutputS0xD(141)(0);
  CNStageIntLLRInputS1xD(173)(2) <= VNStageIntLLROutputS0xD(141)(1);
  CNStageIntLLRInputS1xD(269)(2) <= VNStageIntLLROutputS0xD(141)(2);
  CNStageIntLLRInputS1xD(332)(2) <= VNStageIntLLROutputS0xD(141)(3);
  CNStageIntLLRInputS1xD(347)(2) <= VNStageIntLLROutputS0xD(141)(4);
  CNStageIntLLRInputS1xD(40)(2) <= VNStageIntLLROutputS0xD(142)(0);
  CNStageIntLLRInputS1xD(96)(2) <= VNStageIntLLROutputS0xD(142)(1);
  CNStageIntLLRInputS1xD(118)(2) <= VNStageIntLLROutputS0xD(142)(2);
  CNStageIntLLRInputS1xD(256)(2) <= VNStageIntLLROutputS0xD(142)(3);
  CNStageIntLLRInputS1xD(382)(2) <= VNStageIntLLROutputS0xD(142)(4);
  CNStageIntLLRInputS1xD(39)(2) <= VNStageIntLLROutputS0xD(143)(0);
  CNStageIntLLRInputS1xD(83)(2) <= VNStageIntLLROutputS0xD(143)(1);
  CNStageIntLLRInputS1xD(158)(2) <= VNStageIntLLROutputS0xD(143)(2);
  CNStageIntLLRInputS1xD(192)(2) <= VNStageIntLLROutputS0xD(143)(3);
  CNStageIntLLRInputS1xD(273)(2) <= VNStageIntLLROutputS0xD(143)(4);
  CNStageIntLLRInputS1xD(287)(2) <= VNStageIntLLROutputS0xD(143)(5);
  CNStageIntLLRInputS1xD(373)(2) <= VNStageIntLLROutputS0xD(143)(6);
  CNStageIntLLRInputS1xD(38)(2) <= VNStageIntLLROutputS0xD(144)(0);
  CNStageIntLLRInputS1xD(98)(2) <= VNStageIntLLROutputS0xD(144)(1);
  CNStageIntLLRInputS1xD(166)(2) <= VNStageIntLLROutputS0xD(144)(2);
  CNStageIntLLRInputS1xD(219)(2) <= VNStageIntLLROutputS0xD(144)(3);
  CNStageIntLLRInputS1xD(249)(2) <= VNStageIntLLROutputS0xD(144)(4);
  CNStageIntLLRInputS1xD(324)(2) <= VNStageIntLLROutputS0xD(144)(5);
  CNStageIntLLRInputS1xD(333)(2) <= VNStageIntLLROutputS0xD(144)(6);
  CNStageIntLLRInputS1xD(37)(2) <= VNStageIntLLROutputS0xD(145)(0);
  CNStageIntLLRInputS1xD(61)(2) <= VNStageIntLLROutputS0xD(145)(1);
  CNStageIntLLRInputS1xD(130)(2) <= VNStageIntLLROutputS0xD(145)(2);
  CNStageIntLLRInputS1xD(181)(2) <= VNStageIntLLROutputS0xD(145)(3);
  CNStageIntLLRInputS1xD(247)(2) <= VNStageIntLLROutputS0xD(145)(4);
  CNStageIntLLRInputS1xD(331)(2) <= VNStageIntLLROutputS0xD(145)(5);
  CNStageIntLLRInputS1xD(336)(2) <= VNStageIntLLROutputS0xD(145)(6);
  CNStageIntLLRInputS1xD(36)(2) <= VNStageIntLLROutputS0xD(146)(0);
  CNStageIntLLRInputS1xD(71)(2) <= VNStageIntLLROutputS0xD(146)(1);
  CNStageIntLLRInputS1xD(128)(2) <= VNStageIntLLROutputS0xD(146)(2);
  CNStageIntLLRInputS1xD(261)(2) <= VNStageIntLLROutputS0xD(146)(3);
  CNStageIntLLRInputS1xD(299)(2) <= VNStageIntLLROutputS0xD(146)(4);
  CNStageIntLLRInputS1xD(35)(2) <= VNStageIntLLROutputS0xD(147)(0);
  CNStageIntLLRInputS1xD(66)(2) <= VNStageIntLLROutputS0xD(147)(1);
  CNStageIntLLRInputS1xD(164)(2) <= VNStageIntLLROutputS0xD(147)(2);
  CNStageIntLLRInputS1xD(187)(2) <= VNStageIntLLROutputS0xD(147)(3);
  CNStageIntLLRInputS1xD(253)(2) <= VNStageIntLLROutputS0xD(147)(4);
  CNStageIntLLRInputS1xD(297)(2) <= VNStageIntLLROutputS0xD(147)(5);
  CNStageIntLLRInputS1xD(335)(2) <= VNStageIntLLROutputS0xD(147)(6);
  CNStageIntLLRInputS1xD(34)(2) <= VNStageIntLLROutputS0xD(148)(0);
  CNStageIntLLRInputS1xD(72)(2) <= VNStageIntLLROutputS0xD(148)(1);
  CNStageIntLLRInputS1xD(143)(2) <= VNStageIntLLROutputS0xD(148)(2);
  CNStageIntLLRInputS1xD(207)(2) <= VNStageIntLLROutputS0xD(148)(3);
  CNStageIntLLRInputS1xD(231)(2) <= VNStageIntLLROutputS0xD(148)(4);
  CNStageIntLLRInputS1xD(329)(2) <= VNStageIntLLROutputS0xD(148)(5);
  CNStageIntLLRInputS1xD(33)(2) <= VNStageIntLLROutputS0xD(149)(0);
  CNStageIntLLRInputS1xD(60)(2) <= VNStageIntLLROutputS0xD(149)(1);
  CNStageIntLLRInputS1xD(146)(2) <= VNStageIntLLROutputS0xD(149)(2);
  CNStageIntLLRInputS1xD(221)(2) <= VNStageIntLLROutputS0xD(149)(3);
  CNStageIntLLRInputS1xD(241)(2) <= VNStageIntLLROutputS0xD(149)(4);
  CNStageIntLLRInputS1xD(309)(2) <= VNStageIntLLROutputS0xD(149)(5);
  CNStageIntLLRInputS1xD(370)(2) <= VNStageIntLLROutputS0xD(149)(6);
  CNStageIntLLRInputS1xD(32)(2) <= VNStageIntLLROutputS0xD(150)(0);
  CNStageIntLLRInputS1xD(86)(2) <= VNStageIntLLROutputS0xD(150)(1);
  CNStageIntLLRInputS1xD(131)(2) <= VNStageIntLLROutputS0xD(150)(2);
  CNStageIntLLRInputS1xD(217)(2) <= VNStageIntLLROutputS0xD(150)(3);
  CNStageIntLLRInputS1xD(312)(2) <= VNStageIntLLROutputS0xD(150)(4);
  CNStageIntLLRInputS1xD(378)(2) <= VNStageIntLLROutputS0xD(150)(5);
  CNStageIntLLRInputS1xD(31)(2) <= VNStageIntLLROutputS0xD(151)(0);
  CNStageIntLLRInputS1xD(92)(2) <= VNStageIntLLROutputS0xD(151)(1);
  CNStageIntLLRInputS1xD(165)(2) <= VNStageIntLLROutputS0xD(151)(2);
  CNStageIntLLRInputS1xD(184)(2) <= VNStageIntLLROutputS0xD(151)(3);
  CNStageIntLLRInputS1xD(238)(2) <= VNStageIntLLROutputS0xD(151)(4);
  CNStageIntLLRInputS1xD(342)(2) <= VNStageIntLLROutputS0xD(151)(5);
  CNStageIntLLRInputS1xD(30)(2) <= VNStageIntLLROutputS0xD(152)(0);
  CNStageIntLLRInputS1xD(76)(2) <= VNStageIntLLROutputS0xD(152)(1);
  CNStageIntLLRInputS1xD(127)(2) <= VNStageIntLLROutputS0xD(152)(2);
  CNStageIntLLRInputS1xD(202)(2) <= VNStageIntLLROutputS0xD(152)(3);
  CNStageIntLLRInputS1xD(228)(2) <= VNStageIntLLROutputS0xD(152)(4);
  CNStageIntLLRInputS1xD(330)(2) <= VNStageIntLLROutputS0xD(152)(5);
  CNStageIntLLRInputS1xD(340)(2) <= VNStageIntLLROutputS0xD(152)(6);
  CNStageIntLLRInputS1xD(29)(2) <= VNStageIntLLROutputS0xD(153)(0);
  CNStageIntLLRInputS1xD(78)(2) <= VNStageIntLLROutputS0xD(153)(1);
  CNStageIntLLRInputS1xD(155)(2) <= VNStageIntLLROutputS0xD(153)(2);
  CNStageIntLLRInputS1xD(203)(2) <= VNStageIntLLROutputS0xD(153)(3);
  CNStageIntLLRInputS1xD(262)(2) <= VNStageIntLLROutputS0xD(153)(4);
  CNStageIntLLRInputS1xD(296)(2) <= VNStageIntLLROutputS0xD(153)(5);
  CNStageIntLLRInputS1xD(376)(2) <= VNStageIntLLROutputS0xD(153)(6);
  CNStageIntLLRInputS1xD(28)(2) <= VNStageIntLLROutputS0xD(154)(0);
  CNStageIntLLRInputS1xD(139)(2) <= VNStageIntLLROutputS0xD(154)(1);
  CNStageIntLLRInputS1xD(183)(2) <= VNStageIntLLROutputS0xD(154)(2);
  CNStageIntLLRInputS1xD(246)(2) <= VNStageIntLLROutputS0xD(154)(3);
  CNStageIntLLRInputS1xD(322)(2) <= VNStageIntLLROutputS0xD(154)(4);
  CNStageIntLLRInputS1xD(27)(2) <= VNStageIntLLROutputS0xD(155)(0);
  CNStageIntLLRInputS1xD(84)(2) <= VNStageIntLLROutputS0xD(155)(1);
  CNStageIntLLRInputS1xD(167)(2) <= VNStageIntLLROutputS0xD(155)(2);
  CNStageIntLLRInputS1xD(174)(2) <= VNStageIntLLROutputS0xD(155)(3);
  CNStageIntLLRInputS1xD(257)(2) <= VNStageIntLLROutputS0xD(155)(4);
  CNStageIntLLRInputS1xD(306)(2) <= VNStageIntLLROutputS0xD(155)(5);
  CNStageIntLLRInputS1xD(357)(2) <= VNStageIntLLROutputS0xD(155)(6);
  CNStageIntLLRInputS1xD(26)(2) <= VNStageIntLLROutputS0xD(156)(0);
  CNStageIntLLRInputS1xD(95)(2) <= VNStageIntLLROutputS0xD(156)(1);
  CNStageIntLLRInputS1xD(157)(2) <= VNStageIntLLROutputS0xD(156)(2);
  CNStageIntLLRInputS1xD(343)(2) <= VNStageIntLLROutputS0xD(156)(3);
  CNStageIntLLRInputS1xD(25)(2) <= VNStageIntLLROutputS0xD(157)(0);
  CNStageIntLLRInputS1xD(102)(2) <= VNStageIntLLROutputS0xD(157)(1);
  CNStageIntLLRInputS1xD(144)(2) <= VNStageIntLLROutputS0xD(157)(2);
  CNStageIntLLRInputS1xD(194)(2) <= VNStageIntLLROutputS0xD(157)(3);
  CNStageIntLLRInputS1xD(323)(2) <= VNStageIntLLROutputS0xD(157)(4);
  CNStageIntLLRInputS1xD(377)(2) <= VNStageIntLLROutputS0xD(157)(5);
  CNStageIntLLRInputS1xD(24)(2) <= VNStageIntLLROutputS0xD(158)(0);
  CNStageIntLLRInputS1xD(77)(2) <= VNStageIntLLROutputS0xD(158)(1);
  CNStageIntLLRInputS1xD(163)(2) <= VNStageIntLLROutputS0xD(158)(2);
  CNStageIntLLRInputS1xD(224)(2) <= VNStageIntLLROutputS0xD(158)(3);
  CNStageIntLLRInputS1xD(230)(2) <= VNStageIntLLROutputS0xD(158)(4);
  CNStageIntLLRInputS1xD(310)(2) <= VNStageIntLLROutputS0xD(158)(5);
  CNStageIntLLRInputS1xD(339)(2) <= VNStageIntLLROutputS0xD(158)(6);
  CNStageIntLLRInputS1xD(23)(2) <= VNStageIntLLROutputS0xD(159)(0);
  CNStageIntLLRInputS1xD(91)(2) <= VNStageIntLLROutputS0xD(159)(1);
  CNStageIntLLRInputS1xD(136)(2) <= VNStageIntLLROutputS0xD(159)(2);
  CNStageIntLLRInputS1xD(271)(2) <= VNStageIntLLROutputS0xD(159)(3);
  CNStageIntLLRInputS1xD(367)(2) <= VNStageIntLLROutputS0xD(159)(4);
  CNStageIntLLRInputS1xD(22)(2) <= VNStageIntLLROutputS0xD(160)(0);
  CNStageIntLLRInputS1xD(62)(2) <= VNStageIntLLROutputS0xD(160)(1);
  CNStageIntLLRInputS1xD(133)(2) <= VNStageIntLLROutputS0xD(160)(2);
  CNStageIntLLRInputS1xD(189)(2) <= VNStageIntLLROutputS0xD(160)(3);
  CNStageIntLLRInputS1xD(233)(2) <= VNStageIntLLROutputS0xD(160)(4);
  CNStageIntLLRInputS1xD(302)(2) <= VNStageIntLLROutputS0xD(160)(5);
  CNStageIntLLRInputS1xD(351)(2) <= VNStageIntLLROutputS0xD(160)(6);
  CNStageIntLLRInputS1xD(21)(2) <= VNStageIntLLROutputS0xD(161)(0);
  CNStageIntLLRInputS1xD(97)(2) <= VNStageIntLLROutputS0xD(161)(1);
  CNStageIntLLRInputS1xD(149)(2) <= VNStageIntLLROutputS0xD(161)(2);
  CNStageIntLLRInputS1xD(171)(2) <= VNStageIntLLROutputS0xD(161)(3);
  CNStageIntLLRInputS1xD(250)(2) <= VNStageIntLLROutputS0xD(161)(4);
  CNStageIntLLRInputS1xD(300)(2) <= VNStageIntLLROutputS0xD(161)(5);
  CNStageIntLLRInputS1xD(379)(2) <= VNStageIntLLROutputS0xD(161)(6);
  CNStageIntLLRInputS1xD(20)(2) <= VNStageIntLLROutputS0xD(162)(0);
  CNStageIntLLRInputS1xD(64)(2) <= VNStageIntLLROutputS0xD(162)(1);
  CNStageIntLLRInputS1xD(141)(2) <= VNStageIntLLROutputS0xD(162)(2);
  CNStageIntLLRInputS1xD(179)(2) <= VNStageIntLLROutputS0xD(162)(3);
  CNStageIntLLRInputS1xD(259)(2) <= VNStageIntLLROutputS0xD(162)(4);
  CNStageIntLLRInputS1xD(315)(2) <= VNStageIntLLROutputS0xD(162)(5);
  CNStageIntLLRInputS1xD(369)(2) <= VNStageIntLLROutputS0xD(162)(6);
  CNStageIntLLRInputS1xD(19)(2) <= VNStageIntLLROutputS0xD(163)(0);
  CNStageIntLLRInputS1xD(79)(2) <= VNStageIntLLROutputS0xD(163)(1);
  CNStageIntLLRInputS1xD(115)(2) <= VNStageIntLLROutputS0xD(163)(2);
  CNStageIntLLRInputS1xD(254)(2) <= VNStageIntLLROutputS0xD(163)(3);
  CNStageIntLLRInputS1xD(355)(2) <= VNStageIntLLROutputS0xD(163)(4);
  CNStageIntLLRInputS1xD(18)(2) <= VNStageIntLLROutputS0xD(164)(0);
  CNStageIntLLRInputS1xD(75)(2) <= VNStageIntLLROutputS0xD(164)(1);
  CNStageIntLLRInputS1xD(125)(2) <= VNStageIntLLROutputS0xD(164)(2);
  CNStageIntLLRInputS1xD(197)(2) <= VNStageIntLLROutputS0xD(164)(3);
  CNStageIntLLRInputS1xD(260)(2) <= VNStageIntLLROutputS0xD(164)(4);
  CNStageIntLLRInputS1xD(375)(2) <= VNStageIntLLROutputS0xD(164)(5);
  CNStageIntLLRInputS1xD(17)(2) <= VNStageIntLLROutputS0xD(165)(0);
  CNStageIntLLRInputS1xD(93)(2) <= VNStageIntLLROutputS0xD(165)(1);
  CNStageIntLLRInputS1xD(119)(2) <= VNStageIntLLROutputS0xD(165)(2);
  CNStageIntLLRInputS1xD(177)(2) <= VNStageIntLLROutputS0xD(165)(3);
  CNStageIntLLRInputS1xD(294)(2) <= VNStageIntLLROutputS0xD(165)(4);
  CNStageIntLLRInputS1xD(348)(2) <= VNStageIntLLROutputS0xD(165)(5);
  CNStageIntLLRInputS1xD(16)(2) <= VNStageIntLLROutputS0xD(166)(0);
  CNStageIntLLRInputS1xD(57)(2) <= VNStageIntLLROutputS0xD(166)(1);
  CNStageIntLLRInputS1xD(122)(2) <= VNStageIntLLROutputS0xD(166)(2);
  CNStageIntLLRInputS1xD(210)(2) <= VNStageIntLLROutputS0xD(166)(3);
  CNStageIntLLRInputS1xD(288)(2) <= VNStageIntLLROutputS0xD(166)(4);
  CNStageIntLLRInputS1xD(345)(2) <= VNStageIntLLROutputS0xD(166)(5);
  CNStageIntLLRInputS1xD(15)(2) <= VNStageIntLLROutputS0xD(167)(0);
  CNStageIntLLRInputS1xD(58)(2) <= VNStageIntLLROutputS0xD(167)(1);
  CNStageIntLLRInputS1xD(112)(2) <= VNStageIntLLROutputS0xD(167)(2);
  CNStageIntLLRInputS1xD(213)(2) <= VNStageIntLLROutputS0xD(167)(3);
  CNStageIntLLRInputS1xD(225)(2) <= VNStageIntLLROutputS0xD(167)(4);
  CNStageIntLLRInputS1xD(292)(2) <= VNStageIntLLROutputS0xD(167)(5);
  CNStageIntLLRInputS1xD(360)(2) <= VNStageIntLLROutputS0xD(167)(6);
  CNStageIntLLRInputS1xD(14)(2) <= VNStageIntLLROutputS0xD(168)(0);
  CNStageIntLLRInputS1xD(150)(2) <= VNStageIntLLROutputS0xD(168)(1);
  CNStageIntLLRInputS1xD(199)(2) <= VNStageIntLLROutputS0xD(168)(2);
  CNStageIntLLRInputS1xD(264)(2) <= VNStageIntLLROutputS0xD(168)(3);
  CNStageIntLLRInputS1xD(283)(2) <= VNStageIntLLROutputS0xD(168)(4);
  CNStageIntLLRInputS1xD(353)(2) <= VNStageIntLLROutputS0xD(168)(5);
  CNStageIntLLRInputS1xD(13)(2) <= VNStageIntLLROutputS0xD(169)(0);
  CNStageIntLLRInputS1xD(85)(2) <= VNStageIntLLROutputS0xD(169)(1);
  CNStageIntLLRInputS1xD(132)(2) <= VNStageIntLLROutputS0xD(169)(2);
  CNStageIntLLRInputS1xD(178)(2) <= VNStageIntLLROutputS0xD(169)(3);
  CNStageIntLLRInputS1xD(266)(2) <= VNStageIntLLROutputS0xD(169)(4);
  CNStageIntLLRInputS1xD(316)(2) <= VNStageIntLLROutputS0xD(169)(5);
  CNStageIntLLRInputS1xD(12)(2) <= VNStageIntLLROutputS0xD(170)(0);
  CNStageIntLLRInputS1xD(101)(2) <= VNStageIntLLROutputS0xD(170)(1);
  CNStageIntLLRInputS1xD(145)(2) <= VNStageIntLLROutputS0xD(170)(2);
  CNStageIntLLRInputS1xD(236)(2) <= VNStageIntLLROutputS0xD(170)(3);
  CNStageIntLLRInputS1xD(337)(2) <= VNStageIntLLROutputS0xD(170)(4);
  CNStageIntLLRInputS1xD(105)(2) <= VNStageIntLLROutputS0xD(171)(0);
  CNStageIntLLRInputS1xD(156)(2) <= VNStageIntLLROutputS0xD(171)(1);
  CNStageIntLLRInputS1xD(222)(2) <= VNStageIntLLROutputS0xD(171)(2);
  CNStageIntLLRInputS1xD(311)(2) <= VNStageIntLLROutputS0xD(171)(3);
  CNStageIntLLRInputS1xD(11)(2) <= VNStageIntLLROutputS0xD(172)(0);
  CNStageIntLLRInputS1xD(110)(2) <= VNStageIntLLROutputS0xD(172)(1);
  CNStageIntLLRInputS1xD(126)(2) <= VNStageIntLLROutputS0xD(172)(2);
  CNStageIntLLRInputS1xD(229)(2) <= VNStageIntLLROutputS0xD(172)(3);
  CNStageIntLLRInputS1xD(10)(2) <= VNStageIntLLROutputS0xD(173)(0);
  CNStageIntLLRInputS1xD(104)(2) <= VNStageIntLLROutputS0xD(173)(1);
  CNStageIntLLRInputS1xD(114)(2) <= VNStageIntLLROutputS0xD(173)(2);
  CNStageIntLLRInputS1xD(180)(2) <= VNStageIntLLROutputS0xD(173)(3);
  CNStageIntLLRInputS1xD(237)(2) <= VNStageIntLLROutputS0xD(173)(4);
  CNStageIntLLRInputS1xD(295)(2) <= VNStageIntLLROutputS0xD(173)(5);
  CNStageIntLLRInputS1xD(9)(2) <= VNStageIntLLROutputS0xD(174)(0);
  CNStageIntLLRInputS1xD(99)(2) <= VNStageIntLLROutputS0xD(174)(1);
  CNStageIntLLRInputS1xD(159)(2) <= VNStageIntLLROutputS0xD(174)(2);
  CNStageIntLLRInputS1xD(265)(2) <= VNStageIntLLROutputS0xD(174)(3);
  CNStageIntLLRInputS1xD(361)(2) <= VNStageIntLLROutputS0xD(174)(4);
  CNStageIntLLRInputS1xD(8)(2) <= VNStageIntLLROutputS0xD(175)(0);
  CNStageIntLLRInputS1xD(82)(2) <= VNStageIntLLROutputS0xD(175)(1);
  CNStageIntLLRInputS1xD(117)(2) <= VNStageIntLLROutputS0xD(175)(2);
  CNStageIntLLRInputS1xD(211)(2) <= VNStageIntLLROutputS0xD(175)(3);
  CNStageIntLLRInputS1xD(278)(2) <= VNStageIntLLROutputS0xD(175)(4);
  CNStageIntLLRInputS1xD(325)(2) <= VNStageIntLLROutputS0xD(175)(5);
  CNStageIntLLRInputS1xD(344)(2) <= VNStageIntLLROutputS0xD(175)(6);
  CNStageIntLLRInputS1xD(7)(2) <= VNStageIntLLROutputS0xD(176)(0);
  CNStageIntLLRInputS1xD(89)(2) <= VNStageIntLLROutputS0xD(176)(1);
  CNStageIntLLRInputS1xD(137)(2) <= VNStageIntLLROutputS0xD(176)(2);
  CNStageIntLLRInputS1xD(176)(2) <= VNStageIntLLROutputS0xD(176)(3);
  CNStageIntLLRInputS1xD(251)(2) <= VNStageIntLLROutputS0xD(176)(4);
  CNStageIntLLRInputS1xD(286)(2) <= VNStageIntLLROutputS0xD(176)(5);
  CNStageIntLLRInputS1xD(356)(2) <= VNStageIntLLROutputS0xD(176)(6);
  CNStageIntLLRInputS1xD(6)(2) <= VNStageIntLLROutputS0xD(177)(0);
  CNStageIntLLRInputS1xD(109)(2) <= VNStageIntLLROutputS0xD(177)(1);
  CNStageIntLLRInputS1xD(147)(2) <= VNStageIntLLROutputS0xD(177)(2);
  CNStageIntLLRInputS1xD(204)(2) <= VNStageIntLLROutputS0xD(177)(3);
  CNStageIntLLRInputS1xD(232)(2) <= VNStageIntLLROutputS0xD(177)(4);
  CNStageIntLLRInputS1xD(304)(2) <= VNStageIntLLROutputS0xD(177)(5);
  CNStageIntLLRInputS1xD(368)(2) <= VNStageIntLLROutputS0xD(177)(6);
  CNStageIntLLRInputS1xD(5)(2) <= VNStageIntLLROutputS0xD(178)(0);
  CNStageIntLLRInputS1xD(107)(2) <= VNStageIntLLROutputS0xD(178)(1);
  CNStageIntLLRInputS1xD(142)(2) <= VNStageIntLLROutputS0xD(178)(2);
  CNStageIntLLRInputS1xD(201)(2) <= VNStageIntLLROutputS0xD(178)(3);
  CNStageIntLLRInputS1xD(313)(2) <= VNStageIntLLROutputS0xD(178)(4);
  CNStageIntLLRInputS1xD(338)(2) <= VNStageIntLLROutputS0xD(178)(5);
  CNStageIntLLRInputS1xD(4)(2) <= VNStageIntLLROutputS0xD(179)(0);
  CNStageIntLLRInputS1xD(87)(2) <= VNStageIntLLROutputS0xD(179)(1);
  CNStageIntLLRInputS1xD(148)(2) <= VNStageIntLLROutputS0xD(179)(2);
  CNStageIntLLRInputS1xD(215)(2) <= VNStageIntLLROutputS0xD(179)(3);
  CNStageIntLLRInputS1xD(267)(2) <= VNStageIntLLROutputS0xD(179)(4);
  CNStageIntLLRInputS1xD(308)(2) <= VNStageIntLLROutputS0xD(179)(5);
  CNStageIntLLRInputS1xD(67)(2) <= VNStageIntLLROutputS0xD(180)(0);
  CNStageIntLLRInputS1xD(208)(2) <= VNStageIntLLROutputS0xD(180)(1);
  CNStageIntLLRInputS1xD(263)(2) <= VNStageIntLLROutputS0xD(180)(2);
  CNStageIntLLRInputS1xD(314)(2) <= VNStageIntLLROutputS0xD(180)(3);
  CNStageIntLLRInputS1xD(371)(2) <= VNStageIntLLROutputS0xD(180)(4);
  CNStageIntLLRInputS1xD(3)(2) <= VNStageIntLLROutputS0xD(181)(0);
  CNStageIntLLRInputS1xD(70)(2) <= VNStageIntLLROutputS0xD(181)(1);
  CNStageIntLLRInputS1xD(162)(2) <= VNStageIntLLROutputS0xD(181)(2);
  CNStageIntLLRInputS1xD(186)(2) <= VNStageIntLLROutputS0xD(181)(3);
  CNStageIntLLRInputS1xD(227)(2) <= VNStageIntLLROutputS0xD(181)(4);
  CNStageIntLLRInputS1xD(303)(2) <= VNStageIntLLROutputS0xD(181)(5);
  CNStageIntLLRInputS1xD(2)(2) <= VNStageIntLLROutputS0xD(182)(0);
  CNStageIntLLRInputS1xD(54)(2) <= VNStageIntLLROutputS0xD(182)(1);
  CNStageIntLLRInputS1xD(169)(2) <= VNStageIntLLROutputS0xD(182)(2);
  CNStageIntLLRInputS1xD(195)(2) <= VNStageIntLLROutputS0xD(182)(3);
  CNStageIntLLRInputS1xD(248)(2) <= VNStageIntLLROutputS0xD(182)(4);
  CNStageIntLLRInputS1xD(328)(2) <= VNStageIntLLROutputS0xD(182)(5);
  CNStageIntLLRInputS1xD(350)(2) <= VNStageIntLLROutputS0xD(182)(6);
  CNStageIntLLRInputS1xD(1)(2) <= VNStageIntLLROutputS0xD(183)(0);
  CNStageIntLLRInputS1xD(88)(2) <= VNStageIntLLROutputS0xD(183)(1);
  CNStageIntLLRInputS1xD(190)(2) <= VNStageIntLLROutputS0xD(183)(2);
  CNStageIntLLRInputS1xD(281)(2) <= VNStageIntLLROutputS0xD(183)(3);
  CNStageIntLLRInputS1xD(358)(2) <= VNStageIntLLROutputS0xD(183)(4);
  CNStageIntLLRInputS1xD(0)(2) <= VNStageIntLLROutputS0xD(184)(0);
  CNStageIntLLRInputS1xD(106)(2) <= VNStageIntLLROutputS0xD(184)(1);
  CNStageIntLLRInputS1xD(153)(2) <= VNStageIntLLROutputS0xD(184)(2);
  CNStageIntLLRInputS1xD(193)(2) <= VNStageIntLLROutputS0xD(184)(3);
  CNStageIntLLRInputS1xD(226)(2) <= VNStageIntLLROutputS0xD(184)(4);
  CNStageIntLLRInputS1xD(318)(2) <= VNStageIntLLROutputS0xD(184)(5);
  CNStageIntLLRInputS1xD(354)(2) <= VNStageIntLLROutputS0xD(184)(6);
  CNStageIntLLRInputS1xD(121)(2) <= VNStageIntLLROutputS0xD(185)(0);
  CNStageIntLLRInputS1xD(272)(2) <= VNStageIntLLROutputS0xD(185)(1);
  CNStageIntLLRInputS1xD(320)(2) <= VNStageIntLLROutputS0xD(185)(2);
  CNStageIntLLRInputS1xD(359)(2) <= VNStageIntLLROutputS0xD(185)(3);
  CNStageIntLLRInputS1xD(63)(2) <= VNStageIntLLROutputS0xD(186)(0);
  CNStageIntLLRInputS1xD(160)(2) <= VNStageIntLLROutputS0xD(186)(1);
  CNStageIntLLRInputS1xD(216)(2) <= VNStageIntLLROutputS0xD(186)(2);
  CNStageIntLLRInputS1xD(235)(2) <= VNStageIntLLROutputS0xD(186)(3);
  CNStageIntLLRInputS1xD(290)(2) <= VNStageIntLLROutputS0xD(186)(4);
  CNStageIntLLRInputS1xD(349)(2) <= VNStageIntLLROutputS0xD(186)(5);
  CNStageIntLLRInputS1xD(90)(2) <= VNStageIntLLROutputS0xD(187)(0);
  CNStageIntLLRInputS1xD(113)(2) <= VNStageIntLLROutputS0xD(187)(1);
  CNStageIntLLRInputS1xD(200)(2) <= VNStageIntLLROutputS0xD(187)(2);
  CNStageIntLLRInputS1xD(240)(2) <= VNStageIntLLROutputS0xD(187)(3);
  CNStageIntLLRInputS1xD(326)(2) <= VNStageIntLLROutputS0xD(187)(4);
  CNStageIntLLRInputS1xD(374)(2) <= VNStageIntLLROutputS0xD(187)(5);
  CNStageIntLLRInputS1xD(81)(2) <= VNStageIntLLROutputS0xD(188)(0);
  CNStageIntLLRInputS1xD(212)(2) <= VNStageIntLLROutputS0xD(188)(1);
  CNStageIntLLRInputS1xD(279)(2) <= VNStageIntLLROutputS0xD(188)(2);
  CNStageIntLLRInputS1xD(284)(2) <= VNStageIntLLROutputS0xD(188)(3);
  CNStageIntLLRInputS1xD(381)(2) <= VNStageIntLLROutputS0xD(188)(4);
  CNStageIntLLRInputS1xD(68)(2) <= VNStageIntLLROutputS0xD(189)(0);
  CNStageIntLLRInputS1xD(152)(2) <= VNStageIntLLROutputS0xD(189)(1);
  CNStageIntLLRInputS1xD(223)(2) <= VNStageIntLLROutputS0xD(189)(2);
  CNStageIntLLRInputS1xD(239)(2) <= VNStageIntLLROutputS0xD(189)(3);
  CNStageIntLLRInputS1xD(291)(2) <= VNStageIntLLROutputS0xD(189)(4);
  CNStageIntLLRInputS1xD(363)(2) <= VNStageIntLLROutputS0xD(189)(5);
  CNStageIntLLRInputS1xD(168)(2) <= VNStageIntLLROutputS0xD(190)(0);
  CNStageIntLLRInputS1xD(196)(2) <= VNStageIntLLROutputS0xD(190)(1);
  CNStageIntLLRInputS1xD(234)(2) <= VNStageIntLLROutputS0xD(190)(2);
  CNStageIntLLRInputS1xD(319)(2) <= VNStageIntLLROutputS0xD(190)(3);
  CNStageIntLLRInputS1xD(365)(2) <= VNStageIntLLROutputS0xD(190)(4);
  CNStageIntLLRInputS1xD(52)(2) <= VNStageIntLLROutputS0xD(191)(0);
  CNStageIntLLRInputS1xD(59)(2) <= VNStageIntLLROutputS0xD(191)(1);
  CNStageIntLLRInputS1xD(138)(2) <= VNStageIntLLROutputS0xD(191)(2);
  CNStageIntLLRInputS1xD(185)(2) <= VNStageIntLLROutputS0xD(191)(3);
  CNStageIntLLRInputS1xD(270)(2) <= VNStageIntLLROutputS0xD(191)(4);
  CNStageIntLLRInputS1xD(280)(2) <= VNStageIntLLROutputS0xD(191)(5);
  CNStageIntLLRInputS1xD(53)(3) <= VNStageIntLLROutputS0xD(192)(0);
  CNStageIntLLRInputS1xD(107)(3) <= VNStageIntLLROutputS0xD(192)(1);
  CNStageIntLLRInputS1xD(128)(3) <= VNStageIntLLROutputS0xD(192)(2);
  CNStageIntLLRInputS1xD(197)(3) <= VNStageIntLLROutputS0xD(192)(3);
  CNStageIntLLRInputS1xD(243)(3) <= VNStageIntLLROutputS0xD(192)(4);
  CNStageIntLLRInputS1xD(297)(3) <= VNStageIntLLROutputS0xD(192)(5);
  CNStageIntLLRInputS1xD(340)(3) <= VNStageIntLLROutputS0xD(192)(6);
  CNStageIntLLRInputS1xD(51)(3) <= VNStageIntLLROutputS0xD(193)(0);
  CNStageIntLLRInputS1xD(58)(3) <= VNStageIntLLROutputS0xD(193)(1);
  CNStageIntLLRInputS1xD(137)(3) <= VNStageIntLLROutputS0xD(193)(2);
  CNStageIntLLRInputS1xD(269)(3) <= VNStageIntLLROutputS0xD(193)(3);
  CNStageIntLLRInputS1xD(333)(3) <= VNStageIntLLROutputS0xD(193)(4);
  CNStageIntLLRInputS1xD(50)(3) <= VNStageIntLLROutputS0xD(194)(0);
  CNStageIntLLRInputS1xD(55)(3) <= VNStageIntLLROutputS0xD(194)(1);
  CNStageIntLLRInputS1xD(115)(3) <= VNStageIntLLROutputS0xD(194)(2);
  CNStageIntLLRInputS1xD(171)(3) <= VNStageIntLLROutputS0xD(194)(3);
  CNStageIntLLRInputS1xD(275)(3) <= VNStageIntLLROutputS0xD(194)(4);
  CNStageIntLLRInputS1xD(304)(3) <= VNStageIntLLROutputS0xD(194)(5);
  CNStageIntLLRInputS1xD(371)(3) <= VNStageIntLLROutputS0xD(194)(6);
  CNStageIntLLRInputS1xD(72)(3) <= VNStageIntLLROutputS0xD(195)(0);
  CNStageIntLLRInputS1xD(139)(3) <= VNStageIntLLROutputS0xD(195)(1);
  CNStageIntLLRInputS1xD(187)(3) <= VNStageIntLLROutputS0xD(195)(2);
  CNStageIntLLRInputS1xD(244)(3) <= VNStageIntLLROutputS0xD(195)(3);
  CNStageIntLLRInputS1xD(49)(3) <= VNStageIntLLROutputS0xD(196)(0);
  CNStageIntLLRInputS1xD(64)(3) <= VNStageIntLLROutputS0xD(196)(1);
  CNStageIntLLRInputS1xD(153)(3) <= VNStageIntLLROutputS0xD(196)(2);
  CNStageIntLLRInputS1xD(205)(3) <= VNStageIntLLROutputS0xD(196)(3);
  CNStageIntLLRInputS1xD(242)(3) <= VNStageIntLLROutputS0xD(196)(4);
  CNStageIntLLRInputS1xD(306)(3) <= VNStageIntLLROutputS0xD(196)(5);
  CNStageIntLLRInputS1xD(48)(3) <= VNStageIntLLROutputS0xD(197)(0);
  CNStageIntLLRInputS1xD(96)(3) <= VNStageIntLLROutputS0xD(197)(1);
  CNStageIntLLRInputS1xD(150)(3) <= VNStageIntLLROutputS0xD(197)(2);
  CNStageIntLLRInputS1xD(213)(3) <= VNStageIntLLROutputS0xD(197)(3);
  CNStageIntLLRInputS1xD(273)(3) <= VNStageIntLLROutputS0xD(197)(4);
  CNStageIntLLRInputS1xD(320)(3) <= VNStageIntLLROutputS0xD(197)(5);
  CNStageIntLLRInputS1xD(363)(3) <= VNStageIntLLROutputS0xD(197)(6);
  CNStageIntLLRInputS1xD(47)(3) <= VNStageIntLLROutputS0xD(198)(0);
  CNStageIntLLRInputS1xD(105)(3) <= VNStageIntLLROutputS0xD(198)(1);
  CNStageIntLLRInputS1xD(111)(3) <= VNStageIntLLROutputS0xD(198)(2);
  CNStageIntLLRInputS1xD(208)(3) <= VNStageIntLLROutputS0xD(198)(3);
  CNStageIntLLRInputS1xD(254)(3) <= VNStageIntLLROutputS0xD(198)(4);
  CNStageIntLLRInputS1xD(316)(3) <= VNStageIntLLROutputS0xD(198)(5);
  CNStageIntLLRInputS1xD(379)(3) <= VNStageIntLLROutputS0xD(198)(6);
  CNStageIntLLRInputS1xD(46)(3) <= VNStageIntLLROutputS0xD(199)(0);
  CNStageIntLLRInputS1xD(99)(3) <= VNStageIntLLROutputS0xD(199)(1);
  CNStageIntLLRInputS1xD(133)(3) <= VNStageIntLLROutputS0xD(199)(2);
  CNStageIntLLRInputS1xD(214)(3) <= VNStageIntLLROutputS0xD(199)(3);
  CNStageIntLLRInputS1xD(257)(3) <= VNStageIntLLROutputS0xD(199)(4);
  CNStageIntLLRInputS1xD(282)(3) <= VNStageIntLLROutputS0xD(199)(5);
  CNStageIntLLRInputS1xD(350)(3) <= VNStageIntLLROutputS0xD(199)(6);
  CNStageIntLLRInputS1xD(45)(3) <= VNStageIntLLROutputS0xD(200)(0);
  CNStageIntLLRInputS1xD(102)(3) <= VNStageIntLLROutputS0xD(200)(1);
  CNStageIntLLRInputS1xD(134)(3) <= VNStageIntLLROutputS0xD(200)(2);
  CNStageIntLLRInputS1xD(204)(3) <= VNStageIntLLROutputS0xD(200)(3);
  CNStageIntLLRInputS1xD(245)(3) <= VNStageIntLLROutputS0xD(200)(4);
  CNStageIntLLRInputS1xD(300)(3) <= VNStageIntLLROutputS0xD(200)(5);
  CNStageIntLLRInputS1xD(44)(3) <= VNStageIntLLROutputS0xD(201)(0);
  CNStageIntLLRInputS1xD(93)(3) <= VNStageIntLLROutputS0xD(201)(1);
  CNStageIntLLRInputS1xD(169)(3) <= VNStageIntLLROutputS0xD(201)(2);
  CNStageIntLLRInputS1xD(174)(3) <= VNStageIntLLROutputS0xD(201)(3);
  CNStageIntLLRInputS1xD(274)(3) <= VNStageIntLLROutputS0xD(201)(4);
  CNStageIntLLRInputS1xD(351)(3) <= VNStageIntLLROutputS0xD(201)(5);
  CNStageIntLLRInputS1xD(43)(3) <= VNStageIntLLROutputS0xD(202)(0);
  CNStageIntLLRInputS1xD(73)(3) <= VNStageIntLLROutputS0xD(202)(1);
  CNStageIntLLRInputS1xD(160)(3) <= VNStageIntLLROutputS0xD(202)(2);
  CNStageIntLLRInputS1xD(181)(3) <= VNStageIntLLROutputS0xD(202)(3);
  CNStageIntLLRInputS1xD(281)(3) <= VNStageIntLLROutputS0xD(202)(4);
  CNStageIntLLRInputS1xD(365)(3) <= VNStageIntLLROutputS0xD(202)(5);
  CNStageIntLLRInputS1xD(42)(3) <= VNStageIntLLROutputS0xD(203)(0);
  CNStageIntLLRInputS1xD(54)(3) <= VNStageIntLLROutputS0xD(203)(1);
  CNStageIntLLRInputS1xD(119)(3) <= VNStageIntLLROutputS0xD(203)(2);
  CNStageIntLLRInputS1xD(217)(3) <= VNStageIntLLROutputS0xD(203)(3);
  CNStageIntLLRInputS1xD(267)(3) <= VNStageIntLLROutputS0xD(203)(4);
  CNStageIntLLRInputS1xD(326)(3) <= VNStageIntLLROutputS0xD(203)(5);
  CNStageIntLLRInputS1xD(361)(3) <= VNStageIntLLROutputS0xD(203)(6);
  CNStageIntLLRInputS1xD(41)(3) <= VNStageIntLLROutputS0xD(204)(0);
  CNStageIntLLRInputS1xD(68)(3) <= VNStageIntLLROutputS0xD(204)(1);
  CNStageIntLLRInputS1xD(123)(3) <= VNStageIntLLROutputS0xD(204)(2);
  CNStageIntLLRInputS1xD(219)(3) <= VNStageIntLLROutputS0xD(204)(3);
  CNStageIntLLRInputS1xD(251)(3) <= VNStageIntLLROutputS0xD(204)(4);
  CNStageIntLLRInputS1xD(288)(3) <= VNStageIntLLROutputS0xD(204)(5);
  CNStageIntLLRInputS1xD(382)(3) <= VNStageIntLLROutputS0xD(204)(6);
  CNStageIntLLRInputS1xD(170)(3) <= VNStageIntLLROutputS0xD(205)(0);
  CNStageIntLLRInputS1xD(276)(3) <= VNStageIntLLROutputS0xD(205)(1);
  CNStageIntLLRInputS1xD(345)(3) <= VNStageIntLLROutputS0xD(205)(2);
  CNStageIntLLRInputS1xD(40)(3) <= VNStageIntLLROutputS0xD(206)(0);
  CNStageIntLLRInputS1xD(122)(3) <= VNStageIntLLROutputS0xD(206)(1);
  CNStageIntLLRInputS1xD(172)(3) <= VNStageIntLLROutputS0xD(206)(2);
  CNStageIntLLRInputS1xD(332)(3) <= VNStageIntLLROutputS0xD(206)(3);
  CNStageIntLLRInputS1xD(346)(3) <= VNStageIntLLROutputS0xD(206)(4);
  CNStageIntLLRInputS1xD(39)(3) <= VNStageIntLLROutputS0xD(207)(0);
  CNStageIntLLRInputS1xD(95)(3) <= VNStageIntLLROutputS0xD(207)(1);
  CNStageIntLLRInputS1xD(117)(3) <= VNStageIntLLROutputS0xD(207)(2);
  CNStageIntLLRInputS1xD(255)(3) <= VNStageIntLLROutputS0xD(207)(3);
  CNStageIntLLRInputS1xD(292)(3) <= VNStageIntLLROutputS0xD(207)(4);
  CNStageIntLLRInputS1xD(381)(3) <= VNStageIntLLROutputS0xD(207)(5);
  CNStageIntLLRInputS1xD(38)(3) <= VNStageIntLLROutputS0xD(208)(0);
  CNStageIntLLRInputS1xD(82)(3) <= VNStageIntLLROutputS0xD(208)(1);
  CNStageIntLLRInputS1xD(157)(3) <= VNStageIntLLROutputS0xD(208)(2);
  CNStageIntLLRInputS1xD(191)(3) <= VNStageIntLLROutputS0xD(208)(3);
  CNStageIntLLRInputS1xD(286)(3) <= VNStageIntLLROutputS0xD(208)(4);
  CNStageIntLLRInputS1xD(372)(3) <= VNStageIntLLROutputS0xD(208)(5);
  CNStageIntLLRInputS1xD(37)(3) <= VNStageIntLLROutputS0xD(209)(0);
  CNStageIntLLRInputS1xD(97)(3) <= VNStageIntLLROutputS0xD(209)(1);
  CNStageIntLLRInputS1xD(165)(3) <= VNStageIntLLROutputS0xD(209)(2);
  CNStageIntLLRInputS1xD(218)(3) <= VNStageIntLLROutputS0xD(209)(3);
  CNStageIntLLRInputS1xD(323)(3) <= VNStageIntLLROutputS0xD(209)(4);
  CNStageIntLLRInputS1xD(36)(3) <= VNStageIntLLROutputS0xD(210)(0);
  CNStageIntLLRInputS1xD(60)(3) <= VNStageIntLLROutputS0xD(210)(1);
  CNStageIntLLRInputS1xD(129)(3) <= VNStageIntLLROutputS0xD(210)(2);
  CNStageIntLLRInputS1xD(180)(3) <= VNStageIntLLROutputS0xD(210)(3);
  CNStageIntLLRInputS1xD(246)(3) <= VNStageIntLLROutputS0xD(210)(4);
  CNStageIntLLRInputS1xD(330)(3) <= VNStageIntLLROutputS0xD(210)(5);
  CNStageIntLLRInputS1xD(335)(3) <= VNStageIntLLROutputS0xD(210)(6);
  CNStageIntLLRInputS1xD(35)(3) <= VNStageIntLLROutputS0xD(211)(0);
  CNStageIntLLRInputS1xD(70)(3) <= VNStageIntLLROutputS0xD(211)(1);
  CNStageIntLLRInputS1xD(127)(3) <= VNStageIntLLROutputS0xD(211)(2);
  CNStageIntLLRInputS1xD(206)(3) <= VNStageIntLLROutputS0xD(211)(3);
  CNStageIntLLRInputS1xD(260)(3) <= VNStageIntLLROutputS0xD(211)(4);
  CNStageIntLLRInputS1xD(298)(3) <= VNStageIntLLROutputS0xD(211)(5);
  CNStageIntLLRInputS1xD(34)(3) <= VNStageIntLLROutputS0xD(212)(0);
  CNStageIntLLRInputS1xD(65)(3) <= VNStageIntLLROutputS0xD(212)(1);
  CNStageIntLLRInputS1xD(163)(3) <= VNStageIntLLROutputS0xD(212)(2);
  CNStageIntLLRInputS1xD(186)(3) <= VNStageIntLLROutputS0xD(212)(3);
  CNStageIntLLRInputS1xD(296)(3) <= VNStageIntLLROutputS0xD(212)(4);
  CNStageIntLLRInputS1xD(33)(3) <= VNStageIntLLROutputS0xD(213)(0);
  CNStageIntLLRInputS1xD(71)(3) <= VNStageIntLLROutputS0xD(213)(1);
  CNStageIntLLRInputS1xD(142)(3) <= VNStageIntLLROutputS0xD(213)(2);
  CNStageIntLLRInputS1xD(230)(3) <= VNStageIntLLROutputS0xD(213)(3);
  CNStageIntLLRInputS1xD(32)(3) <= VNStageIntLLROutputS0xD(214)(0);
  CNStageIntLLRInputS1xD(59)(3) <= VNStageIntLLROutputS0xD(214)(1);
  CNStageIntLLRInputS1xD(145)(3) <= VNStageIntLLROutputS0xD(214)(2);
  CNStageIntLLRInputS1xD(220)(3) <= VNStageIntLLROutputS0xD(214)(3);
  CNStageIntLLRInputS1xD(240)(3) <= VNStageIntLLROutputS0xD(214)(4);
  CNStageIntLLRInputS1xD(308)(3) <= VNStageIntLLROutputS0xD(214)(5);
  CNStageIntLLRInputS1xD(369)(3) <= VNStageIntLLROutputS0xD(214)(6);
  CNStageIntLLRInputS1xD(31)(3) <= VNStageIntLLROutputS0xD(215)(0);
  CNStageIntLLRInputS1xD(85)(3) <= VNStageIntLLROutputS0xD(215)(1);
  CNStageIntLLRInputS1xD(130)(3) <= VNStageIntLLROutputS0xD(215)(2);
  CNStageIntLLRInputS1xD(216)(3) <= VNStageIntLLROutputS0xD(215)(3);
  CNStageIntLLRInputS1xD(234)(3) <= VNStageIntLLROutputS0xD(215)(4);
  CNStageIntLLRInputS1xD(311)(3) <= VNStageIntLLROutputS0xD(215)(5);
  CNStageIntLLRInputS1xD(377)(3) <= VNStageIntLLROutputS0xD(215)(6);
  CNStageIntLLRInputS1xD(30)(3) <= VNStageIntLLROutputS0xD(216)(0);
  CNStageIntLLRInputS1xD(91)(3) <= VNStageIntLLROutputS0xD(216)(1);
  CNStageIntLLRInputS1xD(164)(3) <= VNStageIntLLROutputS0xD(216)(2);
  CNStageIntLLRInputS1xD(183)(3) <= VNStageIntLLROutputS0xD(216)(3);
  CNStageIntLLRInputS1xD(237)(3) <= VNStageIntLLROutputS0xD(216)(4);
  CNStageIntLLRInputS1xD(299)(3) <= VNStageIntLLROutputS0xD(216)(5);
  CNStageIntLLRInputS1xD(341)(3) <= VNStageIntLLROutputS0xD(216)(6);
  CNStageIntLLRInputS1xD(29)(3) <= VNStageIntLLROutputS0xD(217)(0);
  CNStageIntLLRInputS1xD(75)(3) <= VNStageIntLLROutputS0xD(217)(1);
  CNStageIntLLRInputS1xD(126)(3) <= VNStageIntLLROutputS0xD(217)(2);
  CNStageIntLLRInputS1xD(201)(3) <= VNStageIntLLROutputS0xD(217)(3);
  CNStageIntLLRInputS1xD(227)(3) <= VNStageIntLLROutputS0xD(217)(4);
  CNStageIntLLRInputS1xD(329)(3) <= VNStageIntLLROutputS0xD(217)(5);
  CNStageIntLLRInputS1xD(339)(3) <= VNStageIntLLROutputS0xD(217)(6);
  CNStageIntLLRInputS1xD(28)(3) <= VNStageIntLLROutputS0xD(218)(0);
  CNStageIntLLRInputS1xD(77)(3) <= VNStageIntLLROutputS0xD(218)(1);
  CNStageIntLLRInputS1xD(154)(3) <= VNStageIntLLROutputS0xD(218)(2);
  CNStageIntLLRInputS1xD(202)(3) <= VNStageIntLLROutputS0xD(218)(3);
  CNStageIntLLRInputS1xD(261)(3) <= VNStageIntLLROutputS0xD(218)(4);
  CNStageIntLLRInputS1xD(295)(3) <= VNStageIntLLROutputS0xD(218)(5);
  CNStageIntLLRInputS1xD(375)(3) <= VNStageIntLLROutputS0xD(218)(6);
  CNStageIntLLRInputS1xD(27)(3) <= VNStageIntLLROutputS0xD(219)(0);
  CNStageIntLLRInputS1xD(101)(3) <= VNStageIntLLROutputS0xD(219)(1);
  CNStageIntLLRInputS1xD(138)(3) <= VNStageIntLLROutputS0xD(219)(2);
  CNStageIntLLRInputS1xD(182)(3) <= VNStageIntLLROutputS0xD(219)(3);
  CNStageIntLLRInputS1xD(321)(3) <= VNStageIntLLROutputS0xD(219)(4);
  CNStageIntLLRInputS1xD(354)(3) <= VNStageIntLLROutputS0xD(219)(5);
  CNStageIntLLRInputS1xD(26)(3) <= VNStageIntLLROutputS0xD(220)(0);
  CNStageIntLLRInputS1xD(83)(3) <= VNStageIntLLROutputS0xD(220)(1);
  CNStageIntLLRInputS1xD(166)(3) <= VNStageIntLLROutputS0xD(220)(2);
  CNStageIntLLRInputS1xD(173)(3) <= VNStageIntLLROutputS0xD(220)(3);
  CNStageIntLLRInputS1xD(256)(3) <= VNStageIntLLROutputS0xD(220)(4);
  CNStageIntLLRInputS1xD(305)(3) <= VNStageIntLLROutputS0xD(220)(5);
  CNStageIntLLRInputS1xD(356)(3) <= VNStageIntLLROutputS0xD(220)(6);
  CNStageIntLLRInputS1xD(25)(3) <= VNStageIntLLROutputS0xD(221)(0);
  CNStageIntLLRInputS1xD(94)(3) <= VNStageIntLLROutputS0xD(221)(1);
  CNStageIntLLRInputS1xD(156)(3) <= VNStageIntLLROutputS0xD(221)(2);
  CNStageIntLLRInputS1xD(190)(3) <= VNStageIntLLROutputS0xD(221)(3);
  CNStageIntLLRInputS1xD(268)(3) <= VNStageIntLLROutputS0xD(221)(4);
  CNStageIntLLRInputS1xD(331)(3) <= VNStageIntLLROutputS0xD(221)(5);
  CNStageIntLLRInputS1xD(342)(3) <= VNStageIntLLROutputS0xD(221)(6);
  CNStageIntLLRInputS1xD(24)(3) <= VNStageIntLLROutputS0xD(222)(0);
  CNStageIntLLRInputS1xD(143)(3) <= VNStageIntLLROutputS0xD(222)(1);
  CNStageIntLLRInputS1xD(241)(3) <= VNStageIntLLROutputS0xD(222)(2);
  CNStageIntLLRInputS1xD(376)(3) <= VNStageIntLLROutputS0xD(222)(3);
  CNStageIntLLRInputS1xD(23)(3) <= VNStageIntLLROutputS0xD(223)(0);
  CNStageIntLLRInputS1xD(76)(3) <= VNStageIntLLROutputS0xD(223)(1);
  CNStageIntLLRInputS1xD(162)(3) <= VNStageIntLLROutputS0xD(223)(2);
  CNStageIntLLRInputS1xD(224)(3) <= VNStageIntLLROutputS0xD(223)(3);
  CNStageIntLLRInputS1xD(229)(3) <= VNStageIntLLROutputS0xD(223)(4);
  CNStageIntLLRInputS1xD(309)(3) <= VNStageIntLLROutputS0xD(223)(5);
  CNStageIntLLRInputS1xD(338)(3) <= VNStageIntLLROutputS0xD(223)(6);
  CNStageIntLLRInputS1xD(22)(3) <= VNStageIntLLROutputS0xD(224)(0);
  CNStageIntLLRInputS1xD(90)(3) <= VNStageIntLLROutputS0xD(224)(1);
  CNStageIntLLRInputS1xD(135)(3) <= VNStageIntLLROutputS0xD(224)(2);
  CNStageIntLLRInputS1xD(193)(3) <= VNStageIntLLROutputS0xD(224)(3);
  CNStageIntLLRInputS1xD(270)(3) <= VNStageIntLLROutputS0xD(224)(4);
  CNStageIntLLRInputS1xD(328)(3) <= VNStageIntLLROutputS0xD(224)(5);
  CNStageIntLLRInputS1xD(366)(3) <= VNStageIntLLROutputS0xD(224)(6);
  CNStageIntLLRInputS1xD(21)(3) <= VNStageIntLLROutputS0xD(225)(0);
  CNStageIntLLRInputS1xD(61)(3) <= VNStageIntLLROutputS0xD(225)(1);
  CNStageIntLLRInputS1xD(132)(3) <= VNStageIntLLROutputS0xD(225)(2);
  CNStageIntLLRInputS1xD(188)(3) <= VNStageIntLLROutputS0xD(225)(3);
  CNStageIntLLRInputS1xD(232)(3) <= VNStageIntLLROutputS0xD(225)(4);
  CNStageIntLLRInputS1xD(301)(3) <= VNStageIntLLROutputS0xD(225)(5);
  CNStageIntLLRInputS1xD(20)(3) <= VNStageIntLLROutputS0xD(226)(0);
  CNStageIntLLRInputS1xD(148)(3) <= VNStageIntLLROutputS0xD(226)(1);
  CNStageIntLLRInputS1xD(378)(3) <= VNStageIntLLROutputS0xD(226)(2);
  CNStageIntLLRInputS1xD(19)(3) <= VNStageIntLLROutputS0xD(227)(0);
  CNStageIntLLRInputS1xD(63)(3) <= VNStageIntLLROutputS0xD(227)(1);
  CNStageIntLLRInputS1xD(140)(3) <= VNStageIntLLROutputS0xD(227)(2);
  CNStageIntLLRInputS1xD(178)(3) <= VNStageIntLLROutputS0xD(227)(3);
  CNStageIntLLRInputS1xD(258)(3) <= VNStageIntLLROutputS0xD(227)(4);
  CNStageIntLLRInputS1xD(314)(3) <= VNStageIntLLROutputS0xD(227)(5);
  CNStageIntLLRInputS1xD(368)(3) <= VNStageIntLLROutputS0xD(227)(6);
  CNStageIntLLRInputS1xD(18)(3) <= VNStageIntLLROutputS0xD(228)(0);
  CNStageIntLLRInputS1xD(78)(3) <= VNStageIntLLROutputS0xD(228)(1);
  CNStageIntLLRInputS1xD(114)(3) <= VNStageIntLLROutputS0xD(228)(2);
  CNStageIntLLRInputS1xD(198)(3) <= VNStageIntLLROutputS0xD(228)(3);
  CNStageIntLLRInputS1xD(253)(3) <= VNStageIntLLROutputS0xD(228)(4);
  CNStageIntLLRInputS1xD(307)(3) <= VNStageIntLLROutputS0xD(228)(5);
  CNStageIntLLRInputS1xD(17)(3) <= VNStageIntLLROutputS0xD(229)(0);
  CNStageIntLLRInputS1xD(74)(3) <= VNStageIntLLROutputS0xD(229)(1);
  CNStageIntLLRInputS1xD(124)(3) <= VNStageIntLLROutputS0xD(229)(2);
  CNStageIntLLRInputS1xD(259)(3) <= VNStageIntLLROutputS0xD(229)(3);
  CNStageIntLLRInputS1xD(374)(3) <= VNStageIntLLROutputS0xD(229)(4);
  CNStageIntLLRInputS1xD(16)(3) <= VNStageIntLLROutputS0xD(230)(0);
  CNStageIntLLRInputS1xD(118)(3) <= VNStageIntLLROutputS0xD(230)(1);
  CNStageIntLLRInputS1xD(176)(3) <= VNStageIntLLROutputS0xD(230)(2);
  CNStageIntLLRInputS1xD(249)(3) <= VNStageIntLLROutputS0xD(230)(3);
  CNStageIntLLRInputS1xD(293)(3) <= VNStageIntLLROutputS0xD(230)(4);
  CNStageIntLLRInputS1xD(347)(3) <= VNStageIntLLROutputS0xD(230)(5);
  CNStageIntLLRInputS1xD(15)(3) <= VNStageIntLLROutputS0xD(231)(0);
  CNStageIntLLRInputS1xD(56)(3) <= VNStageIntLLROutputS0xD(231)(1);
  CNStageIntLLRInputS1xD(209)(3) <= VNStageIntLLROutputS0xD(231)(2);
  CNStageIntLLRInputS1xD(272)(3) <= VNStageIntLLROutputS0xD(231)(3);
  CNStageIntLLRInputS1xD(287)(3) <= VNStageIntLLROutputS0xD(231)(4);
  CNStageIntLLRInputS1xD(344)(3) <= VNStageIntLLROutputS0xD(231)(5);
  CNStageIntLLRInputS1xD(14)(3) <= VNStageIntLLROutputS0xD(232)(0);
  CNStageIntLLRInputS1xD(57)(3) <= VNStageIntLLROutputS0xD(232)(1);
  CNStageIntLLRInputS1xD(212)(3) <= VNStageIntLLROutputS0xD(232)(2);
  CNStageIntLLRInputS1xD(278)(3) <= VNStageIntLLROutputS0xD(232)(3);
  CNStageIntLLRInputS1xD(291)(3) <= VNStageIntLLROutputS0xD(232)(4);
  CNStageIntLLRInputS1xD(359)(3) <= VNStageIntLLROutputS0xD(232)(5);
  CNStageIntLLRInputS1xD(13)(3) <= VNStageIntLLROutputS0xD(233)(0);
  CNStageIntLLRInputS1xD(92)(3) <= VNStageIntLLROutputS0xD(233)(1);
  CNStageIntLLRInputS1xD(149)(3) <= VNStageIntLLROutputS0xD(233)(2);
  CNStageIntLLRInputS1xD(263)(3) <= VNStageIntLLROutputS0xD(233)(3);
  CNStageIntLLRInputS1xD(352)(3) <= VNStageIntLLROutputS0xD(233)(4);
  CNStageIntLLRInputS1xD(12)(3) <= VNStageIntLLROutputS0xD(234)(0);
  CNStageIntLLRInputS1xD(84)(3) <= VNStageIntLLROutputS0xD(234)(1);
  CNStageIntLLRInputS1xD(131)(3) <= VNStageIntLLROutputS0xD(234)(2);
  CNStageIntLLRInputS1xD(177)(3) <= VNStageIntLLROutputS0xD(234)(3);
  CNStageIntLLRInputS1xD(265)(3) <= VNStageIntLLROutputS0xD(234)(4);
  CNStageIntLLRInputS1xD(315)(3) <= VNStageIntLLROutputS0xD(234)(5);
  CNStageIntLLRInputS1xD(100)(3) <= VNStageIntLLROutputS0xD(235)(0);
  CNStageIntLLRInputS1xD(144)(3) <= VNStageIntLLROutputS0xD(235)(1);
  CNStageIntLLRInputS1xD(196)(3) <= VNStageIntLLROutputS0xD(235)(2);
  CNStageIntLLRInputS1xD(235)(3) <= VNStageIntLLROutputS0xD(235)(3);
  CNStageIntLLRInputS1xD(336)(3) <= VNStageIntLLROutputS0xD(235)(4);
  CNStageIntLLRInputS1xD(11)(3) <= VNStageIntLLROutputS0xD(236)(0);
  CNStageIntLLRInputS1xD(104)(3) <= VNStageIntLLROutputS0xD(236)(1);
  CNStageIntLLRInputS1xD(155)(3) <= VNStageIntLLROutputS0xD(236)(2);
  CNStageIntLLRInputS1xD(221)(3) <= VNStageIntLLROutputS0xD(236)(3);
  CNStageIntLLRInputS1xD(271)(3) <= VNStageIntLLROutputS0xD(236)(4);
  CNStageIntLLRInputS1xD(310)(3) <= VNStageIntLLROutputS0xD(236)(5);
  CNStageIntLLRInputS1xD(10)(3) <= VNStageIntLLROutputS0xD(237)(0);
  CNStageIntLLRInputS1xD(110)(3) <= VNStageIntLLROutputS0xD(237)(1);
  CNStageIntLLRInputS1xD(125)(3) <= VNStageIntLLROutputS0xD(237)(2);
  CNStageIntLLRInputS1xD(228)(3) <= VNStageIntLLROutputS0xD(237)(3);
  CNStageIntLLRInputS1xD(322)(3) <= VNStageIntLLROutputS0xD(237)(4);
  CNStageIntLLRInputS1xD(334)(3) <= VNStageIntLLROutputS0xD(237)(5);
  CNStageIntLLRInputS1xD(9)(3) <= VNStageIntLLROutputS0xD(238)(0);
  CNStageIntLLRInputS1xD(103)(3) <= VNStageIntLLROutputS0xD(238)(1);
  CNStageIntLLRInputS1xD(113)(3) <= VNStageIntLLROutputS0xD(238)(2);
  CNStageIntLLRInputS1xD(179)(3) <= VNStageIntLLROutputS0xD(238)(3);
  CNStageIntLLRInputS1xD(236)(3) <= VNStageIntLLROutputS0xD(238)(4);
  CNStageIntLLRInputS1xD(294)(3) <= VNStageIntLLROutputS0xD(238)(5);
  CNStageIntLLRInputS1xD(383)(3) <= VNStageIntLLROutputS0xD(238)(6);
  CNStageIntLLRInputS1xD(8)(3) <= VNStageIntLLROutputS0xD(239)(0);
  CNStageIntLLRInputS1xD(98)(3) <= VNStageIntLLROutputS0xD(239)(1);
  CNStageIntLLRInputS1xD(158)(3) <= VNStageIntLLROutputS0xD(239)(2);
  CNStageIntLLRInputS1xD(223)(3) <= VNStageIntLLROutputS0xD(239)(3);
  CNStageIntLLRInputS1xD(264)(3) <= VNStageIntLLROutputS0xD(239)(4);
  CNStageIntLLRInputS1xD(284)(3) <= VNStageIntLLROutputS0xD(239)(5);
  CNStageIntLLRInputS1xD(360)(3) <= VNStageIntLLROutputS0xD(239)(6);
  CNStageIntLLRInputS1xD(7)(3) <= VNStageIntLLROutputS0xD(240)(0);
  CNStageIntLLRInputS1xD(81)(3) <= VNStageIntLLROutputS0xD(240)(1);
  CNStageIntLLRInputS1xD(116)(3) <= VNStageIntLLROutputS0xD(240)(2);
  CNStageIntLLRInputS1xD(210)(3) <= VNStageIntLLROutputS0xD(240)(3);
  CNStageIntLLRInputS1xD(277)(3) <= VNStageIntLLROutputS0xD(240)(4);
  CNStageIntLLRInputS1xD(324)(3) <= VNStageIntLLROutputS0xD(240)(5);
  CNStageIntLLRInputS1xD(343)(3) <= VNStageIntLLROutputS0xD(240)(6);
  CNStageIntLLRInputS1xD(6)(3) <= VNStageIntLLROutputS0xD(241)(0);
  CNStageIntLLRInputS1xD(88)(3) <= VNStageIntLLROutputS0xD(241)(1);
  CNStageIntLLRInputS1xD(175)(3) <= VNStageIntLLROutputS0xD(241)(2);
  CNStageIntLLRInputS1xD(250)(3) <= VNStageIntLLROutputS0xD(241)(3);
  CNStageIntLLRInputS1xD(285)(3) <= VNStageIntLLROutputS0xD(241)(4);
  CNStageIntLLRInputS1xD(355)(3) <= VNStageIntLLROutputS0xD(241)(5);
  CNStageIntLLRInputS1xD(5)(3) <= VNStageIntLLROutputS0xD(242)(0);
  CNStageIntLLRInputS1xD(108)(3) <= VNStageIntLLROutputS0xD(242)(1);
  CNStageIntLLRInputS1xD(146)(3) <= VNStageIntLLROutputS0xD(242)(2);
  CNStageIntLLRInputS1xD(203)(3) <= VNStageIntLLROutputS0xD(242)(3);
  CNStageIntLLRInputS1xD(231)(3) <= VNStageIntLLROutputS0xD(242)(4);
  CNStageIntLLRInputS1xD(303)(3) <= VNStageIntLLROutputS0xD(242)(5);
  CNStageIntLLRInputS1xD(367)(3) <= VNStageIntLLROutputS0xD(242)(6);
  CNStageIntLLRInputS1xD(4)(3) <= VNStageIntLLROutputS0xD(243)(0);
  CNStageIntLLRInputS1xD(106)(3) <= VNStageIntLLROutputS0xD(243)(1);
  CNStageIntLLRInputS1xD(141)(3) <= VNStageIntLLROutputS0xD(243)(2);
  CNStageIntLLRInputS1xD(200)(3) <= VNStageIntLLROutputS0xD(243)(3);
  CNStageIntLLRInputS1xD(252)(3) <= VNStageIntLLROutputS0xD(243)(4);
  CNStageIntLLRInputS1xD(312)(3) <= VNStageIntLLROutputS0xD(243)(5);
  CNStageIntLLRInputS1xD(337)(3) <= VNStageIntLLROutputS0xD(243)(6);
  CNStageIntLLRInputS1xD(147)(3) <= VNStageIntLLROutputS0xD(244)(0);
  CNStageIntLLRInputS1xD(266)(3) <= VNStageIntLLROutputS0xD(244)(1);
  CNStageIntLLRInputS1xD(3)(3) <= VNStageIntLLROutputS0xD(245)(0);
  CNStageIntLLRInputS1xD(66)(3) <= VNStageIntLLROutputS0xD(245)(1);
  CNStageIntLLRInputS1xD(136)(3) <= VNStageIntLLROutputS0xD(245)(2);
  CNStageIntLLRInputS1xD(207)(3) <= VNStageIntLLROutputS0xD(245)(3);
  CNStageIntLLRInputS1xD(262)(3) <= VNStageIntLLROutputS0xD(245)(4);
  CNStageIntLLRInputS1xD(313)(3) <= VNStageIntLLROutputS0xD(245)(5);
  CNStageIntLLRInputS1xD(370)(3) <= VNStageIntLLROutputS0xD(245)(6);
  CNStageIntLLRInputS1xD(2)(3) <= VNStageIntLLROutputS0xD(246)(0);
  CNStageIntLLRInputS1xD(69)(3) <= VNStageIntLLROutputS0xD(246)(1);
  CNStageIntLLRInputS1xD(161)(3) <= VNStageIntLLROutputS0xD(246)(2);
  CNStageIntLLRInputS1xD(185)(3) <= VNStageIntLLROutputS0xD(246)(3);
  CNStageIntLLRInputS1xD(226)(3) <= VNStageIntLLROutputS0xD(246)(4);
  CNStageIntLLRInputS1xD(302)(3) <= VNStageIntLLROutputS0xD(246)(5);
  CNStageIntLLRInputS1xD(1)(3) <= VNStageIntLLROutputS0xD(247)(0);
  CNStageIntLLRInputS1xD(109)(3) <= VNStageIntLLROutputS0xD(247)(1);
  CNStageIntLLRInputS1xD(168)(3) <= VNStageIntLLROutputS0xD(247)(2);
  CNStageIntLLRInputS1xD(194)(3) <= VNStageIntLLROutputS0xD(247)(3);
  CNStageIntLLRInputS1xD(247)(3) <= VNStageIntLLROutputS0xD(247)(4);
  CNStageIntLLRInputS1xD(327)(3) <= VNStageIntLLROutputS0xD(247)(5);
  CNStageIntLLRInputS1xD(349)(3) <= VNStageIntLLROutputS0xD(247)(6);
  CNStageIntLLRInputS1xD(0)(3) <= VNStageIntLLROutputS0xD(248)(0);
  CNStageIntLLRInputS1xD(87)(3) <= VNStageIntLLROutputS0xD(248)(1);
  CNStageIntLLRInputS1xD(151)(3) <= VNStageIntLLROutputS0xD(248)(2);
  CNStageIntLLRInputS1xD(189)(3) <= VNStageIntLLROutputS0xD(248)(3);
  CNStageIntLLRInputS1xD(248)(3) <= VNStageIntLLROutputS0xD(248)(4);
  CNStageIntLLRInputS1xD(280)(3) <= VNStageIntLLROutputS0xD(248)(5);
  CNStageIntLLRInputS1xD(357)(3) <= VNStageIntLLROutputS0xD(248)(6);
  CNStageIntLLRInputS1xD(152)(3) <= VNStageIntLLROutputS0xD(249)(0);
  CNStageIntLLRInputS1xD(192)(3) <= VNStageIntLLROutputS0xD(249)(1);
  CNStageIntLLRInputS1xD(225)(3) <= VNStageIntLLROutputS0xD(249)(2);
  CNStageIntLLRInputS1xD(317)(3) <= VNStageIntLLROutputS0xD(249)(3);
  CNStageIntLLRInputS1xD(353)(3) <= VNStageIntLLROutputS0xD(249)(4);
  CNStageIntLLRInputS1xD(79)(3) <= VNStageIntLLROutputS0xD(250)(0);
  CNStageIntLLRInputS1xD(120)(3) <= VNStageIntLLROutputS0xD(250)(1);
  CNStageIntLLRInputS1xD(184)(3) <= VNStageIntLLROutputS0xD(250)(2);
  CNStageIntLLRInputS1xD(319)(3) <= VNStageIntLLROutputS0xD(250)(3);
  CNStageIntLLRInputS1xD(358)(3) <= VNStageIntLLROutputS0xD(250)(4);
  CNStageIntLLRInputS1xD(62)(3) <= VNStageIntLLROutputS0xD(251)(0);
  CNStageIntLLRInputS1xD(159)(3) <= VNStageIntLLROutputS0xD(251)(1);
  CNStageIntLLRInputS1xD(215)(3) <= VNStageIntLLROutputS0xD(251)(2);
  CNStageIntLLRInputS1xD(289)(3) <= VNStageIntLLROutputS0xD(251)(3);
  CNStageIntLLRInputS1xD(348)(3) <= VNStageIntLLROutputS0xD(251)(4);
  CNStageIntLLRInputS1xD(89)(3) <= VNStageIntLLROutputS0xD(252)(0);
  CNStageIntLLRInputS1xD(112)(3) <= VNStageIntLLROutputS0xD(252)(1);
  CNStageIntLLRInputS1xD(199)(3) <= VNStageIntLLROutputS0xD(252)(2);
  CNStageIntLLRInputS1xD(239)(3) <= VNStageIntLLROutputS0xD(252)(3);
  CNStageIntLLRInputS1xD(325)(3) <= VNStageIntLLROutputS0xD(252)(4);
  CNStageIntLLRInputS1xD(373)(3) <= VNStageIntLLROutputS0xD(252)(5);
  CNStageIntLLRInputS1xD(80)(3) <= VNStageIntLLROutputS0xD(253)(0);
  CNStageIntLLRInputS1xD(121)(3) <= VNStageIntLLROutputS0xD(253)(1);
  CNStageIntLLRInputS1xD(211)(3) <= VNStageIntLLROutputS0xD(253)(2);
  CNStageIntLLRInputS1xD(279)(3) <= VNStageIntLLROutputS0xD(253)(3);
  CNStageIntLLRInputS1xD(283)(3) <= VNStageIntLLROutputS0xD(253)(4);
  CNStageIntLLRInputS1xD(380)(3) <= VNStageIntLLROutputS0xD(253)(5);
  CNStageIntLLRInputS1xD(67)(3) <= VNStageIntLLROutputS0xD(254)(0);
  CNStageIntLLRInputS1xD(222)(3) <= VNStageIntLLROutputS0xD(254)(1);
  CNStageIntLLRInputS1xD(238)(3) <= VNStageIntLLROutputS0xD(254)(2);
  CNStageIntLLRInputS1xD(290)(3) <= VNStageIntLLROutputS0xD(254)(3);
  CNStageIntLLRInputS1xD(362)(3) <= VNStageIntLLROutputS0xD(254)(4);
  CNStageIntLLRInputS1xD(52)(3) <= VNStageIntLLROutputS0xD(255)(0);
  CNStageIntLLRInputS1xD(86)(3) <= VNStageIntLLROutputS0xD(255)(1);
  CNStageIntLLRInputS1xD(167)(3) <= VNStageIntLLROutputS0xD(255)(2);
  CNStageIntLLRInputS1xD(195)(3) <= VNStageIntLLROutputS0xD(255)(3);
  CNStageIntLLRInputS1xD(233)(3) <= VNStageIntLLROutputS0xD(255)(4);
  CNStageIntLLRInputS1xD(318)(3) <= VNStageIntLLROutputS0xD(255)(5);
  CNStageIntLLRInputS1xD(364)(3) <= VNStageIntLLROutputS0xD(255)(6);
  CNStageIntLLRInputS1xD(53)(4) <= VNStageIntLLROutputS0xD(256)(0);
  CNStageIntLLRInputS1xD(106)(4) <= VNStageIntLLROutputS0xD(256)(1);
  CNStageIntLLRInputS1xD(127)(4) <= VNStageIntLLROutputS0xD(256)(2);
  CNStageIntLLRInputS1xD(242)(4) <= VNStageIntLLROutputS0xD(256)(3);
  CNStageIntLLRInputS1xD(296)(4) <= VNStageIntLLROutputS0xD(256)(4);
  CNStageIntLLRInputS1xD(339)(4) <= VNStageIntLLROutputS0xD(256)(5);
  CNStageIntLLRInputS1xD(51)(4) <= VNStageIntLLROutputS0xD(257)(0);
  CNStageIntLLRInputS1xD(85)(4) <= VNStageIntLLROutputS0xD(257)(1);
  CNStageIntLLRInputS1xD(166)(4) <= VNStageIntLLROutputS0xD(257)(2);
  CNStageIntLLRInputS1xD(194)(4) <= VNStageIntLLROutputS0xD(257)(3);
  CNStageIntLLRInputS1xD(232)(4) <= VNStageIntLLROutputS0xD(257)(4);
  CNStageIntLLRInputS1xD(317)(4) <= VNStageIntLLROutputS0xD(257)(5);
  CNStageIntLLRInputS1xD(363)(4) <= VNStageIntLLROutputS0xD(257)(6);
  CNStageIntLLRInputS1xD(50)(4) <= VNStageIntLLROutputS0xD(258)(0);
  CNStageIntLLRInputS1xD(57)(4) <= VNStageIntLLROutputS0xD(258)(1);
  CNStageIntLLRInputS1xD(331)(4) <= VNStageIntLLROutputS0xD(258)(2);
  CNStageIntLLRInputS1xD(54)(4) <= VNStageIntLLROutputS0xD(259)(0);
  CNStageIntLLRInputS1xD(114)(4) <= VNStageIntLLROutputS0xD(259)(1);
  CNStageIntLLRInputS1xD(274)(4) <= VNStageIntLLROutputS0xD(259)(2);
  CNStageIntLLRInputS1xD(303)(4) <= VNStageIntLLROutputS0xD(259)(3);
  CNStageIntLLRInputS1xD(370)(4) <= VNStageIntLLROutputS0xD(259)(4);
  CNStageIntLLRInputS1xD(49)(4) <= VNStageIntLLROutputS0xD(260)(0);
  CNStageIntLLRInputS1xD(71)(4) <= VNStageIntLLROutputS0xD(260)(1);
  CNStageIntLLRInputS1xD(138)(4) <= VNStageIntLLROutputS0xD(260)(2);
  CNStageIntLLRInputS1xD(186)(4) <= VNStageIntLLROutputS0xD(260)(3);
  CNStageIntLLRInputS1xD(243)(4) <= VNStageIntLLROutputS0xD(260)(4);
  CNStageIntLLRInputS1xD(383)(4) <= VNStageIntLLROutputS0xD(260)(5);
  CNStageIntLLRInputS1xD(48)(4) <= VNStageIntLLROutputS0xD(261)(0);
  CNStageIntLLRInputS1xD(63)(4) <= VNStageIntLLROutputS0xD(261)(1);
  CNStageIntLLRInputS1xD(152)(4) <= VNStageIntLLROutputS0xD(261)(2);
  CNStageIntLLRInputS1xD(204)(4) <= VNStageIntLLROutputS0xD(261)(3);
  CNStageIntLLRInputS1xD(305)(4) <= VNStageIntLLROutputS0xD(261)(4);
  CNStageIntLLRInputS1xD(333)(4) <= VNStageIntLLROutputS0xD(261)(5);
  CNStageIntLLRInputS1xD(47)(4) <= VNStageIntLLROutputS0xD(262)(0);
  CNStageIntLLRInputS1xD(95)(4) <= VNStageIntLLROutputS0xD(262)(1);
  CNStageIntLLRInputS1xD(149)(4) <= VNStageIntLLROutputS0xD(262)(2);
  CNStageIntLLRInputS1xD(212)(4) <= VNStageIntLLROutputS0xD(262)(3);
  CNStageIntLLRInputS1xD(319)(4) <= VNStageIntLLROutputS0xD(262)(4);
  CNStageIntLLRInputS1xD(362)(4) <= VNStageIntLLROutputS0xD(262)(5);
  CNStageIntLLRInputS1xD(46)(4) <= VNStageIntLLROutputS0xD(263)(0);
  CNStageIntLLRInputS1xD(104)(4) <= VNStageIntLLROutputS0xD(263)(1);
  CNStageIntLLRInputS1xD(169)(4) <= VNStageIntLLROutputS0xD(263)(2);
  CNStageIntLLRInputS1xD(207)(4) <= VNStageIntLLROutputS0xD(263)(3);
  CNStageIntLLRInputS1xD(253)(4) <= VNStageIntLLROutputS0xD(263)(4);
  CNStageIntLLRInputS1xD(315)(4) <= VNStageIntLLROutputS0xD(263)(5);
  CNStageIntLLRInputS1xD(378)(4) <= VNStageIntLLROutputS0xD(263)(6);
  CNStageIntLLRInputS1xD(45)(4) <= VNStageIntLLROutputS0xD(264)(0);
  CNStageIntLLRInputS1xD(98)(4) <= VNStageIntLLROutputS0xD(264)(1);
  CNStageIntLLRInputS1xD(132)(4) <= VNStageIntLLROutputS0xD(264)(2);
  CNStageIntLLRInputS1xD(213)(4) <= VNStageIntLLROutputS0xD(264)(3);
  CNStageIntLLRInputS1xD(256)(4) <= VNStageIntLLROutputS0xD(264)(4);
  CNStageIntLLRInputS1xD(281)(4) <= VNStageIntLLROutputS0xD(264)(5);
  CNStageIntLLRInputS1xD(349)(4) <= VNStageIntLLROutputS0xD(264)(6);
  CNStageIntLLRInputS1xD(44)(4) <= VNStageIntLLROutputS0xD(265)(0);
  CNStageIntLLRInputS1xD(133)(4) <= VNStageIntLLROutputS0xD(265)(1);
  CNStageIntLLRInputS1xD(203)(4) <= VNStageIntLLROutputS0xD(265)(2);
  CNStageIntLLRInputS1xD(244)(4) <= VNStageIntLLROutputS0xD(265)(3);
  CNStageIntLLRInputS1xD(43)(4) <= VNStageIntLLROutputS0xD(266)(0);
  CNStageIntLLRInputS1xD(168)(4) <= VNStageIntLLROutputS0xD(266)(1);
  CNStageIntLLRInputS1xD(173)(4) <= VNStageIntLLROutputS0xD(266)(2);
  CNStageIntLLRInputS1xD(273)(4) <= VNStageIntLLROutputS0xD(266)(3);
  CNStageIntLLRInputS1xD(300)(4) <= VNStageIntLLROutputS0xD(266)(4);
  CNStageIntLLRInputS1xD(42)(4) <= VNStageIntLLROutputS0xD(267)(0);
  CNStageIntLLRInputS1xD(72)(4) <= VNStageIntLLROutputS0xD(267)(1);
  CNStageIntLLRInputS1xD(159)(4) <= VNStageIntLLROutputS0xD(267)(2);
  CNStageIntLLRInputS1xD(180)(4) <= VNStageIntLLROutputS0xD(267)(3);
  CNStageIntLLRInputS1xD(241)(4) <= VNStageIntLLROutputS0xD(267)(4);
  CNStageIntLLRInputS1xD(280)(4) <= VNStageIntLLROutputS0xD(267)(5);
  CNStageIntLLRInputS1xD(364)(4) <= VNStageIntLLROutputS0xD(267)(6);
  CNStageIntLLRInputS1xD(41)(4) <= VNStageIntLLROutputS0xD(268)(0);
  CNStageIntLLRInputS1xD(109)(4) <= VNStageIntLLROutputS0xD(268)(1);
  CNStageIntLLRInputS1xD(118)(4) <= VNStageIntLLROutputS0xD(268)(2);
  CNStageIntLLRInputS1xD(216)(4) <= VNStageIntLLROutputS0xD(268)(3);
  CNStageIntLLRInputS1xD(266)(4) <= VNStageIntLLROutputS0xD(268)(4);
  CNStageIntLLRInputS1xD(325)(4) <= VNStageIntLLROutputS0xD(268)(5);
  CNStageIntLLRInputS1xD(360)(4) <= VNStageIntLLROutputS0xD(268)(6);
  CNStageIntLLRInputS1xD(67)(4) <= VNStageIntLLROutputS0xD(269)(0);
  CNStageIntLLRInputS1xD(122)(4) <= VNStageIntLLROutputS0xD(269)(1);
  CNStageIntLLRInputS1xD(218)(4) <= VNStageIntLLROutputS0xD(269)(2);
  CNStageIntLLRInputS1xD(250)(4) <= VNStageIntLLROutputS0xD(269)(3);
  CNStageIntLLRInputS1xD(287)(4) <= VNStageIntLLROutputS0xD(269)(4);
  CNStageIntLLRInputS1xD(381)(4) <= VNStageIntLLROutputS0xD(269)(5);
  CNStageIntLLRInputS1xD(40)(4) <= VNStageIntLLROutputS0xD(270)(0);
  CNStageIntLLRInputS1xD(79)(4) <= VNStageIntLLROutputS0xD(270)(1);
  CNStageIntLLRInputS1xD(170)(4) <= VNStageIntLLROutputS0xD(270)(2);
  CNStageIntLLRInputS1xD(190)(4) <= VNStageIntLLROutputS0xD(270)(3);
  CNStageIntLLRInputS1xD(275)(4) <= VNStageIntLLROutputS0xD(270)(4);
  CNStageIntLLRInputS1xD(292)(4) <= VNStageIntLLROutputS0xD(270)(5);
  CNStageIntLLRInputS1xD(344)(4) <= VNStageIntLLROutputS0xD(270)(6);
  CNStageIntLLRInputS1xD(39)(4) <= VNStageIntLLROutputS0xD(271)(0);
  CNStageIntLLRInputS1xD(105)(4) <= VNStageIntLLROutputS0xD(271)(1);
  CNStageIntLLRInputS1xD(171)(4) <= VNStageIntLLROutputS0xD(271)(2);
  CNStageIntLLRInputS1xD(268)(4) <= VNStageIntLLROutputS0xD(271)(3);
  CNStageIntLLRInputS1xD(332)(4) <= VNStageIntLLROutputS0xD(271)(4);
  CNStageIntLLRInputS1xD(345)(4) <= VNStageIntLLROutputS0xD(271)(5);
  CNStageIntLLRInputS1xD(38)(4) <= VNStageIntLLROutputS0xD(272)(0);
  CNStageIntLLRInputS1xD(94)(4) <= VNStageIntLLROutputS0xD(272)(1);
  CNStageIntLLRInputS1xD(116)(4) <= VNStageIntLLROutputS0xD(272)(2);
  CNStageIntLLRInputS1xD(184)(4) <= VNStageIntLLROutputS0xD(272)(3);
  CNStageIntLLRInputS1xD(254)(4) <= VNStageIntLLROutputS0xD(272)(4);
  CNStageIntLLRInputS1xD(291)(4) <= VNStageIntLLROutputS0xD(272)(5);
  CNStageIntLLRInputS1xD(380)(4) <= VNStageIntLLROutputS0xD(272)(6);
  CNStageIntLLRInputS1xD(37)(4) <= VNStageIntLLROutputS0xD(273)(0);
  CNStageIntLLRInputS1xD(81)(4) <= VNStageIntLLROutputS0xD(273)(1);
  CNStageIntLLRInputS1xD(156)(4) <= VNStageIntLLROutputS0xD(273)(2);
  CNStageIntLLRInputS1xD(272)(4) <= VNStageIntLLROutputS0xD(273)(3);
  CNStageIntLLRInputS1xD(285)(4) <= VNStageIntLLROutputS0xD(273)(4);
  CNStageIntLLRInputS1xD(371)(4) <= VNStageIntLLROutputS0xD(273)(5);
  CNStageIntLLRInputS1xD(36)(4) <= VNStageIntLLROutputS0xD(274)(0);
  CNStageIntLLRInputS1xD(164)(4) <= VNStageIntLLROutputS0xD(274)(1);
  CNStageIntLLRInputS1xD(217)(4) <= VNStageIntLLROutputS0xD(274)(2);
  CNStageIntLLRInputS1xD(248)(4) <= VNStageIntLLROutputS0xD(274)(3);
  CNStageIntLLRInputS1xD(35)(4) <= VNStageIntLLROutputS0xD(275)(0);
  CNStageIntLLRInputS1xD(59)(4) <= VNStageIntLLROutputS0xD(275)(1);
  CNStageIntLLRInputS1xD(128)(4) <= VNStageIntLLROutputS0xD(275)(2);
  CNStageIntLLRInputS1xD(179)(4) <= VNStageIntLLROutputS0xD(275)(3);
  CNStageIntLLRInputS1xD(329)(4) <= VNStageIntLLROutputS0xD(275)(4);
  CNStageIntLLRInputS1xD(34)(4) <= VNStageIntLLROutputS0xD(276)(0);
  CNStageIntLLRInputS1xD(69)(4) <= VNStageIntLLROutputS0xD(276)(1);
  CNStageIntLLRInputS1xD(126)(4) <= VNStageIntLLROutputS0xD(276)(2);
  CNStageIntLLRInputS1xD(205)(4) <= VNStageIntLLROutputS0xD(276)(3);
  CNStageIntLLRInputS1xD(259)(4) <= VNStageIntLLROutputS0xD(276)(4);
  CNStageIntLLRInputS1xD(297)(4) <= VNStageIntLLROutputS0xD(276)(5);
  CNStageIntLLRInputS1xD(33)(4) <= VNStageIntLLROutputS0xD(277)(0);
  CNStageIntLLRInputS1xD(64)(4) <= VNStageIntLLROutputS0xD(277)(1);
  CNStageIntLLRInputS1xD(162)(4) <= VNStageIntLLROutputS0xD(277)(2);
  CNStageIntLLRInputS1xD(185)(4) <= VNStageIntLLROutputS0xD(277)(3);
  CNStageIntLLRInputS1xD(252)(4) <= VNStageIntLLROutputS0xD(277)(4);
  CNStageIntLLRInputS1xD(295)(4) <= VNStageIntLLROutputS0xD(277)(5);
  CNStageIntLLRInputS1xD(334)(4) <= VNStageIntLLROutputS0xD(277)(6);
  CNStageIntLLRInputS1xD(32)(4) <= VNStageIntLLROutputS0xD(278)(0);
  CNStageIntLLRInputS1xD(70)(4) <= VNStageIntLLROutputS0xD(278)(1);
  CNStageIntLLRInputS1xD(141)(4) <= VNStageIntLLROutputS0xD(278)(2);
  CNStageIntLLRInputS1xD(229)(4) <= VNStageIntLLROutputS0xD(278)(3);
  CNStageIntLLRInputS1xD(328)(4) <= VNStageIntLLROutputS0xD(278)(4);
  CNStageIntLLRInputS1xD(31)(4) <= VNStageIntLLROutputS0xD(279)(0);
  CNStageIntLLRInputS1xD(58)(4) <= VNStageIntLLROutputS0xD(279)(1);
  CNStageIntLLRInputS1xD(144)(4) <= VNStageIntLLROutputS0xD(279)(2);
  CNStageIntLLRInputS1xD(219)(4) <= VNStageIntLLROutputS0xD(279)(3);
  CNStageIntLLRInputS1xD(239)(4) <= VNStageIntLLROutputS0xD(279)(4);
  CNStageIntLLRInputS1xD(368)(4) <= VNStageIntLLROutputS0xD(279)(5);
  CNStageIntLLRInputS1xD(30)(4) <= VNStageIntLLROutputS0xD(280)(0);
  CNStageIntLLRInputS1xD(84)(4) <= VNStageIntLLROutputS0xD(280)(1);
  CNStageIntLLRInputS1xD(129)(4) <= VNStageIntLLROutputS0xD(280)(2);
  CNStageIntLLRInputS1xD(215)(4) <= VNStageIntLLROutputS0xD(280)(3);
  CNStageIntLLRInputS1xD(233)(4) <= VNStageIntLLROutputS0xD(280)(4);
  CNStageIntLLRInputS1xD(310)(4) <= VNStageIntLLROutputS0xD(280)(5);
  CNStageIntLLRInputS1xD(376)(4) <= VNStageIntLLROutputS0xD(280)(6);
  CNStageIntLLRInputS1xD(29)(4) <= VNStageIntLLROutputS0xD(281)(0);
  CNStageIntLLRInputS1xD(90)(4) <= VNStageIntLLROutputS0xD(281)(1);
  CNStageIntLLRInputS1xD(163)(4) <= VNStageIntLLROutputS0xD(281)(2);
  CNStageIntLLRInputS1xD(182)(4) <= VNStageIntLLROutputS0xD(281)(3);
  CNStageIntLLRInputS1xD(236)(4) <= VNStageIntLLROutputS0xD(281)(4);
  CNStageIntLLRInputS1xD(298)(4) <= VNStageIntLLROutputS0xD(281)(5);
  CNStageIntLLRInputS1xD(340)(4) <= VNStageIntLLROutputS0xD(281)(6);
  CNStageIntLLRInputS1xD(28)(4) <= VNStageIntLLROutputS0xD(282)(0);
  CNStageIntLLRInputS1xD(74)(4) <= VNStageIntLLROutputS0xD(282)(1);
  CNStageIntLLRInputS1xD(125)(4) <= VNStageIntLLROutputS0xD(282)(2);
  CNStageIntLLRInputS1xD(200)(4) <= VNStageIntLLROutputS0xD(282)(3);
  CNStageIntLLRInputS1xD(226)(4) <= VNStageIntLLROutputS0xD(282)(4);
  CNStageIntLLRInputS1xD(338)(4) <= VNStageIntLLROutputS0xD(282)(5);
  CNStageIntLLRInputS1xD(27)(4) <= VNStageIntLLROutputS0xD(283)(0);
  CNStageIntLLRInputS1xD(76)(4) <= VNStageIntLLROutputS0xD(283)(1);
  CNStageIntLLRInputS1xD(153)(4) <= VNStageIntLLROutputS0xD(283)(2);
  CNStageIntLLRInputS1xD(201)(4) <= VNStageIntLLROutputS0xD(283)(3);
  CNStageIntLLRInputS1xD(260)(4) <= VNStageIntLLROutputS0xD(283)(4);
  CNStageIntLLRInputS1xD(294)(4) <= VNStageIntLLROutputS0xD(283)(5);
  CNStageIntLLRInputS1xD(374)(4) <= VNStageIntLLROutputS0xD(283)(6);
  CNStageIntLLRInputS1xD(26)(4) <= VNStageIntLLROutputS0xD(284)(0);
  CNStageIntLLRInputS1xD(100)(4) <= VNStageIntLLROutputS0xD(284)(1);
  CNStageIntLLRInputS1xD(137)(4) <= VNStageIntLLROutputS0xD(284)(2);
  CNStageIntLLRInputS1xD(181)(4) <= VNStageIntLLROutputS0xD(284)(3);
  CNStageIntLLRInputS1xD(245)(4) <= VNStageIntLLROutputS0xD(284)(4);
  CNStageIntLLRInputS1xD(320)(4) <= VNStageIntLLROutputS0xD(284)(5);
  CNStageIntLLRInputS1xD(353)(4) <= VNStageIntLLROutputS0xD(284)(6);
  CNStageIntLLRInputS1xD(25)(4) <= VNStageIntLLROutputS0xD(285)(0);
  CNStageIntLLRInputS1xD(82)(4) <= VNStageIntLLROutputS0xD(285)(1);
  CNStageIntLLRInputS1xD(165)(4) <= VNStageIntLLROutputS0xD(285)(2);
  CNStageIntLLRInputS1xD(172)(4) <= VNStageIntLLROutputS0xD(285)(3);
  CNStageIntLLRInputS1xD(255)(4) <= VNStageIntLLROutputS0xD(285)(4);
  CNStageIntLLRInputS1xD(304)(4) <= VNStageIntLLROutputS0xD(285)(5);
  CNStageIntLLRInputS1xD(355)(4) <= VNStageIntLLROutputS0xD(285)(6);
  CNStageIntLLRInputS1xD(24)(4) <= VNStageIntLLROutputS0xD(286)(0);
  CNStageIntLLRInputS1xD(93)(4) <= VNStageIntLLROutputS0xD(286)(1);
  CNStageIntLLRInputS1xD(155)(4) <= VNStageIntLLROutputS0xD(286)(2);
  CNStageIntLLRInputS1xD(189)(4) <= VNStageIntLLROutputS0xD(286)(3);
  CNStageIntLLRInputS1xD(267)(4) <= VNStageIntLLROutputS0xD(286)(4);
  CNStageIntLLRInputS1xD(330)(4) <= VNStageIntLLROutputS0xD(286)(5);
  CNStageIntLLRInputS1xD(341)(4) <= VNStageIntLLROutputS0xD(286)(6);
  CNStageIntLLRInputS1xD(23)(4) <= VNStageIntLLROutputS0xD(287)(0);
  CNStageIntLLRInputS1xD(101)(4) <= VNStageIntLLROutputS0xD(287)(1);
  CNStageIntLLRInputS1xD(142)(4) <= VNStageIntLLROutputS0xD(287)(2);
  CNStageIntLLRInputS1xD(193)(4) <= VNStageIntLLROutputS0xD(287)(3);
  CNStageIntLLRInputS1xD(240)(4) <= VNStageIntLLROutputS0xD(287)(4);
  CNStageIntLLRInputS1xD(322)(4) <= VNStageIntLLROutputS0xD(287)(5);
  CNStageIntLLRInputS1xD(375)(4) <= VNStageIntLLROutputS0xD(287)(6);
  CNStageIntLLRInputS1xD(22)(4) <= VNStageIntLLROutputS0xD(288)(0);
  CNStageIntLLRInputS1xD(75)(4) <= VNStageIntLLROutputS0xD(288)(1);
  CNStageIntLLRInputS1xD(161)(4) <= VNStageIntLLROutputS0xD(288)(2);
  CNStageIntLLRInputS1xD(224)(4) <= VNStageIntLLROutputS0xD(288)(3);
  CNStageIntLLRInputS1xD(228)(4) <= VNStageIntLLROutputS0xD(288)(4);
  CNStageIntLLRInputS1xD(308)(4) <= VNStageIntLLROutputS0xD(288)(5);
  CNStageIntLLRInputS1xD(337)(4) <= VNStageIntLLROutputS0xD(288)(6);
  CNStageIntLLRInputS1xD(21)(4) <= VNStageIntLLROutputS0xD(289)(0);
  CNStageIntLLRInputS1xD(89)(4) <= VNStageIntLLROutputS0xD(289)(1);
  CNStageIntLLRInputS1xD(134)(4) <= VNStageIntLLROutputS0xD(289)(2);
  CNStageIntLLRInputS1xD(192)(4) <= VNStageIntLLROutputS0xD(289)(3);
  CNStageIntLLRInputS1xD(269)(4) <= VNStageIntLLROutputS0xD(289)(4);
  CNStageIntLLRInputS1xD(327)(4) <= VNStageIntLLROutputS0xD(289)(5);
  CNStageIntLLRInputS1xD(365)(4) <= VNStageIntLLROutputS0xD(289)(6);
  CNStageIntLLRInputS1xD(20)(4) <= VNStageIntLLROutputS0xD(290)(0);
  CNStageIntLLRInputS1xD(60)(4) <= VNStageIntLLROutputS0xD(290)(1);
  CNStageIntLLRInputS1xD(131)(4) <= VNStageIntLLROutputS0xD(290)(2);
  CNStageIntLLRInputS1xD(187)(4) <= VNStageIntLLROutputS0xD(290)(3);
  CNStageIntLLRInputS1xD(231)(4) <= VNStageIntLLROutputS0xD(290)(4);
  CNStageIntLLRInputS1xD(350)(4) <= VNStageIntLLROutputS0xD(290)(5);
  CNStageIntLLRInputS1xD(19)(4) <= VNStageIntLLROutputS0xD(291)(0);
  CNStageIntLLRInputS1xD(96)(4) <= VNStageIntLLROutputS0xD(291)(1);
  CNStageIntLLRInputS1xD(147)(4) <= VNStageIntLLROutputS0xD(291)(2);
  CNStageIntLLRInputS1xD(223)(4) <= VNStageIntLLROutputS0xD(291)(3);
  CNStageIntLLRInputS1xD(249)(4) <= VNStageIntLLROutputS0xD(291)(4);
  CNStageIntLLRInputS1xD(377)(4) <= VNStageIntLLROutputS0xD(291)(5);
  CNStageIntLLRInputS1xD(18)(4) <= VNStageIntLLROutputS0xD(292)(0);
  CNStageIntLLRInputS1xD(62)(4) <= VNStageIntLLROutputS0xD(292)(1);
  CNStageIntLLRInputS1xD(139)(4) <= VNStageIntLLROutputS0xD(292)(2);
  CNStageIntLLRInputS1xD(177)(4) <= VNStageIntLLROutputS0xD(292)(3);
  CNStageIntLLRInputS1xD(257)(4) <= VNStageIntLLROutputS0xD(292)(4);
  CNStageIntLLRInputS1xD(313)(4) <= VNStageIntLLROutputS0xD(292)(5);
  CNStageIntLLRInputS1xD(367)(4) <= VNStageIntLLROutputS0xD(292)(6);
  CNStageIntLLRInputS1xD(17)(4) <= VNStageIntLLROutputS0xD(293)(0);
  CNStageIntLLRInputS1xD(77)(4) <= VNStageIntLLROutputS0xD(293)(1);
  CNStageIntLLRInputS1xD(113)(4) <= VNStageIntLLROutputS0xD(293)(2);
  CNStageIntLLRInputS1xD(197)(4) <= VNStageIntLLROutputS0xD(293)(3);
  CNStageIntLLRInputS1xD(306)(4) <= VNStageIntLLROutputS0xD(293)(4);
  CNStageIntLLRInputS1xD(354)(4) <= VNStageIntLLROutputS0xD(293)(5);
  CNStageIntLLRInputS1xD(16)(4) <= VNStageIntLLROutputS0xD(294)(0);
  CNStageIntLLRInputS1xD(73)(4) <= VNStageIntLLROutputS0xD(294)(1);
  CNStageIntLLRInputS1xD(123)(4) <= VNStageIntLLROutputS0xD(294)(2);
  CNStageIntLLRInputS1xD(196)(4) <= VNStageIntLLROutputS0xD(294)(3);
  CNStageIntLLRInputS1xD(258)(4) <= VNStageIntLLROutputS0xD(294)(4);
  CNStageIntLLRInputS1xD(284)(4) <= VNStageIntLLROutputS0xD(294)(5);
  CNStageIntLLRInputS1xD(373)(4) <= VNStageIntLLROutputS0xD(294)(6);
  CNStageIntLLRInputS1xD(15)(4) <= VNStageIntLLROutputS0xD(295)(0);
  CNStageIntLLRInputS1xD(92)(4) <= VNStageIntLLROutputS0xD(295)(1);
  CNStageIntLLRInputS1xD(117)(4) <= VNStageIntLLROutputS0xD(295)(2);
  CNStageIntLLRInputS1xD(175)(4) <= VNStageIntLLROutputS0xD(295)(3);
  CNStageIntLLRInputS1xD(346)(4) <= VNStageIntLLROutputS0xD(295)(4);
  CNStageIntLLRInputS1xD(14)(4) <= VNStageIntLLROutputS0xD(296)(0);
  CNStageIntLLRInputS1xD(55)(4) <= VNStageIntLLROutputS0xD(296)(1);
  CNStageIntLLRInputS1xD(121)(4) <= VNStageIntLLROutputS0xD(296)(2);
  CNStageIntLLRInputS1xD(208)(4) <= VNStageIntLLROutputS0xD(296)(3);
  CNStageIntLLRInputS1xD(286)(4) <= VNStageIntLLROutputS0xD(296)(4);
  CNStageIntLLRInputS1xD(343)(4) <= VNStageIntLLROutputS0xD(296)(5);
  CNStageIntLLRInputS1xD(13)(4) <= VNStageIntLLROutputS0xD(297)(0);
  CNStageIntLLRInputS1xD(56)(4) <= VNStageIntLLROutputS0xD(297)(1);
  CNStageIntLLRInputS1xD(111)(4) <= VNStageIntLLROutputS0xD(297)(2);
  CNStageIntLLRInputS1xD(211)(4) <= VNStageIntLLROutputS0xD(297)(3);
  CNStageIntLLRInputS1xD(277)(4) <= VNStageIntLLROutputS0xD(297)(4);
  CNStageIntLLRInputS1xD(290)(4) <= VNStageIntLLROutputS0xD(297)(5);
  CNStageIntLLRInputS1xD(358)(4) <= VNStageIntLLROutputS0xD(297)(6);
  CNStageIntLLRInputS1xD(12)(4) <= VNStageIntLLROutputS0xD(298)(0);
  CNStageIntLLRInputS1xD(91)(4) <= VNStageIntLLROutputS0xD(298)(1);
  CNStageIntLLRInputS1xD(148)(4) <= VNStageIntLLROutputS0xD(298)(2);
  CNStageIntLLRInputS1xD(198)(4) <= VNStageIntLLROutputS0xD(298)(3);
  CNStageIntLLRInputS1xD(262)(4) <= VNStageIntLLROutputS0xD(298)(4);
  CNStageIntLLRInputS1xD(282)(4) <= VNStageIntLLROutputS0xD(298)(5);
  CNStageIntLLRInputS1xD(351)(4) <= VNStageIntLLROutputS0xD(298)(6);
  CNStageIntLLRInputS1xD(83)(4) <= VNStageIntLLROutputS0xD(299)(0);
  CNStageIntLLRInputS1xD(130)(4) <= VNStageIntLLROutputS0xD(299)(1);
  CNStageIntLLRInputS1xD(176)(4) <= VNStageIntLLROutputS0xD(299)(2);
  CNStageIntLLRInputS1xD(264)(4) <= VNStageIntLLROutputS0xD(299)(3);
  CNStageIntLLRInputS1xD(314)(4) <= VNStageIntLLROutputS0xD(299)(4);
  CNStageIntLLRInputS1xD(11)(4) <= VNStageIntLLROutputS0xD(300)(0);
  CNStageIntLLRInputS1xD(99)(4) <= VNStageIntLLROutputS0xD(300)(1);
  CNStageIntLLRInputS1xD(143)(4) <= VNStageIntLLROutputS0xD(300)(2);
  CNStageIntLLRInputS1xD(195)(4) <= VNStageIntLLROutputS0xD(300)(3);
  CNStageIntLLRInputS1xD(299)(4) <= VNStageIntLLROutputS0xD(300)(4);
  CNStageIntLLRInputS1xD(335)(4) <= VNStageIntLLROutputS0xD(300)(5);
  CNStageIntLLRInputS1xD(10)(4) <= VNStageIntLLROutputS0xD(301)(0);
  CNStageIntLLRInputS1xD(103)(4) <= VNStageIntLLROutputS0xD(301)(1);
  CNStageIntLLRInputS1xD(154)(4) <= VNStageIntLLROutputS0xD(301)(2);
  CNStageIntLLRInputS1xD(220)(4) <= VNStageIntLLROutputS0xD(301)(3);
  CNStageIntLLRInputS1xD(270)(4) <= VNStageIntLLROutputS0xD(301)(4);
  CNStageIntLLRInputS1xD(309)(4) <= VNStageIntLLROutputS0xD(301)(5);
  CNStageIntLLRInputS1xD(9)(4) <= VNStageIntLLROutputS0xD(302)(0);
  CNStageIntLLRInputS1xD(110)(4) <= VNStageIntLLROutputS0xD(302)(1);
  CNStageIntLLRInputS1xD(124)(4) <= VNStageIntLLROutputS0xD(302)(2);
  CNStageIntLLRInputS1xD(206)(4) <= VNStageIntLLROutputS0xD(302)(3);
  CNStageIntLLRInputS1xD(227)(4) <= VNStageIntLLROutputS0xD(302)(4);
  CNStageIntLLRInputS1xD(321)(4) <= VNStageIntLLROutputS0xD(302)(5);
  CNStageIntLLRInputS1xD(8)(4) <= VNStageIntLLROutputS0xD(303)(0);
  CNStageIntLLRInputS1xD(102)(4) <= VNStageIntLLROutputS0xD(303)(1);
  CNStageIntLLRInputS1xD(112)(4) <= VNStageIntLLROutputS0xD(303)(2);
  CNStageIntLLRInputS1xD(178)(4) <= VNStageIntLLROutputS0xD(303)(3);
  CNStageIntLLRInputS1xD(235)(4) <= VNStageIntLLROutputS0xD(303)(4);
  CNStageIntLLRInputS1xD(293)(4) <= VNStageIntLLROutputS0xD(303)(5);
  CNStageIntLLRInputS1xD(382)(4) <= VNStageIntLLROutputS0xD(303)(6);
  CNStageIntLLRInputS1xD(7)(4) <= VNStageIntLLROutputS0xD(304)(0);
  CNStageIntLLRInputS1xD(97)(4) <= VNStageIntLLROutputS0xD(304)(1);
  CNStageIntLLRInputS1xD(157)(4) <= VNStageIntLLROutputS0xD(304)(2);
  CNStageIntLLRInputS1xD(222)(4) <= VNStageIntLLROutputS0xD(304)(3);
  CNStageIntLLRInputS1xD(263)(4) <= VNStageIntLLROutputS0xD(304)(4);
  CNStageIntLLRInputS1xD(283)(4) <= VNStageIntLLROutputS0xD(304)(5);
  CNStageIntLLRInputS1xD(359)(4) <= VNStageIntLLROutputS0xD(304)(6);
  CNStageIntLLRInputS1xD(6)(4) <= VNStageIntLLROutputS0xD(305)(0);
  CNStageIntLLRInputS1xD(80)(4) <= VNStageIntLLROutputS0xD(305)(1);
  CNStageIntLLRInputS1xD(115)(4) <= VNStageIntLLROutputS0xD(305)(2);
  CNStageIntLLRInputS1xD(209)(4) <= VNStageIntLLROutputS0xD(305)(3);
  CNStageIntLLRInputS1xD(276)(4) <= VNStageIntLLROutputS0xD(305)(4);
  CNStageIntLLRInputS1xD(323)(4) <= VNStageIntLLROutputS0xD(305)(5);
  CNStageIntLLRInputS1xD(342)(4) <= VNStageIntLLROutputS0xD(305)(6);
  CNStageIntLLRInputS1xD(5)(4) <= VNStageIntLLROutputS0xD(306)(0);
  CNStageIntLLRInputS1xD(87)(4) <= VNStageIntLLROutputS0xD(306)(1);
  CNStageIntLLRInputS1xD(136)(4) <= VNStageIntLLROutputS0xD(306)(2);
  CNStageIntLLRInputS1xD(174)(4) <= VNStageIntLLROutputS0xD(306)(3);
  CNStageIntLLRInputS1xD(4)(4) <= VNStageIntLLROutputS0xD(307)(0);
  CNStageIntLLRInputS1xD(107)(4) <= VNStageIntLLROutputS0xD(307)(1);
  CNStageIntLLRInputS1xD(145)(4) <= VNStageIntLLROutputS0xD(307)(2);
  CNStageIntLLRInputS1xD(202)(4) <= VNStageIntLLROutputS0xD(307)(3);
  CNStageIntLLRInputS1xD(230)(4) <= VNStageIntLLROutputS0xD(307)(4);
  CNStageIntLLRInputS1xD(302)(4) <= VNStageIntLLROutputS0xD(307)(5);
  CNStageIntLLRInputS1xD(366)(4) <= VNStageIntLLROutputS0xD(307)(6);
  CNStageIntLLRInputS1xD(140)(4) <= VNStageIntLLROutputS0xD(308)(0);
  CNStageIntLLRInputS1xD(199)(4) <= VNStageIntLLROutputS0xD(308)(1);
  CNStageIntLLRInputS1xD(251)(4) <= VNStageIntLLROutputS0xD(308)(2);
  CNStageIntLLRInputS1xD(311)(4) <= VNStageIntLLROutputS0xD(308)(3);
  CNStageIntLLRInputS1xD(336)(4) <= VNStageIntLLROutputS0xD(308)(4);
  CNStageIntLLRInputS1xD(3)(4) <= VNStageIntLLROutputS0xD(309)(0);
  CNStageIntLLRInputS1xD(86)(4) <= VNStageIntLLROutputS0xD(309)(1);
  CNStageIntLLRInputS1xD(146)(4) <= VNStageIntLLROutputS0xD(309)(2);
  CNStageIntLLRInputS1xD(214)(4) <= VNStageIntLLROutputS0xD(309)(3);
  CNStageIntLLRInputS1xD(265)(4) <= VNStageIntLLROutputS0xD(309)(4);
  CNStageIntLLRInputS1xD(307)(4) <= VNStageIntLLROutputS0xD(309)(5);
  CNStageIntLLRInputS1xD(2)(4) <= VNStageIntLLROutputS0xD(310)(0);
  CNStageIntLLRInputS1xD(65)(4) <= VNStageIntLLROutputS0xD(310)(1);
  CNStageIntLLRInputS1xD(135)(4) <= VNStageIntLLROutputS0xD(310)(2);
  CNStageIntLLRInputS1xD(261)(4) <= VNStageIntLLROutputS0xD(310)(3);
  CNStageIntLLRInputS1xD(312)(4) <= VNStageIntLLROutputS0xD(310)(4);
  CNStageIntLLRInputS1xD(369)(4) <= VNStageIntLLROutputS0xD(310)(5);
  CNStageIntLLRInputS1xD(1)(4) <= VNStageIntLLROutputS0xD(311)(0);
  CNStageIntLLRInputS1xD(68)(4) <= VNStageIntLLROutputS0xD(311)(1);
  CNStageIntLLRInputS1xD(160)(4) <= VNStageIntLLROutputS0xD(311)(2);
  CNStageIntLLRInputS1xD(225)(4) <= VNStageIntLLROutputS0xD(311)(3);
  CNStageIntLLRInputS1xD(301)(4) <= VNStageIntLLROutputS0xD(311)(4);
  CNStageIntLLRInputS1xD(0)(4) <= VNStageIntLLROutputS0xD(312)(0);
  CNStageIntLLRInputS1xD(108)(4) <= VNStageIntLLROutputS0xD(312)(1);
  CNStageIntLLRInputS1xD(167)(4) <= VNStageIntLLROutputS0xD(312)(2);
  CNStageIntLLRInputS1xD(246)(4) <= VNStageIntLLROutputS0xD(312)(3);
  CNStageIntLLRInputS1xD(326)(4) <= VNStageIntLLROutputS0xD(312)(4);
  CNStageIntLLRInputS1xD(348)(4) <= VNStageIntLLROutputS0xD(312)(5);
  CNStageIntLLRInputS1xD(150)(4) <= VNStageIntLLROutputS0xD(313)(0);
  CNStageIntLLRInputS1xD(188)(4) <= VNStageIntLLROutputS0xD(313)(1);
  CNStageIntLLRInputS1xD(247)(4) <= VNStageIntLLROutputS0xD(313)(2);
  CNStageIntLLRInputS1xD(356)(4) <= VNStageIntLLROutputS0xD(313)(3);
  CNStageIntLLRInputS1xD(191)(4) <= VNStageIntLLROutputS0xD(314)(0);
  CNStageIntLLRInputS1xD(278)(4) <= VNStageIntLLROutputS0xD(314)(1);
  CNStageIntLLRInputS1xD(316)(4) <= VNStageIntLLROutputS0xD(314)(2);
  CNStageIntLLRInputS1xD(352)(4) <= VNStageIntLLROutputS0xD(314)(3);
  CNStageIntLLRInputS1xD(78)(4) <= VNStageIntLLROutputS0xD(315)(0);
  CNStageIntLLRInputS1xD(119)(4) <= VNStageIntLLROutputS0xD(315)(1);
  CNStageIntLLRInputS1xD(183)(4) <= VNStageIntLLROutputS0xD(315)(2);
  CNStageIntLLRInputS1xD(271)(4) <= VNStageIntLLROutputS0xD(315)(3);
  CNStageIntLLRInputS1xD(318)(4) <= VNStageIntLLROutputS0xD(315)(4);
  CNStageIntLLRInputS1xD(357)(4) <= VNStageIntLLROutputS0xD(315)(5);
  CNStageIntLLRInputS1xD(61)(4) <= VNStageIntLLROutputS0xD(316)(0);
  CNStageIntLLRInputS1xD(158)(4) <= VNStageIntLLROutputS0xD(316)(1);
  CNStageIntLLRInputS1xD(234)(4) <= VNStageIntLLROutputS0xD(316)(2);
  CNStageIntLLRInputS1xD(288)(4) <= VNStageIntLLROutputS0xD(316)(3);
  CNStageIntLLRInputS1xD(347)(4) <= VNStageIntLLROutputS0xD(316)(4);
  CNStageIntLLRInputS1xD(88)(4) <= VNStageIntLLROutputS0xD(317)(0);
  CNStageIntLLRInputS1xD(238)(4) <= VNStageIntLLROutputS0xD(317)(1);
  CNStageIntLLRInputS1xD(324)(4) <= VNStageIntLLROutputS0xD(317)(2);
  CNStageIntLLRInputS1xD(372)(4) <= VNStageIntLLROutputS0xD(317)(3);
  CNStageIntLLRInputS1xD(120)(4) <= VNStageIntLLROutputS0xD(318)(0);
  CNStageIntLLRInputS1xD(210)(4) <= VNStageIntLLROutputS0xD(318)(1);
  CNStageIntLLRInputS1xD(279)(4) <= VNStageIntLLROutputS0xD(318)(2);
  CNStageIntLLRInputS1xD(379)(4) <= VNStageIntLLROutputS0xD(318)(3);
  CNStageIntLLRInputS1xD(52)(4) <= VNStageIntLLROutputS0xD(319)(0);
  CNStageIntLLRInputS1xD(66)(4) <= VNStageIntLLROutputS0xD(319)(1);
  CNStageIntLLRInputS1xD(151)(4) <= VNStageIntLLROutputS0xD(319)(2);
  CNStageIntLLRInputS1xD(221)(4) <= VNStageIntLLROutputS0xD(319)(3);
  CNStageIntLLRInputS1xD(237)(4) <= VNStageIntLLROutputS0xD(319)(4);
  CNStageIntLLRInputS1xD(289)(4) <= VNStageIntLLROutputS0xD(319)(5);
  CNStageIntLLRInputS1xD(361)(4) <= VNStageIntLLROutputS0xD(319)(6);
  CNStageIntLLRInputS1xD(53)(5) <= VNStageIntLLROutputS0xD(320)(0);
  CNStageIntLLRInputS1xD(126)(5) <= VNStageIntLLROutputS0xD(320)(1);
  CNStageIntLLRInputS1xD(196)(5) <= VNStageIntLLROutputS0xD(320)(2);
  CNStageIntLLRInputS1xD(295)(5) <= VNStageIntLLROutputS0xD(320)(3);
  CNStageIntLLRInputS1xD(338)(5) <= VNStageIntLLROutputS0xD(320)(4);
  CNStageIntLLRInputS1xD(51)(5) <= VNStageIntLLROutputS0xD(321)(0);
  CNStageIntLLRInputS1xD(65)(5) <= VNStageIntLLROutputS0xD(321)(1);
  CNStageIntLLRInputS1xD(150)(5) <= VNStageIntLLROutputS0xD(321)(2);
  CNStageIntLLRInputS1xD(220)(5) <= VNStageIntLLROutputS0xD(321)(3);
  CNStageIntLLRInputS1xD(236)(5) <= VNStageIntLLROutputS0xD(321)(4);
  CNStageIntLLRInputS1xD(288)(5) <= VNStageIntLLROutputS0xD(321)(5);
  CNStageIntLLRInputS1xD(360)(5) <= VNStageIntLLROutputS0xD(321)(6);
  CNStageIntLLRInputS1xD(50)(5) <= VNStageIntLLROutputS0xD(322)(0);
  CNStageIntLLRInputS1xD(84)(5) <= VNStageIntLLROutputS0xD(322)(1);
  CNStageIntLLRInputS1xD(165)(5) <= VNStageIntLLROutputS0xD(322)(2);
  CNStageIntLLRInputS1xD(231)(5) <= VNStageIntLLROutputS0xD(322)(3);
  CNStageIntLLRInputS1xD(316)(5) <= VNStageIntLLROutputS0xD(322)(4);
  CNStageIntLLRInputS1xD(362)(5) <= VNStageIntLLROutputS0xD(322)(5);
  CNStageIntLLRInputS1xD(56)(5) <= VNStageIntLLROutputS0xD(323)(0);
  CNStageIntLLRInputS1xD(136)(5) <= VNStageIntLLROutputS0xD(323)(1);
  CNStageIntLLRInputS1xD(184)(5) <= VNStageIntLLROutputS0xD(323)(2);
  CNStageIntLLRInputS1xD(268)(5) <= VNStageIntLLROutputS0xD(323)(3);
  CNStageIntLLRInputS1xD(330)(5) <= VNStageIntLLROutputS0xD(323)(4);
  CNStageIntLLRInputS1xD(49)(5) <= VNStageIntLLROutputS0xD(324)(0);
  CNStageIntLLRInputS1xD(109)(5) <= VNStageIntLLROutputS0xD(324)(1);
  CNStageIntLLRInputS1xD(113)(5) <= VNStageIntLLROutputS0xD(324)(2);
  CNStageIntLLRInputS1xD(223)(5) <= VNStageIntLLROutputS0xD(324)(3);
  CNStageIntLLRInputS1xD(273)(5) <= VNStageIntLLROutputS0xD(324)(4);
  CNStageIntLLRInputS1xD(302)(5) <= VNStageIntLLROutputS0xD(324)(5);
  CNStageIntLLRInputS1xD(369)(5) <= VNStageIntLLROutputS0xD(324)(6);
  CNStageIntLLRInputS1xD(48)(5) <= VNStageIntLLROutputS0xD(325)(0);
  CNStageIntLLRInputS1xD(70)(5) <= VNStageIntLLROutputS0xD(325)(1);
  CNStageIntLLRInputS1xD(137)(5) <= VNStageIntLLROutputS0xD(325)(2);
  CNStageIntLLRInputS1xD(185)(5) <= VNStageIntLLROutputS0xD(325)(3);
  CNStageIntLLRInputS1xD(242)(5) <= VNStageIntLLROutputS0xD(325)(4);
  CNStageIntLLRInputS1xD(284)(5) <= VNStageIntLLROutputS0xD(325)(5);
  CNStageIntLLRInputS1xD(382)(5) <= VNStageIntLLROutputS0xD(325)(6);
  CNStageIntLLRInputS1xD(47)(5) <= VNStageIntLLROutputS0xD(326)(0);
  CNStageIntLLRInputS1xD(62)(5) <= VNStageIntLLROutputS0xD(326)(1);
  CNStageIntLLRInputS1xD(203)(5) <= VNStageIntLLROutputS0xD(326)(2);
  CNStageIntLLRInputS1xD(241)(5) <= VNStageIntLLROutputS0xD(326)(3);
  CNStageIntLLRInputS1xD(304)(5) <= VNStageIntLLROutputS0xD(326)(4);
  CNStageIntLLRInputS1xD(46)(5) <= VNStageIntLLROutputS0xD(327)(0);
  CNStageIntLLRInputS1xD(94)(5) <= VNStageIntLLROutputS0xD(327)(1);
  CNStageIntLLRInputS1xD(148)(5) <= VNStageIntLLROutputS0xD(327)(2);
  CNStageIntLLRInputS1xD(211)(5) <= VNStageIntLLROutputS0xD(327)(3);
  CNStageIntLLRInputS1xD(272)(5) <= VNStageIntLLROutputS0xD(327)(4);
  CNStageIntLLRInputS1xD(318)(5) <= VNStageIntLLROutputS0xD(327)(5);
  CNStageIntLLRInputS1xD(361)(5) <= VNStageIntLLROutputS0xD(327)(6);
  CNStageIntLLRInputS1xD(45)(5) <= VNStageIntLLROutputS0xD(328)(0);
  CNStageIntLLRInputS1xD(103)(5) <= VNStageIntLLROutputS0xD(328)(1);
  CNStageIntLLRInputS1xD(168)(5) <= VNStageIntLLROutputS0xD(328)(2);
  CNStageIntLLRInputS1xD(314)(5) <= VNStageIntLLROutputS0xD(328)(3);
  CNStageIntLLRInputS1xD(377)(5) <= VNStageIntLLROutputS0xD(328)(4);
  CNStageIntLLRInputS1xD(44)(5) <= VNStageIntLLROutputS0xD(329)(0);
  CNStageIntLLRInputS1xD(97)(5) <= VNStageIntLLROutputS0xD(329)(1);
  CNStageIntLLRInputS1xD(131)(5) <= VNStageIntLLROutputS0xD(329)(2);
  CNStageIntLLRInputS1xD(212)(5) <= VNStageIntLLROutputS0xD(329)(3);
  CNStageIntLLRInputS1xD(255)(5) <= VNStageIntLLROutputS0xD(329)(4);
  CNStageIntLLRInputS1xD(280)(5) <= VNStageIntLLROutputS0xD(329)(5);
  CNStageIntLLRInputS1xD(348)(5) <= VNStageIntLLROutputS0xD(329)(6);
  CNStageIntLLRInputS1xD(43)(5) <= VNStageIntLLROutputS0xD(330)(0);
  CNStageIntLLRInputS1xD(101)(5) <= VNStageIntLLROutputS0xD(330)(1);
  CNStageIntLLRInputS1xD(132)(5) <= VNStageIntLLROutputS0xD(330)(2);
  CNStageIntLLRInputS1xD(202)(5) <= VNStageIntLLROutputS0xD(330)(3);
  CNStageIntLLRInputS1xD(243)(5) <= VNStageIntLLROutputS0xD(330)(4);
  CNStageIntLLRInputS1xD(42)(5) <= VNStageIntLLROutputS0xD(331)(0);
  CNStageIntLLRInputS1xD(92)(5) <= VNStageIntLLROutputS0xD(331)(1);
  CNStageIntLLRInputS1xD(167)(5) <= VNStageIntLLROutputS0xD(331)(2);
  CNStageIntLLRInputS1xD(172)(5) <= VNStageIntLLROutputS0xD(331)(3);
  CNStageIntLLRInputS1xD(350)(5) <= VNStageIntLLROutputS0xD(331)(4);
  CNStageIntLLRInputS1xD(41)(5) <= VNStageIntLLROutputS0xD(332)(0);
  CNStageIntLLRInputS1xD(71)(5) <= VNStageIntLLROutputS0xD(332)(1);
  CNStageIntLLRInputS1xD(158)(5) <= VNStageIntLLROutputS0xD(332)(2);
  CNStageIntLLRInputS1xD(179)(5) <= VNStageIntLLROutputS0xD(332)(3);
  CNStageIntLLRInputS1xD(240)(5) <= VNStageIntLLROutputS0xD(332)(4);
  CNStageIntLLRInputS1xD(363)(5) <= VNStageIntLLROutputS0xD(332)(5);
  CNStageIntLLRInputS1xD(108)(5) <= VNStageIntLLROutputS0xD(333)(0);
  CNStageIntLLRInputS1xD(117)(5) <= VNStageIntLLROutputS0xD(333)(1);
  CNStageIntLLRInputS1xD(215)(5) <= VNStageIntLLROutputS0xD(333)(2);
  CNStageIntLLRInputS1xD(265)(5) <= VNStageIntLLROutputS0xD(333)(3);
  CNStageIntLLRInputS1xD(324)(5) <= VNStageIntLLROutputS0xD(333)(4);
  CNStageIntLLRInputS1xD(359)(5) <= VNStageIntLLROutputS0xD(333)(5);
  CNStageIntLLRInputS1xD(40)(5) <= VNStageIntLLROutputS0xD(334)(0);
  CNStageIntLLRInputS1xD(66)(5) <= VNStageIntLLROutputS0xD(334)(1);
  CNStageIntLLRInputS1xD(217)(5) <= VNStageIntLLROutputS0xD(334)(2);
  CNStageIntLLRInputS1xD(286)(5) <= VNStageIntLLROutputS0xD(334)(3);
  CNStageIntLLRInputS1xD(380)(5) <= VNStageIntLLROutputS0xD(334)(4);
  CNStageIntLLRInputS1xD(39)(5) <= VNStageIntLLROutputS0xD(335)(0);
  CNStageIntLLRInputS1xD(78)(5) <= VNStageIntLLROutputS0xD(335)(1);
  CNStageIntLLRInputS1xD(170)(5) <= VNStageIntLLROutputS0xD(335)(2);
  CNStageIntLLRInputS1xD(189)(5) <= VNStageIntLLROutputS0xD(335)(3);
  CNStageIntLLRInputS1xD(274)(5) <= VNStageIntLLROutputS0xD(335)(4);
  CNStageIntLLRInputS1xD(291)(5) <= VNStageIntLLROutputS0xD(335)(5);
  CNStageIntLLRInputS1xD(343)(5) <= VNStageIntLLROutputS0xD(335)(6);
  CNStageIntLLRInputS1xD(38)(5) <= VNStageIntLLROutputS0xD(336)(0);
  CNStageIntLLRInputS1xD(104)(5) <= VNStageIntLLROutputS0xD(336)(1);
  CNStageIntLLRInputS1xD(121)(5) <= VNStageIntLLROutputS0xD(336)(2);
  CNStageIntLLRInputS1xD(267)(5) <= VNStageIntLLROutputS0xD(336)(3);
  CNStageIntLLRInputS1xD(332)(5) <= VNStageIntLLROutputS0xD(336)(4);
  CNStageIntLLRInputS1xD(344)(5) <= VNStageIntLLROutputS0xD(336)(5);
  CNStageIntLLRInputS1xD(37)(5) <= VNStageIntLLROutputS0xD(337)(0);
  CNStageIntLLRInputS1xD(93)(5) <= VNStageIntLLROutputS0xD(337)(1);
  CNStageIntLLRInputS1xD(115)(5) <= VNStageIntLLROutputS0xD(337)(2);
  CNStageIntLLRInputS1xD(183)(5) <= VNStageIntLLROutputS0xD(337)(3);
  CNStageIntLLRInputS1xD(253)(5) <= VNStageIntLLROutputS0xD(337)(4);
  CNStageIntLLRInputS1xD(290)(5) <= VNStageIntLLROutputS0xD(337)(5);
  CNStageIntLLRInputS1xD(379)(5) <= VNStageIntLLROutputS0xD(337)(6);
  CNStageIntLLRInputS1xD(36)(5) <= VNStageIntLLROutputS0xD(338)(0);
  CNStageIntLLRInputS1xD(80)(5) <= VNStageIntLLROutputS0xD(338)(1);
  CNStageIntLLRInputS1xD(155)(5) <= VNStageIntLLROutputS0xD(338)(2);
  CNStageIntLLRInputS1xD(190)(5) <= VNStageIntLLROutputS0xD(338)(3);
  CNStageIntLLRInputS1xD(370)(5) <= VNStageIntLLROutputS0xD(338)(4);
  CNStageIntLLRInputS1xD(35)(5) <= VNStageIntLLROutputS0xD(339)(0);
  CNStageIntLLRInputS1xD(96)(5) <= VNStageIntLLROutputS0xD(339)(1);
  CNStageIntLLRInputS1xD(163)(5) <= VNStageIntLLROutputS0xD(339)(2);
  CNStageIntLLRInputS1xD(216)(5) <= VNStageIntLLROutputS0xD(339)(3);
  CNStageIntLLRInputS1xD(247)(5) <= VNStageIntLLROutputS0xD(339)(4);
  CNStageIntLLRInputS1xD(322)(5) <= VNStageIntLLROutputS0xD(339)(5);
  CNStageIntLLRInputS1xD(34)(5) <= VNStageIntLLROutputS0xD(340)(0);
  CNStageIntLLRInputS1xD(58)(5) <= VNStageIntLLROutputS0xD(340)(1);
  CNStageIntLLRInputS1xD(127)(5) <= VNStageIntLLROutputS0xD(340)(2);
  CNStageIntLLRInputS1xD(178)(5) <= VNStageIntLLROutputS0xD(340)(3);
  CNStageIntLLRInputS1xD(245)(5) <= VNStageIntLLROutputS0xD(340)(4);
  CNStageIntLLRInputS1xD(334)(5) <= VNStageIntLLROutputS0xD(340)(5);
  CNStageIntLLRInputS1xD(33)(5) <= VNStageIntLLROutputS0xD(341)(0);
  CNStageIntLLRInputS1xD(68)(5) <= VNStageIntLLROutputS0xD(341)(1);
  CNStageIntLLRInputS1xD(125)(5) <= VNStageIntLLROutputS0xD(341)(2);
  CNStageIntLLRInputS1xD(204)(5) <= VNStageIntLLROutputS0xD(341)(3);
  CNStageIntLLRInputS1xD(258)(5) <= VNStageIntLLROutputS0xD(341)(4);
  CNStageIntLLRInputS1xD(296)(5) <= VNStageIntLLROutputS0xD(341)(5);
  CNStageIntLLRInputS1xD(32)(5) <= VNStageIntLLROutputS0xD(342)(0);
  CNStageIntLLRInputS1xD(63)(5) <= VNStageIntLLROutputS0xD(342)(1);
  CNStageIntLLRInputS1xD(161)(5) <= VNStageIntLLROutputS0xD(342)(2);
  CNStageIntLLRInputS1xD(251)(5) <= VNStageIntLLROutputS0xD(342)(3);
  CNStageIntLLRInputS1xD(294)(5) <= VNStageIntLLROutputS0xD(342)(4);
  CNStageIntLLRInputS1xD(31)(5) <= VNStageIntLLROutputS0xD(343)(0);
  CNStageIntLLRInputS1xD(69)(5) <= VNStageIntLLROutputS0xD(343)(1);
  CNStageIntLLRInputS1xD(140)(5) <= VNStageIntLLROutputS0xD(343)(2);
  CNStageIntLLRInputS1xD(206)(5) <= VNStageIntLLROutputS0xD(343)(3);
  CNStageIntLLRInputS1xD(228)(5) <= VNStageIntLLROutputS0xD(343)(4);
  CNStageIntLLRInputS1xD(327)(5) <= VNStageIntLLROutputS0xD(343)(5);
  CNStageIntLLRInputS1xD(30)(5) <= VNStageIntLLROutputS0xD(344)(0);
  CNStageIntLLRInputS1xD(57)(5) <= VNStageIntLLROutputS0xD(344)(1);
  CNStageIntLLRInputS1xD(143)(5) <= VNStageIntLLROutputS0xD(344)(2);
  CNStageIntLLRInputS1xD(218)(5) <= VNStageIntLLROutputS0xD(344)(3);
  CNStageIntLLRInputS1xD(238)(5) <= VNStageIntLLROutputS0xD(344)(4);
  CNStageIntLLRInputS1xD(307)(5) <= VNStageIntLLROutputS0xD(344)(5);
  CNStageIntLLRInputS1xD(367)(5) <= VNStageIntLLROutputS0xD(344)(6);
  CNStageIntLLRInputS1xD(29)(5) <= VNStageIntLLROutputS0xD(345)(0);
  CNStageIntLLRInputS1xD(83)(5) <= VNStageIntLLROutputS0xD(345)(1);
  CNStageIntLLRInputS1xD(128)(5) <= VNStageIntLLROutputS0xD(345)(2);
  CNStageIntLLRInputS1xD(232)(5) <= VNStageIntLLROutputS0xD(345)(3);
  CNStageIntLLRInputS1xD(309)(5) <= VNStageIntLLROutputS0xD(345)(4);
  CNStageIntLLRInputS1xD(375)(5) <= VNStageIntLLROutputS0xD(345)(5);
  CNStageIntLLRInputS1xD(28)(5) <= VNStageIntLLROutputS0xD(346)(0);
  CNStageIntLLRInputS1xD(89)(5) <= VNStageIntLLROutputS0xD(346)(1);
  CNStageIntLLRInputS1xD(162)(5) <= VNStageIntLLROutputS0xD(346)(2);
  CNStageIntLLRInputS1xD(181)(5) <= VNStageIntLLROutputS0xD(346)(3);
  CNStageIntLLRInputS1xD(235)(5) <= VNStageIntLLROutputS0xD(346)(4);
  CNStageIntLLRInputS1xD(297)(5) <= VNStageIntLLROutputS0xD(346)(5);
  CNStageIntLLRInputS1xD(339)(5) <= VNStageIntLLROutputS0xD(346)(6);
  CNStageIntLLRInputS1xD(27)(5) <= VNStageIntLLROutputS0xD(347)(0);
  CNStageIntLLRInputS1xD(73)(5) <= VNStageIntLLROutputS0xD(347)(1);
  CNStageIntLLRInputS1xD(124)(5) <= VNStageIntLLROutputS0xD(347)(2);
  CNStageIntLLRInputS1xD(199)(5) <= VNStageIntLLROutputS0xD(347)(3);
  CNStageIntLLRInputS1xD(225)(5) <= VNStageIntLLROutputS0xD(347)(4);
  CNStageIntLLRInputS1xD(328)(5) <= VNStageIntLLROutputS0xD(347)(5);
  CNStageIntLLRInputS1xD(337)(5) <= VNStageIntLLROutputS0xD(347)(6);
  CNStageIntLLRInputS1xD(26)(5) <= VNStageIntLLROutputS0xD(348)(0);
  CNStageIntLLRInputS1xD(75)(5) <= VNStageIntLLROutputS0xD(348)(1);
  CNStageIntLLRInputS1xD(152)(5) <= VNStageIntLLROutputS0xD(348)(2);
  CNStageIntLLRInputS1xD(200)(5) <= VNStageIntLLROutputS0xD(348)(3);
  CNStageIntLLRInputS1xD(259)(5) <= VNStageIntLLROutputS0xD(348)(4);
  CNStageIntLLRInputS1xD(293)(5) <= VNStageIntLLROutputS0xD(348)(5);
  CNStageIntLLRInputS1xD(373)(5) <= VNStageIntLLROutputS0xD(348)(6);
  CNStageIntLLRInputS1xD(25)(5) <= VNStageIntLLROutputS0xD(349)(0);
  CNStageIntLLRInputS1xD(99)(5) <= VNStageIntLLROutputS0xD(349)(1);
  CNStageIntLLRInputS1xD(180)(5) <= VNStageIntLLROutputS0xD(349)(2);
  CNStageIntLLRInputS1xD(244)(5) <= VNStageIntLLROutputS0xD(349)(3);
  CNStageIntLLRInputS1xD(319)(5) <= VNStageIntLLROutputS0xD(349)(4);
  CNStageIntLLRInputS1xD(352)(5) <= VNStageIntLLROutputS0xD(349)(5);
  CNStageIntLLRInputS1xD(24)(5) <= VNStageIntLLROutputS0xD(350)(0);
  CNStageIntLLRInputS1xD(81)(5) <= VNStageIntLLROutputS0xD(350)(1);
  CNStageIntLLRInputS1xD(164)(5) <= VNStageIntLLROutputS0xD(350)(2);
  CNStageIntLLRInputS1xD(171)(5) <= VNStageIntLLROutputS0xD(350)(3);
  CNStageIntLLRInputS1xD(254)(5) <= VNStageIntLLROutputS0xD(350)(4);
  CNStageIntLLRInputS1xD(303)(5) <= VNStageIntLLROutputS0xD(350)(5);
  CNStageIntLLRInputS1xD(23)(5) <= VNStageIntLLROutputS0xD(351)(0);
  CNStageIntLLRInputS1xD(154)(5) <= VNStageIntLLROutputS0xD(351)(1);
  CNStageIntLLRInputS1xD(188)(5) <= VNStageIntLLROutputS0xD(351)(2);
  CNStageIntLLRInputS1xD(266)(5) <= VNStageIntLLROutputS0xD(351)(3);
  CNStageIntLLRInputS1xD(329)(5) <= VNStageIntLLROutputS0xD(351)(4);
  CNStageIntLLRInputS1xD(340)(5) <= VNStageIntLLROutputS0xD(351)(5);
  CNStageIntLLRInputS1xD(22)(5) <= VNStageIntLLROutputS0xD(352)(0);
  CNStageIntLLRInputS1xD(100)(5) <= VNStageIntLLROutputS0xD(352)(1);
  CNStageIntLLRInputS1xD(141)(5) <= VNStageIntLLROutputS0xD(352)(2);
  CNStageIntLLRInputS1xD(192)(5) <= VNStageIntLLROutputS0xD(352)(3);
  CNStageIntLLRInputS1xD(239)(5) <= VNStageIntLLROutputS0xD(352)(4);
  CNStageIntLLRInputS1xD(321)(5) <= VNStageIntLLROutputS0xD(352)(5);
  CNStageIntLLRInputS1xD(374)(5) <= VNStageIntLLROutputS0xD(352)(6);
  CNStageIntLLRInputS1xD(21)(5) <= VNStageIntLLROutputS0xD(353)(0);
  CNStageIntLLRInputS1xD(74)(5) <= VNStageIntLLROutputS0xD(353)(1);
  CNStageIntLLRInputS1xD(160)(5) <= VNStageIntLLROutputS0xD(353)(2);
  CNStageIntLLRInputS1xD(224)(5) <= VNStageIntLLROutputS0xD(353)(3);
  CNStageIntLLRInputS1xD(227)(5) <= VNStageIntLLROutputS0xD(353)(4);
  CNStageIntLLRInputS1xD(336)(5) <= VNStageIntLLROutputS0xD(353)(5);
  CNStageIntLLRInputS1xD(20)(5) <= VNStageIntLLROutputS0xD(354)(0);
  CNStageIntLLRInputS1xD(88)(5) <= VNStageIntLLROutputS0xD(354)(1);
  CNStageIntLLRInputS1xD(133)(5) <= VNStageIntLLROutputS0xD(354)(2);
  CNStageIntLLRInputS1xD(191)(5) <= VNStageIntLLROutputS0xD(354)(3);
  CNStageIntLLRInputS1xD(326)(5) <= VNStageIntLLROutputS0xD(354)(4);
  CNStageIntLLRInputS1xD(364)(5) <= VNStageIntLLROutputS0xD(354)(5);
  CNStageIntLLRInputS1xD(19)(5) <= VNStageIntLLROutputS0xD(355)(0);
  CNStageIntLLRInputS1xD(59)(5) <= VNStageIntLLROutputS0xD(355)(1);
  CNStageIntLLRInputS1xD(130)(5) <= VNStageIntLLROutputS0xD(355)(2);
  CNStageIntLLRInputS1xD(186)(5) <= VNStageIntLLROutputS0xD(355)(3);
  CNStageIntLLRInputS1xD(230)(5) <= VNStageIntLLROutputS0xD(355)(4);
  CNStageIntLLRInputS1xD(300)(5) <= VNStageIntLLROutputS0xD(355)(5);
  CNStageIntLLRInputS1xD(349)(5) <= VNStageIntLLROutputS0xD(355)(6);
  CNStageIntLLRInputS1xD(18)(5) <= VNStageIntLLROutputS0xD(356)(0);
  CNStageIntLLRInputS1xD(95)(5) <= VNStageIntLLROutputS0xD(356)(1);
  CNStageIntLLRInputS1xD(146)(5) <= VNStageIntLLROutputS0xD(356)(2);
  CNStageIntLLRInputS1xD(222)(5) <= VNStageIntLLROutputS0xD(356)(3);
  CNStageIntLLRInputS1xD(299)(5) <= VNStageIntLLROutputS0xD(356)(4);
  CNStageIntLLRInputS1xD(376)(5) <= VNStageIntLLROutputS0xD(356)(5);
  CNStageIntLLRInputS1xD(17)(5) <= VNStageIntLLROutputS0xD(357)(0);
  CNStageIntLLRInputS1xD(61)(5) <= VNStageIntLLROutputS0xD(357)(1);
  CNStageIntLLRInputS1xD(138)(5) <= VNStageIntLLROutputS0xD(357)(2);
  CNStageIntLLRInputS1xD(176)(5) <= VNStageIntLLROutputS0xD(357)(3);
  CNStageIntLLRInputS1xD(256)(5) <= VNStageIntLLROutputS0xD(357)(4);
  CNStageIntLLRInputS1xD(312)(5) <= VNStageIntLLROutputS0xD(357)(5);
  CNStageIntLLRInputS1xD(366)(5) <= VNStageIntLLROutputS0xD(357)(6);
  CNStageIntLLRInputS1xD(16)(5) <= VNStageIntLLROutputS0xD(358)(0);
  CNStageIntLLRInputS1xD(76)(5) <= VNStageIntLLROutputS0xD(358)(1);
  CNStageIntLLRInputS1xD(112)(5) <= VNStageIntLLROutputS0xD(358)(2);
  CNStageIntLLRInputS1xD(252)(5) <= VNStageIntLLROutputS0xD(358)(3);
  CNStageIntLLRInputS1xD(305)(5) <= VNStageIntLLROutputS0xD(358)(4);
  CNStageIntLLRInputS1xD(353)(5) <= VNStageIntLLROutputS0xD(358)(5);
  CNStageIntLLRInputS1xD(15)(5) <= VNStageIntLLROutputS0xD(359)(0);
  CNStageIntLLRInputS1xD(72)(5) <= VNStageIntLLROutputS0xD(359)(1);
  CNStageIntLLRInputS1xD(122)(5) <= VNStageIntLLROutputS0xD(359)(2);
  CNStageIntLLRInputS1xD(195)(5) <= VNStageIntLLROutputS0xD(359)(3);
  CNStageIntLLRInputS1xD(257)(5) <= VNStageIntLLROutputS0xD(359)(4);
  CNStageIntLLRInputS1xD(283)(5) <= VNStageIntLLROutputS0xD(359)(5);
  CNStageIntLLRInputS1xD(372)(5) <= VNStageIntLLROutputS0xD(359)(6);
  CNStageIntLLRInputS1xD(14)(5) <= VNStageIntLLROutputS0xD(360)(0);
  CNStageIntLLRInputS1xD(91)(5) <= VNStageIntLLROutputS0xD(360)(1);
  CNStageIntLLRInputS1xD(116)(5) <= VNStageIntLLROutputS0xD(360)(2);
  CNStageIntLLRInputS1xD(174)(5) <= VNStageIntLLROutputS0xD(360)(3);
  CNStageIntLLRInputS1xD(248)(5) <= VNStageIntLLROutputS0xD(360)(4);
  CNStageIntLLRInputS1xD(292)(5) <= VNStageIntLLROutputS0xD(360)(5);
  CNStageIntLLRInputS1xD(345)(5) <= VNStageIntLLROutputS0xD(360)(6);
  CNStageIntLLRInputS1xD(13)(5) <= VNStageIntLLROutputS0xD(361)(0);
  CNStageIntLLRInputS1xD(54)(5) <= VNStageIntLLROutputS0xD(361)(1);
  CNStageIntLLRInputS1xD(120)(5) <= VNStageIntLLROutputS0xD(361)(2);
  CNStageIntLLRInputS1xD(207)(5) <= VNStageIntLLROutputS0xD(361)(3);
  CNStageIntLLRInputS1xD(271)(5) <= VNStageIntLLROutputS0xD(361)(4);
  CNStageIntLLRInputS1xD(285)(5) <= VNStageIntLLROutputS0xD(361)(5);
  CNStageIntLLRInputS1xD(342)(5) <= VNStageIntLLROutputS0xD(361)(6);
  CNStageIntLLRInputS1xD(12)(5) <= VNStageIntLLROutputS0xD(362)(0);
  CNStageIntLLRInputS1xD(55)(5) <= VNStageIntLLROutputS0xD(362)(1);
  CNStageIntLLRInputS1xD(169)(5) <= VNStageIntLLROutputS0xD(362)(2);
  CNStageIntLLRInputS1xD(210)(5) <= VNStageIntLLROutputS0xD(362)(3);
  CNStageIntLLRInputS1xD(276)(5) <= VNStageIntLLROutputS0xD(362)(4);
  CNStageIntLLRInputS1xD(289)(5) <= VNStageIntLLROutputS0xD(362)(5);
  CNStageIntLLRInputS1xD(357)(5) <= VNStageIntLLROutputS0xD(362)(6);
  CNStageIntLLRInputS1xD(90)(5) <= VNStageIntLLROutputS0xD(363)(0);
  CNStageIntLLRInputS1xD(147)(5) <= VNStageIntLLROutputS0xD(363)(1);
  CNStageIntLLRInputS1xD(197)(5) <= VNStageIntLLROutputS0xD(363)(2);
  CNStageIntLLRInputS1xD(261)(5) <= VNStageIntLLROutputS0xD(363)(3);
  CNStageIntLLRInputS1xD(281)(5) <= VNStageIntLLROutputS0xD(363)(4);
  CNStageIntLLRInputS1xD(11)(5) <= VNStageIntLLROutputS0xD(364)(0);
  CNStageIntLLRInputS1xD(82)(5) <= VNStageIntLLROutputS0xD(364)(1);
  CNStageIntLLRInputS1xD(129)(5) <= VNStageIntLLROutputS0xD(364)(2);
  CNStageIntLLRInputS1xD(175)(5) <= VNStageIntLLROutputS0xD(364)(3);
  CNStageIntLLRInputS1xD(263)(5) <= VNStageIntLLROutputS0xD(364)(4);
  CNStageIntLLRInputS1xD(313)(5) <= VNStageIntLLROutputS0xD(364)(5);
  CNStageIntLLRInputS1xD(10)(5) <= VNStageIntLLROutputS0xD(365)(0);
  CNStageIntLLRInputS1xD(98)(5) <= VNStageIntLLROutputS0xD(365)(1);
  CNStageIntLLRInputS1xD(142)(5) <= VNStageIntLLROutputS0xD(365)(2);
  CNStageIntLLRInputS1xD(194)(5) <= VNStageIntLLROutputS0xD(365)(3);
  CNStageIntLLRInputS1xD(234)(5) <= VNStageIntLLROutputS0xD(365)(4);
  CNStageIntLLRInputS1xD(298)(5) <= VNStageIntLLROutputS0xD(365)(5);
  CNStageIntLLRInputS1xD(9)(5) <= VNStageIntLLROutputS0xD(366)(0);
  CNStageIntLLRInputS1xD(102)(5) <= VNStageIntLLROutputS0xD(366)(1);
  CNStageIntLLRInputS1xD(153)(5) <= VNStageIntLLROutputS0xD(366)(2);
  CNStageIntLLRInputS1xD(219)(5) <= VNStageIntLLROutputS0xD(366)(3);
  CNStageIntLLRInputS1xD(269)(5) <= VNStageIntLLROutputS0xD(366)(4);
  CNStageIntLLRInputS1xD(308)(5) <= VNStageIntLLROutputS0xD(366)(5);
  CNStageIntLLRInputS1xD(8)(5) <= VNStageIntLLROutputS0xD(367)(0);
  CNStageIntLLRInputS1xD(110)(5) <= VNStageIntLLROutputS0xD(367)(1);
  CNStageIntLLRInputS1xD(123)(5) <= VNStageIntLLROutputS0xD(367)(2);
  CNStageIntLLRInputS1xD(205)(5) <= VNStageIntLLROutputS0xD(367)(3);
  CNStageIntLLRInputS1xD(226)(5) <= VNStageIntLLROutputS0xD(367)(4);
  CNStageIntLLRInputS1xD(320)(5) <= VNStageIntLLROutputS0xD(367)(5);
  CNStageIntLLRInputS1xD(333)(5) <= VNStageIntLLROutputS0xD(367)(6);
  CNStageIntLLRInputS1xD(7)(5) <= VNStageIntLLROutputS0xD(368)(0);
  CNStageIntLLRInputS1xD(177)(5) <= VNStageIntLLROutputS0xD(368)(1);
  CNStageIntLLRInputS1xD(381)(5) <= VNStageIntLLROutputS0xD(368)(2);
  CNStageIntLLRInputS1xD(6)(5) <= VNStageIntLLROutputS0xD(369)(0);
  CNStageIntLLRInputS1xD(156)(5) <= VNStageIntLLROutputS0xD(369)(1);
  CNStageIntLLRInputS1xD(221)(5) <= VNStageIntLLROutputS0xD(369)(2);
  CNStageIntLLRInputS1xD(262)(5) <= VNStageIntLLROutputS0xD(369)(3);
  CNStageIntLLRInputS1xD(358)(5) <= VNStageIntLLROutputS0xD(369)(4);
  CNStageIntLLRInputS1xD(5)(5) <= VNStageIntLLROutputS0xD(370)(0);
  CNStageIntLLRInputS1xD(114)(5) <= VNStageIntLLROutputS0xD(370)(1);
  CNStageIntLLRInputS1xD(208)(5) <= VNStageIntLLROutputS0xD(370)(2);
  CNStageIntLLRInputS1xD(275)(5) <= VNStageIntLLROutputS0xD(370)(3);
  CNStageIntLLRInputS1xD(341)(5) <= VNStageIntLLROutputS0xD(370)(4);
  CNStageIntLLRInputS1xD(4)(5) <= VNStageIntLLROutputS0xD(371)(0);
  CNStageIntLLRInputS1xD(135)(5) <= VNStageIntLLROutputS0xD(371)(1);
  CNStageIntLLRInputS1xD(173)(5) <= VNStageIntLLROutputS0xD(371)(2);
  CNStageIntLLRInputS1xD(249)(5) <= VNStageIntLLROutputS0xD(371)(3);
  CNStageIntLLRInputS1xD(354)(5) <= VNStageIntLLROutputS0xD(371)(4);
  CNStageIntLLRInputS1xD(106)(5) <= VNStageIntLLROutputS0xD(372)(0);
  CNStageIntLLRInputS1xD(144)(5) <= VNStageIntLLROutputS0xD(372)(1);
  CNStageIntLLRInputS1xD(201)(5) <= VNStageIntLLROutputS0xD(372)(2);
  CNStageIntLLRInputS1xD(229)(5) <= VNStageIntLLROutputS0xD(372)(3);
  CNStageIntLLRInputS1xD(301)(5) <= VNStageIntLLROutputS0xD(372)(4);
  CNStageIntLLRInputS1xD(365)(5) <= VNStageIntLLROutputS0xD(372)(5);
  CNStageIntLLRInputS1xD(3)(5) <= VNStageIntLLROutputS0xD(373)(0);
  CNStageIntLLRInputS1xD(139)(5) <= VNStageIntLLROutputS0xD(373)(1);
  CNStageIntLLRInputS1xD(250)(5) <= VNStageIntLLROutputS0xD(373)(2);
  CNStageIntLLRInputS1xD(310)(5) <= VNStageIntLLROutputS0xD(373)(3);
  CNStageIntLLRInputS1xD(335)(5) <= VNStageIntLLROutputS0xD(373)(4);
  CNStageIntLLRInputS1xD(2)(5) <= VNStageIntLLROutputS0xD(374)(0);
  CNStageIntLLRInputS1xD(85)(5) <= VNStageIntLLROutputS0xD(374)(1);
  CNStageIntLLRInputS1xD(145)(5) <= VNStageIntLLROutputS0xD(374)(2);
  CNStageIntLLRInputS1xD(213)(5) <= VNStageIntLLROutputS0xD(374)(3);
  CNStageIntLLRInputS1xD(264)(5) <= VNStageIntLLROutputS0xD(374)(4);
  CNStageIntLLRInputS1xD(306)(5) <= VNStageIntLLROutputS0xD(374)(5);
  CNStageIntLLRInputS1xD(383)(5) <= VNStageIntLLROutputS0xD(374)(6);
  CNStageIntLLRInputS1xD(1)(5) <= VNStageIntLLROutputS0xD(375)(0);
  CNStageIntLLRInputS1xD(64)(5) <= VNStageIntLLROutputS0xD(375)(1);
  CNStageIntLLRInputS1xD(134)(5) <= VNStageIntLLROutputS0xD(375)(2);
  CNStageIntLLRInputS1xD(260)(5) <= VNStageIntLLROutputS0xD(375)(3);
  CNStageIntLLRInputS1xD(311)(5) <= VNStageIntLLROutputS0xD(375)(4);
  CNStageIntLLRInputS1xD(368)(5) <= VNStageIntLLROutputS0xD(375)(5);
  CNStageIntLLRInputS1xD(0)(5) <= VNStageIntLLROutputS0xD(376)(0);
  CNStageIntLLRInputS1xD(67)(5) <= VNStageIntLLROutputS0xD(376)(1);
  CNStageIntLLRInputS1xD(159)(5) <= VNStageIntLLROutputS0xD(376)(2);
  CNStageIntLLRInputS1xD(278)(5) <= VNStageIntLLROutputS0xD(376)(3);
  CNStageIntLLRInputS1xD(107)(5) <= VNStageIntLLROutputS0xD(377)(0);
  CNStageIntLLRInputS1xD(166)(5) <= VNStageIntLLROutputS0xD(377)(1);
  CNStageIntLLRInputS1xD(193)(5) <= VNStageIntLLROutputS0xD(377)(2);
  CNStageIntLLRInputS1xD(325)(5) <= VNStageIntLLROutputS0xD(377)(3);
  CNStageIntLLRInputS1xD(347)(5) <= VNStageIntLLROutputS0xD(377)(4);
  CNStageIntLLRInputS1xD(86)(5) <= VNStageIntLLROutputS0xD(378)(0);
  CNStageIntLLRInputS1xD(149)(5) <= VNStageIntLLROutputS0xD(378)(1);
  CNStageIntLLRInputS1xD(187)(5) <= VNStageIntLLROutputS0xD(378)(2);
  CNStageIntLLRInputS1xD(246)(5) <= VNStageIntLLROutputS0xD(378)(3);
  CNStageIntLLRInputS1xD(331)(5) <= VNStageIntLLROutputS0xD(378)(4);
  CNStageIntLLRInputS1xD(355)(5) <= VNStageIntLLROutputS0xD(378)(5);
  CNStageIntLLRInputS1xD(105)(5) <= VNStageIntLLROutputS0xD(379)(0);
  CNStageIntLLRInputS1xD(151)(5) <= VNStageIntLLROutputS0xD(379)(1);
  CNStageIntLLRInputS1xD(277)(5) <= VNStageIntLLROutputS0xD(379)(2);
  CNStageIntLLRInputS1xD(315)(5) <= VNStageIntLLROutputS0xD(379)(3);
  CNStageIntLLRInputS1xD(351)(5) <= VNStageIntLLROutputS0xD(379)(4);
  CNStageIntLLRInputS1xD(77)(5) <= VNStageIntLLROutputS0xD(380)(0);
  CNStageIntLLRInputS1xD(118)(5) <= VNStageIntLLROutputS0xD(380)(1);
  CNStageIntLLRInputS1xD(182)(5) <= VNStageIntLLROutputS0xD(380)(2);
  CNStageIntLLRInputS1xD(270)(5) <= VNStageIntLLROutputS0xD(380)(3);
  CNStageIntLLRInputS1xD(317)(5) <= VNStageIntLLROutputS0xD(380)(4);
  CNStageIntLLRInputS1xD(356)(5) <= VNStageIntLLROutputS0xD(380)(5);
  CNStageIntLLRInputS1xD(60)(5) <= VNStageIntLLROutputS0xD(381)(0);
  CNStageIntLLRInputS1xD(157)(5) <= VNStageIntLLROutputS0xD(381)(1);
  CNStageIntLLRInputS1xD(214)(5) <= VNStageIntLLROutputS0xD(381)(2);
  CNStageIntLLRInputS1xD(233)(5) <= VNStageIntLLROutputS0xD(381)(3);
  CNStageIntLLRInputS1xD(287)(5) <= VNStageIntLLROutputS0xD(381)(4);
  CNStageIntLLRInputS1xD(346)(5) <= VNStageIntLLROutputS0xD(381)(5);
  CNStageIntLLRInputS1xD(87)(5) <= VNStageIntLLROutputS0xD(382)(0);
  CNStageIntLLRInputS1xD(111)(5) <= VNStageIntLLROutputS0xD(382)(1);
  CNStageIntLLRInputS1xD(198)(5) <= VNStageIntLLROutputS0xD(382)(2);
  CNStageIntLLRInputS1xD(237)(5) <= VNStageIntLLROutputS0xD(382)(3);
  CNStageIntLLRInputS1xD(323)(5) <= VNStageIntLLROutputS0xD(382)(4);
  CNStageIntLLRInputS1xD(371)(5) <= VNStageIntLLROutputS0xD(382)(5);
  CNStageIntLLRInputS1xD(52)(5) <= VNStageIntLLROutputS0xD(383)(0);
  CNStageIntLLRInputS1xD(79)(5) <= VNStageIntLLROutputS0xD(383)(1);
  CNStageIntLLRInputS1xD(119)(5) <= VNStageIntLLROutputS0xD(383)(2);
  CNStageIntLLRInputS1xD(209)(5) <= VNStageIntLLROutputS0xD(383)(3);
  CNStageIntLLRInputS1xD(279)(5) <= VNStageIntLLROutputS0xD(383)(4);
  CNStageIntLLRInputS1xD(282)(5) <= VNStageIntLLROutputS0xD(383)(5);
  CNStageIntLLRInputS1xD(378)(5) <= VNStageIntLLROutputS0xD(383)(6);

  -- Variable Nodes (Iteration 1)
  VNStageIntLLRInputS1xD(56)(0) <= CNStageIntLLROutputS1xD(0)(0);
  VNStageIntLLRInputS1xD(120)(0) <= CNStageIntLLROutputS1xD(0)(1);
  VNStageIntLLRInputS1xD(184)(0) <= CNStageIntLLROutputS1xD(0)(2);
  VNStageIntLLRInputS1xD(248)(0) <= CNStageIntLLROutputS1xD(0)(3);
  VNStageIntLLRInputS1xD(312)(0) <= CNStageIntLLROutputS1xD(0)(4);
  VNStageIntLLRInputS1xD(376)(0) <= CNStageIntLLROutputS1xD(0)(5);
  VNStageIntLLRInputS1xD(55)(0) <= CNStageIntLLROutputS1xD(1)(0);
  VNStageIntLLRInputS1xD(119)(0) <= CNStageIntLLROutputS1xD(1)(1);
  VNStageIntLLRInputS1xD(183)(0) <= CNStageIntLLROutputS1xD(1)(2);
  VNStageIntLLRInputS1xD(247)(0) <= CNStageIntLLROutputS1xD(1)(3);
  VNStageIntLLRInputS1xD(311)(0) <= CNStageIntLLROutputS1xD(1)(4);
  VNStageIntLLRInputS1xD(375)(0) <= CNStageIntLLROutputS1xD(1)(5);
  VNStageIntLLRInputS1xD(54)(0) <= CNStageIntLLROutputS1xD(2)(0);
  VNStageIntLLRInputS1xD(118)(0) <= CNStageIntLLROutputS1xD(2)(1);
  VNStageIntLLRInputS1xD(182)(0) <= CNStageIntLLROutputS1xD(2)(2);
  VNStageIntLLRInputS1xD(246)(0) <= CNStageIntLLROutputS1xD(2)(3);
  VNStageIntLLRInputS1xD(310)(0) <= CNStageIntLLROutputS1xD(2)(4);
  VNStageIntLLRInputS1xD(374)(0) <= CNStageIntLLROutputS1xD(2)(5);
  VNStageIntLLRInputS1xD(53)(0) <= CNStageIntLLROutputS1xD(3)(0);
  VNStageIntLLRInputS1xD(117)(0) <= CNStageIntLLROutputS1xD(3)(1);
  VNStageIntLLRInputS1xD(181)(0) <= CNStageIntLLROutputS1xD(3)(2);
  VNStageIntLLRInputS1xD(245)(0) <= CNStageIntLLROutputS1xD(3)(3);
  VNStageIntLLRInputS1xD(309)(0) <= CNStageIntLLROutputS1xD(3)(4);
  VNStageIntLLRInputS1xD(373)(0) <= CNStageIntLLROutputS1xD(3)(5);
  VNStageIntLLRInputS1xD(51)(0) <= CNStageIntLLROutputS1xD(4)(0);
  VNStageIntLLRInputS1xD(115)(0) <= CNStageIntLLROutputS1xD(4)(1);
  VNStageIntLLRInputS1xD(179)(0) <= CNStageIntLLROutputS1xD(4)(2);
  VNStageIntLLRInputS1xD(243)(0) <= CNStageIntLLROutputS1xD(4)(3);
  VNStageIntLLRInputS1xD(307)(0) <= CNStageIntLLROutputS1xD(4)(4);
  VNStageIntLLRInputS1xD(371)(0) <= CNStageIntLLROutputS1xD(4)(5);
  VNStageIntLLRInputS1xD(50)(0) <= CNStageIntLLROutputS1xD(5)(0);
  VNStageIntLLRInputS1xD(114)(0) <= CNStageIntLLROutputS1xD(5)(1);
  VNStageIntLLRInputS1xD(178)(0) <= CNStageIntLLROutputS1xD(5)(2);
  VNStageIntLLRInputS1xD(242)(0) <= CNStageIntLLROutputS1xD(5)(3);
  VNStageIntLLRInputS1xD(306)(0) <= CNStageIntLLROutputS1xD(5)(4);
  VNStageIntLLRInputS1xD(370)(0) <= CNStageIntLLROutputS1xD(5)(5);
  VNStageIntLLRInputS1xD(49)(0) <= CNStageIntLLROutputS1xD(6)(0);
  VNStageIntLLRInputS1xD(113)(0) <= CNStageIntLLROutputS1xD(6)(1);
  VNStageIntLLRInputS1xD(177)(0) <= CNStageIntLLROutputS1xD(6)(2);
  VNStageIntLLRInputS1xD(241)(0) <= CNStageIntLLROutputS1xD(6)(3);
  VNStageIntLLRInputS1xD(305)(0) <= CNStageIntLLROutputS1xD(6)(4);
  VNStageIntLLRInputS1xD(369)(0) <= CNStageIntLLROutputS1xD(6)(5);
  VNStageIntLLRInputS1xD(48)(0) <= CNStageIntLLROutputS1xD(7)(0);
  VNStageIntLLRInputS1xD(112)(0) <= CNStageIntLLROutputS1xD(7)(1);
  VNStageIntLLRInputS1xD(176)(0) <= CNStageIntLLROutputS1xD(7)(2);
  VNStageIntLLRInputS1xD(240)(0) <= CNStageIntLLROutputS1xD(7)(3);
  VNStageIntLLRInputS1xD(304)(0) <= CNStageIntLLROutputS1xD(7)(4);
  VNStageIntLLRInputS1xD(368)(0) <= CNStageIntLLROutputS1xD(7)(5);
  VNStageIntLLRInputS1xD(47)(0) <= CNStageIntLLROutputS1xD(8)(0);
  VNStageIntLLRInputS1xD(111)(0) <= CNStageIntLLROutputS1xD(8)(1);
  VNStageIntLLRInputS1xD(175)(0) <= CNStageIntLLROutputS1xD(8)(2);
  VNStageIntLLRInputS1xD(239)(0) <= CNStageIntLLROutputS1xD(8)(3);
  VNStageIntLLRInputS1xD(303)(0) <= CNStageIntLLROutputS1xD(8)(4);
  VNStageIntLLRInputS1xD(367)(0) <= CNStageIntLLROutputS1xD(8)(5);
  VNStageIntLLRInputS1xD(46)(0) <= CNStageIntLLROutputS1xD(9)(0);
  VNStageIntLLRInputS1xD(110)(0) <= CNStageIntLLROutputS1xD(9)(1);
  VNStageIntLLRInputS1xD(174)(0) <= CNStageIntLLROutputS1xD(9)(2);
  VNStageIntLLRInputS1xD(238)(0) <= CNStageIntLLROutputS1xD(9)(3);
  VNStageIntLLRInputS1xD(302)(0) <= CNStageIntLLROutputS1xD(9)(4);
  VNStageIntLLRInputS1xD(366)(0) <= CNStageIntLLROutputS1xD(9)(5);
  VNStageIntLLRInputS1xD(45)(0) <= CNStageIntLLROutputS1xD(10)(0);
  VNStageIntLLRInputS1xD(109)(0) <= CNStageIntLLROutputS1xD(10)(1);
  VNStageIntLLRInputS1xD(173)(0) <= CNStageIntLLROutputS1xD(10)(2);
  VNStageIntLLRInputS1xD(237)(0) <= CNStageIntLLROutputS1xD(10)(3);
  VNStageIntLLRInputS1xD(301)(0) <= CNStageIntLLROutputS1xD(10)(4);
  VNStageIntLLRInputS1xD(365)(0) <= CNStageIntLLROutputS1xD(10)(5);
  VNStageIntLLRInputS1xD(44)(0) <= CNStageIntLLROutputS1xD(11)(0);
  VNStageIntLLRInputS1xD(108)(0) <= CNStageIntLLROutputS1xD(11)(1);
  VNStageIntLLRInputS1xD(172)(0) <= CNStageIntLLROutputS1xD(11)(2);
  VNStageIntLLRInputS1xD(236)(0) <= CNStageIntLLROutputS1xD(11)(3);
  VNStageIntLLRInputS1xD(300)(0) <= CNStageIntLLROutputS1xD(11)(4);
  VNStageIntLLRInputS1xD(364)(0) <= CNStageIntLLROutputS1xD(11)(5);
  VNStageIntLLRInputS1xD(42)(0) <= CNStageIntLLROutputS1xD(12)(0);
  VNStageIntLLRInputS1xD(106)(0) <= CNStageIntLLROutputS1xD(12)(1);
  VNStageIntLLRInputS1xD(170)(0) <= CNStageIntLLROutputS1xD(12)(2);
  VNStageIntLLRInputS1xD(234)(0) <= CNStageIntLLROutputS1xD(12)(3);
  VNStageIntLLRInputS1xD(298)(0) <= CNStageIntLLROutputS1xD(12)(4);
  VNStageIntLLRInputS1xD(362)(0) <= CNStageIntLLROutputS1xD(12)(5);
  VNStageIntLLRInputS1xD(41)(0) <= CNStageIntLLROutputS1xD(13)(0);
  VNStageIntLLRInputS1xD(105)(0) <= CNStageIntLLROutputS1xD(13)(1);
  VNStageIntLLRInputS1xD(169)(0) <= CNStageIntLLROutputS1xD(13)(2);
  VNStageIntLLRInputS1xD(233)(0) <= CNStageIntLLROutputS1xD(13)(3);
  VNStageIntLLRInputS1xD(297)(0) <= CNStageIntLLROutputS1xD(13)(4);
  VNStageIntLLRInputS1xD(361)(0) <= CNStageIntLLROutputS1xD(13)(5);
  VNStageIntLLRInputS1xD(40)(0) <= CNStageIntLLROutputS1xD(14)(0);
  VNStageIntLLRInputS1xD(104)(0) <= CNStageIntLLROutputS1xD(14)(1);
  VNStageIntLLRInputS1xD(168)(0) <= CNStageIntLLROutputS1xD(14)(2);
  VNStageIntLLRInputS1xD(232)(0) <= CNStageIntLLROutputS1xD(14)(3);
  VNStageIntLLRInputS1xD(296)(0) <= CNStageIntLLROutputS1xD(14)(4);
  VNStageIntLLRInputS1xD(360)(0) <= CNStageIntLLROutputS1xD(14)(5);
  VNStageIntLLRInputS1xD(39)(0) <= CNStageIntLLROutputS1xD(15)(0);
  VNStageIntLLRInputS1xD(103)(0) <= CNStageIntLLROutputS1xD(15)(1);
  VNStageIntLLRInputS1xD(167)(0) <= CNStageIntLLROutputS1xD(15)(2);
  VNStageIntLLRInputS1xD(231)(0) <= CNStageIntLLROutputS1xD(15)(3);
  VNStageIntLLRInputS1xD(295)(0) <= CNStageIntLLROutputS1xD(15)(4);
  VNStageIntLLRInputS1xD(359)(0) <= CNStageIntLLROutputS1xD(15)(5);
  VNStageIntLLRInputS1xD(38)(0) <= CNStageIntLLROutputS1xD(16)(0);
  VNStageIntLLRInputS1xD(102)(0) <= CNStageIntLLROutputS1xD(16)(1);
  VNStageIntLLRInputS1xD(166)(0) <= CNStageIntLLROutputS1xD(16)(2);
  VNStageIntLLRInputS1xD(230)(0) <= CNStageIntLLROutputS1xD(16)(3);
  VNStageIntLLRInputS1xD(294)(0) <= CNStageIntLLROutputS1xD(16)(4);
  VNStageIntLLRInputS1xD(358)(0) <= CNStageIntLLROutputS1xD(16)(5);
  VNStageIntLLRInputS1xD(37)(0) <= CNStageIntLLROutputS1xD(17)(0);
  VNStageIntLLRInputS1xD(101)(0) <= CNStageIntLLROutputS1xD(17)(1);
  VNStageIntLLRInputS1xD(165)(0) <= CNStageIntLLROutputS1xD(17)(2);
  VNStageIntLLRInputS1xD(229)(0) <= CNStageIntLLROutputS1xD(17)(3);
  VNStageIntLLRInputS1xD(293)(0) <= CNStageIntLLROutputS1xD(17)(4);
  VNStageIntLLRInputS1xD(357)(0) <= CNStageIntLLROutputS1xD(17)(5);
  VNStageIntLLRInputS1xD(36)(0) <= CNStageIntLLROutputS1xD(18)(0);
  VNStageIntLLRInputS1xD(100)(0) <= CNStageIntLLROutputS1xD(18)(1);
  VNStageIntLLRInputS1xD(164)(0) <= CNStageIntLLROutputS1xD(18)(2);
  VNStageIntLLRInputS1xD(228)(0) <= CNStageIntLLROutputS1xD(18)(3);
  VNStageIntLLRInputS1xD(292)(0) <= CNStageIntLLROutputS1xD(18)(4);
  VNStageIntLLRInputS1xD(356)(0) <= CNStageIntLLROutputS1xD(18)(5);
  VNStageIntLLRInputS1xD(35)(0) <= CNStageIntLLROutputS1xD(19)(0);
  VNStageIntLLRInputS1xD(99)(0) <= CNStageIntLLROutputS1xD(19)(1);
  VNStageIntLLRInputS1xD(163)(0) <= CNStageIntLLROutputS1xD(19)(2);
  VNStageIntLLRInputS1xD(227)(0) <= CNStageIntLLROutputS1xD(19)(3);
  VNStageIntLLRInputS1xD(291)(0) <= CNStageIntLLROutputS1xD(19)(4);
  VNStageIntLLRInputS1xD(355)(0) <= CNStageIntLLROutputS1xD(19)(5);
  VNStageIntLLRInputS1xD(34)(0) <= CNStageIntLLROutputS1xD(20)(0);
  VNStageIntLLRInputS1xD(98)(0) <= CNStageIntLLROutputS1xD(20)(1);
  VNStageIntLLRInputS1xD(162)(0) <= CNStageIntLLROutputS1xD(20)(2);
  VNStageIntLLRInputS1xD(226)(0) <= CNStageIntLLROutputS1xD(20)(3);
  VNStageIntLLRInputS1xD(290)(0) <= CNStageIntLLROutputS1xD(20)(4);
  VNStageIntLLRInputS1xD(354)(0) <= CNStageIntLLROutputS1xD(20)(5);
  VNStageIntLLRInputS1xD(33)(0) <= CNStageIntLLROutputS1xD(21)(0);
  VNStageIntLLRInputS1xD(97)(0) <= CNStageIntLLROutputS1xD(21)(1);
  VNStageIntLLRInputS1xD(161)(0) <= CNStageIntLLROutputS1xD(21)(2);
  VNStageIntLLRInputS1xD(225)(0) <= CNStageIntLLROutputS1xD(21)(3);
  VNStageIntLLRInputS1xD(289)(0) <= CNStageIntLLROutputS1xD(21)(4);
  VNStageIntLLRInputS1xD(353)(0) <= CNStageIntLLROutputS1xD(21)(5);
  VNStageIntLLRInputS1xD(32)(0) <= CNStageIntLLROutputS1xD(22)(0);
  VNStageIntLLRInputS1xD(96)(0) <= CNStageIntLLROutputS1xD(22)(1);
  VNStageIntLLRInputS1xD(160)(0) <= CNStageIntLLROutputS1xD(22)(2);
  VNStageIntLLRInputS1xD(224)(0) <= CNStageIntLLROutputS1xD(22)(3);
  VNStageIntLLRInputS1xD(288)(0) <= CNStageIntLLROutputS1xD(22)(4);
  VNStageIntLLRInputS1xD(352)(0) <= CNStageIntLLROutputS1xD(22)(5);
  VNStageIntLLRInputS1xD(31)(0) <= CNStageIntLLROutputS1xD(23)(0);
  VNStageIntLLRInputS1xD(95)(0) <= CNStageIntLLROutputS1xD(23)(1);
  VNStageIntLLRInputS1xD(159)(0) <= CNStageIntLLROutputS1xD(23)(2);
  VNStageIntLLRInputS1xD(223)(0) <= CNStageIntLLROutputS1xD(23)(3);
  VNStageIntLLRInputS1xD(287)(0) <= CNStageIntLLROutputS1xD(23)(4);
  VNStageIntLLRInputS1xD(351)(0) <= CNStageIntLLROutputS1xD(23)(5);
  VNStageIntLLRInputS1xD(30)(0) <= CNStageIntLLROutputS1xD(24)(0);
  VNStageIntLLRInputS1xD(94)(0) <= CNStageIntLLROutputS1xD(24)(1);
  VNStageIntLLRInputS1xD(158)(0) <= CNStageIntLLROutputS1xD(24)(2);
  VNStageIntLLRInputS1xD(222)(0) <= CNStageIntLLROutputS1xD(24)(3);
  VNStageIntLLRInputS1xD(286)(0) <= CNStageIntLLROutputS1xD(24)(4);
  VNStageIntLLRInputS1xD(350)(0) <= CNStageIntLLROutputS1xD(24)(5);
  VNStageIntLLRInputS1xD(29)(0) <= CNStageIntLLROutputS1xD(25)(0);
  VNStageIntLLRInputS1xD(93)(0) <= CNStageIntLLROutputS1xD(25)(1);
  VNStageIntLLRInputS1xD(157)(0) <= CNStageIntLLROutputS1xD(25)(2);
  VNStageIntLLRInputS1xD(221)(0) <= CNStageIntLLROutputS1xD(25)(3);
  VNStageIntLLRInputS1xD(285)(0) <= CNStageIntLLROutputS1xD(25)(4);
  VNStageIntLLRInputS1xD(349)(0) <= CNStageIntLLROutputS1xD(25)(5);
  VNStageIntLLRInputS1xD(28)(0) <= CNStageIntLLROutputS1xD(26)(0);
  VNStageIntLLRInputS1xD(92)(0) <= CNStageIntLLROutputS1xD(26)(1);
  VNStageIntLLRInputS1xD(156)(0) <= CNStageIntLLROutputS1xD(26)(2);
  VNStageIntLLRInputS1xD(220)(0) <= CNStageIntLLROutputS1xD(26)(3);
  VNStageIntLLRInputS1xD(284)(0) <= CNStageIntLLROutputS1xD(26)(4);
  VNStageIntLLRInputS1xD(348)(0) <= CNStageIntLLROutputS1xD(26)(5);
  VNStageIntLLRInputS1xD(27)(0) <= CNStageIntLLROutputS1xD(27)(0);
  VNStageIntLLRInputS1xD(91)(0) <= CNStageIntLLROutputS1xD(27)(1);
  VNStageIntLLRInputS1xD(155)(0) <= CNStageIntLLROutputS1xD(27)(2);
  VNStageIntLLRInputS1xD(219)(0) <= CNStageIntLLROutputS1xD(27)(3);
  VNStageIntLLRInputS1xD(283)(0) <= CNStageIntLLROutputS1xD(27)(4);
  VNStageIntLLRInputS1xD(347)(0) <= CNStageIntLLROutputS1xD(27)(5);
  VNStageIntLLRInputS1xD(26)(0) <= CNStageIntLLROutputS1xD(28)(0);
  VNStageIntLLRInputS1xD(90)(0) <= CNStageIntLLROutputS1xD(28)(1);
  VNStageIntLLRInputS1xD(154)(0) <= CNStageIntLLROutputS1xD(28)(2);
  VNStageIntLLRInputS1xD(218)(0) <= CNStageIntLLROutputS1xD(28)(3);
  VNStageIntLLRInputS1xD(282)(0) <= CNStageIntLLROutputS1xD(28)(4);
  VNStageIntLLRInputS1xD(346)(0) <= CNStageIntLLROutputS1xD(28)(5);
  VNStageIntLLRInputS1xD(25)(0) <= CNStageIntLLROutputS1xD(29)(0);
  VNStageIntLLRInputS1xD(89)(0) <= CNStageIntLLROutputS1xD(29)(1);
  VNStageIntLLRInputS1xD(153)(0) <= CNStageIntLLROutputS1xD(29)(2);
  VNStageIntLLRInputS1xD(217)(0) <= CNStageIntLLROutputS1xD(29)(3);
  VNStageIntLLRInputS1xD(281)(0) <= CNStageIntLLROutputS1xD(29)(4);
  VNStageIntLLRInputS1xD(345)(0) <= CNStageIntLLROutputS1xD(29)(5);
  VNStageIntLLRInputS1xD(24)(0) <= CNStageIntLLROutputS1xD(30)(0);
  VNStageIntLLRInputS1xD(88)(0) <= CNStageIntLLROutputS1xD(30)(1);
  VNStageIntLLRInputS1xD(152)(0) <= CNStageIntLLROutputS1xD(30)(2);
  VNStageIntLLRInputS1xD(216)(0) <= CNStageIntLLROutputS1xD(30)(3);
  VNStageIntLLRInputS1xD(280)(0) <= CNStageIntLLROutputS1xD(30)(4);
  VNStageIntLLRInputS1xD(344)(0) <= CNStageIntLLROutputS1xD(30)(5);
  VNStageIntLLRInputS1xD(23)(0) <= CNStageIntLLROutputS1xD(31)(0);
  VNStageIntLLRInputS1xD(87)(0) <= CNStageIntLLROutputS1xD(31)(1);
  VNStageIntLLRInputS1xD(151)(0) <= CNStageIntLLROutputS1xD(31)(2);
  VNStageIntLLRInputS1xD(215)(0) <= CNStageIntLLROutputS1xD(31)(3);
  VNStageIntLLRInputS1xD(279)(0) <= CNStageIntLLROutputS1xD(31)(4);
  VNStageIntLLRInputS1xD(343)(0) <= CNStageIntLLROutputS1xD(31)(5);
  VNStageIntLLRInputS1xD(22)(0) <= CNStageIntLLROutputS1xD(32)(0);
  VNStageIntLLRInputS1xD(86)(0) <= CNStageIntLLROutputS1xD(32)(1);
  VNStageIntLLRInputS1xD(150)(0) <= CNStageIntLLROutputS1xD(32)(2);
  VNStageIntLLRInputS1xD(214)(0) <= CNStageIntLLROutputS1xD(32)(3);
  VNStageIntLLRInputS1xD(278)(0) <= CNStageIntLLROutputS1xD(32)(4);
  VNStageIntLLRInputS1xD(342)(0) <= CNStageIntLLROutputS1xD(32)(5);
  VNStageIntLLRInputS1xD(21)(0) <= CNStageIntLLROutputS1xD(33)(0);
  VNStageIntLLRInputS1xD(85)(0) <= CNStageIntLLROutputS1xD(33)(1);
  VNStageIntLLRInputS1xD(149)(0) <= CNStageIntLLROutputS1xD(33)(2);
  VNStageIntLLRInputS1xD(213)(0) <= CNStageIntLLROutputS1xD(33)(3);
  VNStageIntLLRInputS1xD(277)(0) <= CNStageIntLLROutputS1xD(33)(4);
  VNStageIntLLRInputS1xD(341)(0) <= CNStageIntLLROutputS1xD(33)(5);
  VNStageIntLLRInputS1xD(20)(0) <= CNStageIntLLROutputS1xD(34)(0);
  VNStageIntLLRInputS1xD(84)(0) <= CNStageIntLLROutputS1xD(34)(1);
  VNStageIntLLRInputS1xD(148)(0) <= CNStageIntLLROutputS1xD(34)(2);
  VNStageIntLLRInputS1xD(212)(0) <= CNStageIntLLROutputS1xD(34)(3);
  VNStageIntLLRInputS1xD(276)(0) <= CNStageIntLLROutputS1xD(34)(4);
  VNStageIntLLRInputS1xD(340)(0) <= CNStageIntLLROutputS1xD(34)(5);
  VNStageIntLLRInputS1xD(19)(0) <= CNStageIntLLROutputS1xD(35)(0);
  VNStageIntLLRInputS1xD(83)(0) <= CNStageIntLLROutputS1xD(35)(1);
  VNStageIntLLRInputS1xD(147)(0) <= CNStageIntLLROutputS1xD(35)(2);
  VNStageIntLLRInputS1xD(211)(0) <= CNStageIntLLROutputS1xD(35)(3);
  VNStageIntLLRInputS1xD(275)(0) <= CNStageIntLLROutputS1xD(35)(4);
  VNStageIntLLRInputS1xD(339)(0) <= CNStageIntLLROutputS1xD(35)(5);
  VNStageIntLLRInputS1xD(18)(0) <= CNStageIntLLROutputS1xD(36)(0);
  VNStageIntLLRInputS1xD(82)(0) <= CNStageIntLLROutputS1xD(36)(1);
  VNStageIntLLRInputS1xD(146)(0) <= CNStageIntLLROutputS1xD(36)(2);
  VNStageIntLLRInputS1xD(210)(0) <= CNStageIntLLROutputS1xD(36)(3);
  VNStageIntLLRInputS1xD(274)(0) <= CNStageIntLLROutputS1xD(36)(4);
  VNStageIntLLRInputS1xD(338)(0) <= CNStageIntLLROutputS1xD(36)(5);
  VNStageIntLLRInputS1xD(17)(0) <= CNStageIntLLROutputS1xD(37)(0);
  VNStageIntLLRInputS1xD(81)(0) <= CNStageIntLLROutputS1xD(37)(1);
  VNStageIntLLRInputS1xD(145)(0) <= CNStageIntLLROutputS1xD(37)(2);
  VNStageIntLLRInputS1xD(209)(0) <= CNStageIntLLROutputS1xD(37)(3);
  VNStageIntLLRInputS1xD(273)(0) <= CNStageIntLLROutputS1xD(37)(4);
  VNStageIntLLRInputS1xD(337)(0) <= CNStageIntLLROutputS1xD(37)(5);
  VNStageIntLLRInputS1xD(16)(0) <= CNStageIntLLROutputS1xD(38)(0);
  VNStageIntLLRInputS1xD(80)(0) <= CNStageIntLLROutputS1xD(38)(1);
  VNStageIntLLRInputS1xD(144)(0) <= CNStageIntLLROutputS1xD(38)(2);
  VNStageIntLLRInputS1xD(208)(0) <= CNStageIntLLROutputS1xD(38)(3);
  VNStageIntLLRInputS1xD(272)(0) <= CNStageIntLLROutputS1xD(38)(4);
  VNStageIntLLRInputS1xD(336)(0) <= CNStageIntLLROutputS1xD(38)(5);
  VNStageIntLLRInputS1xD(15)(0) <= CNStageIntLLROutputS1xD(39)(0);
  VNStageIntLLRInputS1xD(79)(0) <= CNStageIntLLROutputS1xD(39)(1);
  VNStageIntLLRInputS1xD(143)(0) <= CNStageIntLLROutputS1xD(39)(2);
  VNStageIntLLRInputS1xD(207)(0) <= CNStageIntLLROutputS1xD(39)(3);
  VNStageIntLLRInputS1xD(271)(0) <= CNStageIntLLROutputS1xD(39)(4);
  VNStageIntLLRInputS1xD(335)(0) <= CNStageIntLLROutputS1xD(39)(5);
  VNStageIntLLRInputS1xD(14)(0) <= CNStageIntLLROutputS1xD(40)(0);
  VNStageIntLLRInputS1xD(78)(0) <= CNStageIntLLROutputS1xD(40)(1);
  VNStageIntLLRInputS1xD(142)(0) <= CNStageIntLLROutputS1xD(40)(2);
  VNStageIntLLRInputS1xD(206)(0) <= CNStageIntLLROutputS1xD(40)(3);
  VNStageIntLLRInputS1xD(270)(0) <= CNStageIntLLROutputS1xD(40)(4);
  VNStageIntLLRInputS1xD(334)(0) <= CNStageIntLLROutputS1xD(40)(5);
  VNStageIntLLRInputS1xD(12)(0) <= CNStageIntLLROutputS1xD(41)(0);
  VNStageIntLLRInputS1xD(76)(0) <= CNStageIntLLROutputS1xD(41)(1);
  VNStageIntLLRInputS1xD(140)(0) <= CNStageIntLLROutputS1xD(41)(2);
  VNStageIntLLRInputS1xD(204)(0) <= CNStageIntLLROutputS1xD(41)(3);
  VNStageIntLLRInputS1xD(268)(0) <= CNStageIntLLROutputS1xD(41)(4);
  VNStageIntLLRInputS1xD(332)(0) <= CNStageIntLLROutputS1xD(41)(5);
  VNStageIntLLRInputS1xD(11)(0) <= CNStageIntLLROutputS1xD(42)(0);
  VNStageIntLLRInputS1xD(75)(0) <= CNStageIntLLROutputS1xD(42)(1);
  VNStageIntLLRInputS1xD(139)(0) <= CNStageIntLLROutputS1xD(42)(2);
  VNStageIntLLRInputS1xD(203)(0) <= CNStageIntLLROutputS1xD(42)(3);
  VNStageIntLLRInputS1xD(267)(0) <= CNStageIntLLROutputS1xD(42)(4);
  VNStageIntLLRInputS1xD(331)(0) <= CNStageIntLLROutputS1xD(42)(5);
  VNStageIntLLRInputS1xD(10)(0) <= CNStageIntLLROutputS1xD(43)(0);
  VNStageIntLLRInputS1xD(74)(0) <= CNStageIntLLROutputS1xD(43)(1);
  VNStageIntLLRInputS1xD(138)(0) <= CNStageIntLLROutputS1xD(43)(2);
  VNStageIntLLRInputS1xD(202)(0) <= CNStageIntLLROutputS1xD(43)(3);
  VNStageIntLLRInputS1xD(266)(0) <= CNStageIntLLROutputS1xD(43)(4);
  VNStageIntLLRInputS1xD(330)(0) <= CNStageIntLLROutputS1xD(43)(5);
  VNStageIntLLRInputS1xD(9)(0) <= CNStageIntLLROutputS1xD(44)(0);
  VNStageIntLLRInputS1xD(73)(0) <= CNStageIntLLROutputS1xD(44)(1);
  VNStageIntLLRInputS1xD(137)(0) <= CNStageIntLLROutputS1xD(44)(2);
  VNStageIntLLRInputS1xD(201)(0) <= CNStageIntLLROutputS1xD(44)(3);
  VNStageIntLLRInputS1xD(265)(0) <= CNStageIntLLROutputS1xD(44)(4);
  VNStageIntLLRInputS1xD(329)(0) <= CNStageIntLLROutputS1xD(44)(5);
  VNStageIntLLRInputS1xD(8)(0) <= CNStageIntLLROutputS1xD(45)(0);
  VNStageIntLLRInputS1xD(72)(0) <= CNStageIntLLROutputS1xD(45)(1);
  VNStageIntLLRInputS1xD(136)(0) <= CNStageIntLLROutputS1xD(45)(2);
  VNStageIntLLRInputS1xD(200)(0) <= CNStageIntLLROutputS1xD(45)(3);
  VNStageIntLLRInputS1xD(264)(0) <= CNStageIntLLROutputS1xD(45)(4);
  VNStageIntLLRInputS1xD(328)(0) <= CNStageIntLLROutputS1xD(45)(5);
  VNStageIntLLRInputS1xD(7)(0) <= CNStageIntLLROutputS1xD(46)(0);
  VNStageIntLLRInputS1xD(71)(0) <= CNStageIntLLROutputS1xD(46)(1);
  VNStageIntLLRInputS1xD(135)(0) <= CNStageIntLLROutputS1xD(46)(2);
  VNStageIntLLRInputS1xD(199)(0) <= CNStageIntLLROutputS1xD(46)(3);
  VNStageIntLLRInputS1xD(263)(0) <= CNStageIntLLROutputS1xD(46)(4);
  VNStageIntLLRInputS1xD(327)(0) <= CNStageIntLLROutputS1xD(46)(5);
  VNStageIntLLRInputS1xD(6)(0) <= CNStageIntLLROutputS1xD(47)(0);
  VNStageIntLLRInputS1xD(70)(0) <= CNStageIntLLROutputS1xD(47)(1);
  VNStageIntLLRInputS1xD(134)(0) <= CNStageIntLLROutputS1xD(47)(2);
  VNStageIntLLRInputS1xD(198)(0) <= CNStageIntLLROutputS1xD(47)(3);
  VNStageIntLLRInputS1xD(262)(0) <= CNStageIntLLROutputS1xD(47)(4);
  VNStageIntLLRInputS1xD(326)(0) <= CNStageIntLLROutputS1xD(47)(5);
  VNStageIntLLRInputS1xD(5)(0) <= CNStageIntLLROutputS1xD(48)(0);
  VNStageIntLLRInputS1xD(69)(0) <= CNStageIntLLROutputS1xD(48)(1);
  VNStageIntLLRInputS1xD(133)(0) <= CNStageIntLLROutputS1xD(48)(2);
  VNStageIntLLRInputS1xD(197)(0) <= CNStageIntLLROutputS1xD(48)(3);
  VNStageIntLLRInputS1xD(261)(0) <= CNStageIntLLROutputS1xD(48)(4);
  VNStageIntLLRInputS1xD(325)(0) <= CNStageIntLLROutputS1xD(48)(5);
  VNStageIntLLRInputS1xD(4)(0) <= CNStageIntLLROutputS1xD(49)(0);
  VNStageIntLLRInputS1xD(68)(0) <= CNStageIntLLROutputS1xD(49)(1);
  VNStageIntLLRInputS1xD(132)(0) <= CNStageIntLLROutputS1xD(49)(2);
  VNStageIntLLRInputS1xD(196)(0) <= CNStageIntLLROutputS1xD(49)(3);
  VNStageIntLLRInputS1xD(260)(0) <= CNStageIntLLROutputS1xD(49)(4);
  VNStageIntLLRInputS1xD(324)(0) <= CNStageIntLLROutputS1xD(49)(5);
  VNStageIntLLRInputS1xD(2)(0) <= CNStageIntLLROutputS1xD(50)(0);
  VNStageIntLLRInputS1xD(66)(0) <= CNStageIntLLROutputS1xD(50)(1);
  VNStageIntLLRInputS1xD(130)(0) <= CNStageIntLLROutputS1xD(50)(2);
  VNStageIntLLRInputS1xD(194)(0) <= CNStageIntLLROutputS1xD(50)(3);
  VNStageIntLLRInputS1xD(258)(0) <= CNStageIntLLROutputS1xD(50)(4);
  VNStageIntLLRInputS1xD(322)(0) <= CNStageIntLLROutputS1xD(50)(5);
  VNStageIntLLRInputS1xD(1)(0) <= CNStageIntLLROutputS1xD(51)(0);
  VNStageIntLLRInputS1xD(65)(0) <= CNStageIntLLROutputS1xD(51)(1);
  VNStageIntLLRInputS1xD(129)(0) <= CNStageIntLLROutputS1xD(51)(2);
  VNStageIntLLRInputS1xD(193)(0) <= CNStageIntLLROutputS1xD(51)(3);
  VNStageIntLLRInputS1xD(257)(0) <= CNStageIntLLROutputS1xD(51)(4);
  VNStageIntLLRInputS1xD(321)(0) <= CNStageIntLLROutputS1xD(51)(5);
  VNStageIntLLRInputS1xD(63)(0) <= CNStageIntLLROutputS1xD(52)(0);
  VNStageIntLLRInputS1xD(127)(0) <= CNStageIntLLROutputS1xD(52)(1);
  VNStageIntLLRInputS1xD(191)(0) <= CNStageIntLLROutputS1xD(52)(2);
  VNStageIntLLRInputS1xD(255)(0) <= CNStageIntLLROutputS1xD(52)(3);
  VNStageIntLLRInputS1xD(319)(0) <= CNStageIntLLROutputS1xD(52)(4);
  VNStageIntLLRInputS1xD(383)(0) <= CNStageIntLLROutputS1xD(52)(5);
  VNStageIntLLRInputS1xD(0)(0) <= CNStageIntLLROutputS1xD(53)(0);
  VNStageIntLLRInputS1xD(64)(0) <= CNStageIntLLROutputS1xD(53)(1);
  VNStageIntLLRInputS1xD(128)(0) <= CNStageIntLLROutputS1xD(53)(2);
  VNStageIntLLRInputS1xD(192)(0) <= CNStageIntLLROutputS1xD(53)(3);
  VNStageIntLLRInputS1xD(256)(0) <= CNStageIntLLROutputS1xD(53)(4);
  VNStageIntLLRInputS1xD(320)(0) <= CNStageIntLLROutputS1xD(53)(5);
  VNStageIntLLRInputS1xD(42)(1) <= CNStageIntLLROutputS1xD(54)(0);
  VNStageIntLLRInputS1xD(112)(1) <= CNStageIntLLROutputS1xD(54)(1);
  VNStageIntLLRInputS1xD(182)(1) <= CNStageIntLLROutputS1xD(54)(2);
  VNStageIntLLRInputS1xD(203)(1) <= CNStageIntLLROutputS1xD(54)(3);
  VNStageIntLLRInputS1xD(259)(0) <= CNStageIntLLROutputS1xD(54)(4);
  VNStageIntLLRInputS1xD(361)(1) <= CNStageIntLLROutputS1xD(54)(5);
  VNStageIntLLRInputS1xD(41)(1) <= CNStageIntLLROutputS1xD(55)(0);
  VNStageIntLLRInputS1xD(117)(1) <= CNStageIntLLROutputS1xD(55)(1);
  VNStageIntLLRInputS1xD(138)(1) <= CNStageIntLLROutputS1xD(55)(2);
  VNStageIntLLRInputS1xD(194)(1) <= CNStageIntLLROutputS1xD(55)(3);
  VNStageIntLLRInputS1xD(296)(1) <= CNStageIntLLROutputS1xD(55)(4);
  VNStageIntLLRInputS1xD(362)(1) <= CNStageIntLLROutputS1xD(55)(5);
  VNStageIntLLRInputS1xD(40)(1) <= CNStageIntLLROutputS1xD(56)(0);
  VNStageIntLLRInputS1xD(73)(1) <= CNStageIntLLROutputS1xD(56)(1);
  VNStageIntLLRInputS1xD(129)(1) <= CNStageIntLLROutputS1xD(56)(2);
  VNStageIntLLRInputS1xD(231)(1) <= CNStageIntLLROutputS1xD(56)(3);
  VNStageIntLLRInputS1xD(297)(1) <= CNStageIntLLROutputS1xD(56)(4);
  VNStageIntLLRInputS1xD(323)(0) <= CNStageIntLLROutputS1xD(56)(5);
  VNStageIntLLRInputS1xD(39)(1) <= CNStageIntLLROutputS1xD(57)(0);
  VNStageIntLLRInputS1xD(127)(1) <= CNStageIntLLROutputS1xD(57)(1);
  VNStageIntLLRInputS1xD(166)(1) <= CNStageIntLLROutputS1xD(57)(2);
  VNStageIntLLRInputS1xD(232)(1) <= CNStageIntLLROutputS1xD(57)(3);
  VNStageIntLLRInputS1xD(258)(1) <= CNStageIntLLROutputS1xD(57)(4);
  VNStageIntLLRInputS1xD(344)(1) <= CNStageIntLLROutputS1xD(57)(5);
  VNStageIntLLRInputS1xD(38)(1) <= CNStageIntLLROutputS1xD(58)(0);
  VNStageIntLLRInputS1xD(101)(1) <= CNStageIntLLROutputS1xD(58)(1);
  VNStageIntLLRInputS1xD(167)(1) <= CNStageIntLLROutputS1xD(58)(2);
  VNStageIntLLRInputS1xD(193)(1) <= CNStageIntLLROutputS1xD(58)(3);
  VNStageIntLLRInputS1xD(279)(1) <= CNStageIntLLROutputS1xD(58)(4);
  VNStageIntLLRInputS1xD(340)(1) <= CNStageIntLLROutputS1xD(58)(5);
  VNStageIntLLRInputS1xD(37)(1) <= CNStageIntLLROutputS1xD(59)(0);
  VNStageIntLLRInputS1xD(102)(1) <= CNStageIntLLROutputS1xD(59)(1);
  VNStageIntLLRInputS1xD(191)(1) <= CNStageIntLLROutputS1xD(59)(2);
  VNStageIntLLRInputS1xD(214)(1) <= CNStageIntLLROutputS1xD(59)(3);
  VNStageIntLLRInputS1xD(275)(1) <= CNStageIntLLROutputS1xD(59)(4);
  VNStageIntLLRInputS1xD(355)(1) <= CNStageIntLLROutputS1xD(59)(5);
  VNStageIntLLRInputS1xD(36)(1) <= CNStageIntLLROutputS1xD(60)(0);
  VNStageIntLLRInputS1xD(126)(0) <= CNStageIntLLROutputS1xD(60)(1);
  VNStageIntLLRInputS1xD(149)(1) <= CNStageIntLLROutputS1xD(60)(2);
  VNStageIntLLRInputS1xD(210)(1) <= CNStageIntLLROutputS1xD(60)(3);
  VNStageIntLLRInputS1xD(290)(1) <= CNStageIntLLROutputS1xD(60)(4);
  VNStageIntLLRInputS1xD(381)(0) <= CNStageIntLLROutputS1xD(60)(5);
  VNStageIntLLRInputS1xD(35)(1) <= CNStageIntLLROutputS1xD(61)(0);
  VNStageIntLLRInputS1xD(84)(1) <= CNStageIntLLROutputS1xD(61)(1);
  VNStageIntLLRInputS1xD(145)(1) <= CNStageIntLLROutputS1xD(61)(2);
  VNStageIntLLRInputS1xD(225)(1) <= CNStageIntLLROutputS1xD(61)(3);
  VNStageIntLLRInputS1xD(316)(0) <= CNStageIntLLROutputS1xD(61)(4);
  VNStageIntLLRInputS1xD(357)(1) <= CNStageIntLLROutputS1xD(61)(5);
  VNStageIntLLRInputS1xD(34)(1) <= CNStageIntLLROutputS1xD(62)(0);
  VNStageIntLLRInputS1xD(80)(1) <= CNStageIntLLROutputS1xD(62)(1);
  VNStageIntLLRInputS1xD(160)(1) <= CNStageIntLLROutputS1xD(62)(2);
  VNStageIntLLRInputS1xD(251)(0) <= CNStageIntLLROutputS1xD(62)(3);
  VNStageIntLLRInputS1xD(292)(1) <= CNStageIntLLROutputS1xD(62)(4);
  VNStageIntLLRInputS1xD(326)(1) <= CNStageIntLLROutputS1xD(62)(5);
  VNStageIntLLRInputS1xD(33)(1) <= CNStageIntLLROutputS1xD(63)(0);
  VNStageIntLLRInputS1xD(95)(1) <= CNStageIntLLROutputS1xD(63)(1);
  VNStageIntLLRInputS1xD(186)(0) <= CNStageIntLLROutputS1xD(63)(2);
  VNStageIntLLRInputS1xD(227)(1) <= CNStageIntLLROutputS1xD(63)(3);
  VNStageIntLLRInputS1xD(261)(1) <= CNStageIntLLROutputS1xD(63)(4);
  VNStageIntLLRInputS1xD(342)(1) <= CNStageIntLLROutputS1xD(63)(5);
  VNStageIntLLRInputS1xD(32)(1) <= CNStageIntLLROutputS1xD(64)(0);
  VNStageIntLLRInputS1xD(121)(0) <= CNStageIntLLROutputS1xD(64)(1);
  VNStageIntLLRInputS1xD(162)(1) <= CNStageIntLLROutputS1xD(64)(2);
  VNStageIntLLRInputS1xD(196)(1) <= CNStageIntLLROutputS1xD(64)(3);
  VNStageIntLLRInputS1xD(277)(1) <= CNStageIntLLROutputS1xD(64)(4);
  VNStageIntLLRInputS1xD(375)(1) <= CNStageIntLLROutputS1xD(64)(5);
  VNStageIntLLRInputS1xD(31)(1) <= CNStageIntLLROutputS1xD(65)(0);
  VNStageIntLLRInputS1xD(97)(1) <= CNStageIntLLROutputS1xD(65)(1);
  VNStageIntLLRInputS1xD(131)(0) <= CNStageIntLLROutputS1xD(65)(2);
  VNStageIntLLRInputS1xD(212)(1) <= CNStageIntLLROutputS1xD(65)(3);
  VNStageIntLLRInputS1xD(310)(1) <= CNStageIntLLROutputS1xD(65)(4);
  VNStageIntLLRInputS1xD(321)(1) <= CNStageIntLLROutputS1xD(65)(5);
  VNStageIntLLRInputS1xD(30)(1) <= CNStageIntLLROutputS1xD(66)(0);
  VNStageIntLLRInputS1xD(66)(1) <= CNStageIntLLROutputS1xD(66)(1);
  VNStageIntLLRInputS1xD(147)(1) <= CNStageIntLLROutputS1xD(66)(2);
  VNStageIntLLRInputS1xD(245)(1) <= CNStageIntLLROutputS1xD(66)(3);
  VNStageIntLLRInputS1xD(319)(1) <= CNStageIntLLROutputS1xD(66)(4);
  VNStageIntLLRInputS1xD(334)(1) <= CNStageIntLLROutputS1xD(66)(5);
  VNStageIntLLRInputS1xD(29)(1) <= CNStageIntLLROutputS1xD(67)(0);
  VNStageIntLLRInputS1xD(82)(1) <= CNStageIntLLROutputS1xD(67)(1);
  VNStageIntLLRInputS1xD(180)(0) <= CNStageIntLLROutputS1xD(67)(2);
  VNStageIntLLRInputS1xD(254)(0) <= CNStageIntLLROutputS1xD(67)(3);
  VNStageIntLLRInputS1xD(269)(0) <= CNStageIntLLROutputS1xD(67)(4);
  VNStageIntLLRInputS1xD(376)(1) <= CNStageIntLLROutputS1xD(67)(5);
  VNStageIntLLRInputS1xD(28)(1) <= CNStageIntLLROutputS1xD(68)(0);
  VNStageIntLLRInputS1xD(115)(1) <= CNStageIntLLROutputS1xD(68)(1);
  VNStageIntLLRInputS1xD(189)(0) <= CNStageIntLLROutputS1xD(68)(2);
  VNStageIntLLRInputS1xD(204)(1) <= CNStageIntLLROutputS1xD(68)(3);
  VNStageIntLLRInputS1xD(311)(1) <= CNStageIntLLROutputS1xD(68)(4);
  VNStageIntLLRInputS1xD(341)(1) <= CNStageIntLLROutputS1xD(68)(5);
  VNStageIntLLRInputS1xD(27)(1) <= CNStageIntLLROutputS1xD(69)(0);
  VNStageIntLLRInputS1xD(124)(0) <= CNStageIntLLROutputS1xD(69)(1);
  VNStageIntLLRInputS1xD(139)(1) <= CNStageIntLLROutputS1xD(69)(2);
  VNStageIntLLRInputS1xD(246)(1) <= CNStageIntLLROutputS1xD(69)(3);
  VNStageIntLLRInputS1xD(276)(1) <= CNStageIntLLROutputS1xD(69)(4);
  VNStageIntLLRInputS1xD(343)(1) <= CNStageIntLLROutputS1xD(69)(5);
  VNStageIntLLRInputS1xD(26)(1) <= CNStageIntLLROutputS1xD(70)(0);
  VNStageIntLLRInputS1xD(74)(1) <= CNStageIntLLROutputS1xD(70)(1);
  VNStageIntLLRInputS1xD(181)(1) <= CNStageIntLLROutputS1xD(70)(2);
  VNStageIntLLRInputS1xD(211)(1) <= CNStageIntLLROutputS1xD(70)(3);
  VNStageIntLLRInputS1xD(278)(1) <= CNStageIntLLROutputS1xD(70)(4);
  VNStageIntLLRInputS1xD(325)(1) <= CNStageIntLLROutputS1xD(70)(5);
  VNStageIntLLRInputS1xD(25)(1) <= CNStageIntLLROutputS1xD(71)(0);
  VNStageIntLLRInputS1xD(116)(0) <= CNStageIntLLROutputS1xD(71)(1);
  VNStageIntLLRInputS1xD(146)(1) <= CNStageIntLLROutputS1xD(71)(2);
  VNStageIntLLRInputS1xD(213)(1) <= CNStageIntLLROutputS1xD(71)(3);
  VNStageIntLLRInputS1xD(260)(1) <= CNStageIntLLROutputS1xD(71)(4);
  VNStageIntLLRInputS1xD(332)(1) <= CNStageIntLLROutputS1xD(71)(5);
  VNStageIntLLRInputS1xD(24)(1) <= CNStageIntLLROutputS1xD(72)(0);
  VNStageIntLLRInputS1xD(81)(1) <= CNStageIntLLROutputS1xD(72)(1);
  VNStageIntLLRInputS1xD(148)(1) <= CNStageIntLLROutputS1xD(72)(2);
  VNStageIntLLRInputS1xD(195)(0) <= CNStageIntLLROutputS1xD(72)(3);
  VNStageIntLLRInputS1xD(267)(1) <= CNStageIntLLROutputS1xD(72)(4);
  VNStageIntLLRInputS1xD(359)(1) <= CNStageIntLLROutputS1xD(72)(5);
  VNStageIntLLRInputS1xD(23)(1) <= CNStageIntLLROutputS1xD(73)(0);
  VNStageIntLLRInputS1xD(83)(1) <= CNStageIntLLROutputS1xD(73)(1);
  VNStageIntLLRInputS1xD(130)(1) <= CNStageIntLLROutputS1xD(73)(2);
  VNStageIntLLRInputS1xD(202)(1) <= CNStageIntLLROutputS1xD(73)(3);
  VNStageIntLLRInputS1xD(294)(1) <= CNStageIntLLROutputS1xD(73)(4);
  VNStageIntLLRInputS1xD(347)(1) <= CNStageIntLLROutputS1xD(73)(5);
  VNStageIntLLRInputS1xD(22)(1) <= CNStageIntLLROutputS1xD(74)(0);
  VNStageIntLLRInputS1xD(65)(1) <= CNStageIntLLROutputS1xD(74)(1);
  VNStageIntLLRInputS1xD(137)(1) <= CNStageIntLLROutputS1xD(74)(2);
  VNStageIntLLRInputS1xD(229)(1) <= CNStageIntLLROutputS1xD(74)(3);
  VNStageIntLLRInputS1xD(282)(1) <= CNStageIntLLROutputS1xD(74)(4);
  VNStageIntLLRInputS1xD(353)(1) <= CNStageIntLLROutputS1xD(74)(5);
  VNStageIntLLRInputS1xD(21)(1) <= CNStageIntLLROutputS1xD(75)(0);
  VNStageIntLLRInputS1xD(72)(1) <= CNStageIntLLROutputS1xD(75)(1);
  VNStageIntLLRInputS1xD(164)(1) <= CNStageIntLLROutputS1xD(75)(2);
  VNStageIntLLRInputS1xD(217)(1) <= CNStageIntLLROutputS1xD(75)(3);
  VNStageIntLLRInputS1xD(288)(1) <= CNStageIntLLROutputS1xD(75)(4);
  VNStageIntLLRInputS1xD(348)(1) <= CNStageIntLLROutputS1xD(75)(5);
  VNStageIntLLRInputS1xD(20)(1) <= CNStageIntLLROutputS1xD(76)(0);
  VNStageIntLLRInputS1xD(99)(1) <= CNStageIntLLROutputS1xD(76)(1);
  VNStageIntLLRInputS1xD(152)(1) <= CNStageIntLLROutputS1xD(76)(2);
  VNStageIntLLRInputS1xD(223)(1) <= CNStageIntLLROutputS1xD(76)(3);
  VNStageIntLLRInputS1xD(283)(1) <= CNStageIntLLROutputS1xD(76)(4);
  VNStageIntLLRInputS1xD(358)(1) <= CNStageIntLLROutputS1xD(76)(5);
  VNStageIntLLRInputS1xD(19)(1) <= CNStageIntLLROutputS1xD(77)(0);
  VNStageIntLLRInputS1xD(87)(1) <= CNStageIntLLROutputS1xD(77)(1);
  VNStageIntLLRInputS1xD(158)(1) <= CNStageIntLLROutputS1xD(77)(2);
  VNStageIntLLRInputS1xD(218)(1) <= CNStageIntLLROutputS1xD(77)(3);
  VNStageIntLLRInputS1xD(293)(1) <= CNStageIntLLROutputS1xD(77)(4);
  VNStageIntLLRInputS1xD(380)(0) <= CNStageIntLLROutputS1xD(77)(5);
  VNStageIntLLRInputS1xD(18)(1) <= CNStageIntLLROutputS1xD(78)(0);
  VNStageIntLLRInputS1xD(93)(1) <= CNStageIntLLROutputS1xD(78)(1);
  VNStageIntLLRInputS1xD(153)(1) <= CNStageIntLLROutputS1xD(78)(2);
  VNStageIntLLRInputS1xD(228)(1) <= CNStageIntLLROutputS1xD(78)(3);
  VNStageIntLLRInputS1xD(315)(0) <= CNStageIntLLROutputS1xD(78)(4);
  VNStageIntLLRInputS1xD(335)(1) <= CNStageIntLLROutputS1xD(78)(5);
  VNStageIntLLRInputS1xD(17)(1) <= CNStageIntLLROutputS1xD(79)(0);
  VNStageIntLLRInputS1xD(88)(1) <= CNStageIntLLROutputS1xD(79)(1);
  VNStageIntLLRInputS1xD(163)(1) <= CNStageIntLLROutputS1xD(79)(2);
  VNStageIntLLRInputS1xD(250)(0) <= CNStageIntLLROutputS1xD(79)(3);
  VNStageIntLLRInputS1xD(270)(1) <= CNStageIntLLROutputS1xD(79)(4);
  VNStageIntLLRInputS1xD(383)(1) <= CNStageIntLLROutputS1xD(79)(5);
  VNStageIntLLRInputS1xD(15)(1) <= CNStageIntLLROutputS1xD(80)(0);
  VNStageIntLLRInputS1xD(120)(1) <= CNStageIntLLROutputS1xD(80)(1);
  VNStageIntLLRInputS1xD(140)(1) <= CNStageIntLLROutputS1xD(80)(2);
  VNStageIntLLRInputS1xD(253)(0) <= CNStageIntLLROutputS1xD(80)(3);
  VNStageIntLLRInputS1xD(305)(1) <= CNStageIntLLROutputS1xD(80)(4);
  VNStageIntLLRInputS1xD(338)(1) <= CNStageIntLLROutputS1xD(80)(5);
  VNStageIntLLRInputS1xD(14)(1) <= CNStageIntLLROutputS1xD(81)(0);
  VNStageIntLLRInputS1xD(75)(1) <= CNStageIntLLROutputS1xD(81)(1);
  VNStageIntLLRInputS1xD(188)(0) <= CNStageIntLLROutputS1xD(81)(2);
  VNStageIntLLRInputS1xD(240)(1) <= CNStageIntLLROutputS1xD(81)(3);
  VNStageIntLLRInputS1xD(273)(1) <= CNStageIntLLROutputS1xD(81)(4);
  VNStageIntLLRInputS1xD(350)(1) <= CNStageIntLLROutputS1xD(81)(5);
  VNStageIntLLRInputS1xD(13)(0) <= CNStageIntLLROutputS1xD(82)(0);
  VNStageIntLLRInputS1xD(123)(0) <= CNStageIntLLROutputS1xD(82)(1);
  VNStageIntLLRInputS1xD(175)(1) <= CNStageIntLLROutputS1xD(82)(2);
  VNStageIntLLRInputS1xD(208)(1) <= CNStageIntLLROutputS1xD(82)(3);
  VNStageIntLLRInputS1xD(285)(1) <= CNStageIntLLROutputS1xD(82)(4);
  VNStageIntLLRInputS1xD(364)(1) <= CNStageIntLLROutputS1xD(82)(5);
  VNStageIntLLRInputS1xD(12)(1) <= CNStageIntLLROutputS1xD(83)(0);
  VNStageIntLLRInputS1xD(110)(1) <= CNStageIntLLROutputS1xD(83)(1);
  VNStageIntLLRInputS1xD(143)(1) <= CNStageIntLLROutputS1xD(83)(2);
  VNStageIntLLRInputS1xD(220)(1) <= CNStageIntLLROutputS1xD(83)(3);
  VNStageIntLLRInputS1xD(299)(0) <= CNStageIntLLROutputS1xD(83)(4);
  VNStageIntLLRInputS1xD(345)(1) <= CNStageIntLLROutputS1xD(83)(5);
  VNStageIntLLRInputS1xD(11)(1) <= CNStageIntLLROutputS1xD(84)(0);
  VNStageIntLLRInputS1xD(78)(1) <= CNStageIntLLROutputS1xD(84)(1);
  VNStageIntLLRInputS1xD(155)(1) <= CNStageIntLLROutputS1xD(84)(2);
  VNStageIntLLRInputS1xD(234)(1) <= CNStageIntLLROutputS1xD(84)(3);
  VNStageIntLLRInputS1xD(280)(1) <= CNStageIntLLROutputS1xD(84)(4);
  VNStageIntLLRInputS1xD(322)(1) <= CNStageIntLLROutputS1xD(84)(5);
  VNStageIntLLRInputS1xD(10)(1) <= CNStageIntLLROutputS1xD(85)(0);
  VNStageIntLLRInputS1xD(90)(1) <= CNStageIntLLROutputS1xD(85)(1);
  VNStageIntLLRInputS1xD(169)(1) <= CNStageIntLLROutputS1xD(85)(2);
  VNStageIntLLRInputS1xD(215)(1) <= CNStageIntLLROutputS1xD(85)(3);
  VNStageIntLLRInputS1xD(257)(1) <= CNStageIntLLROutputS1xD(85)(4);
  VNStageIntLLRInputS1xD(374)(1) <= CNStageIntLLROutputS1xD(85)(5);
  VNStageIntLLRInputS1xD(9)(1) <= CNStageIntLLROutputS1xD(86)(0);
  VNStageIntLLRInputS1xD(104)(1) <= CNStageIntLLROutputS1xD(86)(1);
  VNStageIntLLRInputS1xD(150)(1) <= CNStageIntLLROutputS1xD(86)(2);
  VNStageIntLLRInputS1xD(255)(1) <= CNStageIntLLROutputS1xD(86)(3);
  VNStageIntLLRInputS1xD(309)(1) <= CNStageIntLLROutputS1xD(86)(4);
  VNStageIntLLRInputS1xD(378)(0) <= CNStageIntLLROutputS1xD(86)(5);
  VNStageIntLLRInputS1xD(7)(1) <= CNStageIntLLROutputS1xD(87)(0);
  VNStageIntLLRInputS1xD(125)(0) <= CNStageIntLLROutputS1xD(87)(1);
  VNStageIntLLRInputS1xD(179)(1) <= CNStageIntLLROutputS1xD(87)(2);
  VNStageIntLLRInputS1xD(248)(1) <= CNStageIntLLROutputS1xD(87)(3);
  VNStageIntLLRInputS1xD(306)(1) <= CNStageIntLLROutputS1xD(87)(4);
  VNStageIntLLRInputS1xD(382)(0) <= CNStageIntLLROutputS1xD(87)(5);
  VNStageIntLLRInputS1xD(6)(1) <= CNStageIntLLROutputS1xD(88)(0);
  VNStageIntLLRInputS1xD(114)(1) <= CNStageIntLLROutputS1xD(88)(1);
  VNStageIntLLRInputS1xD(183)(1) <= CNStageIntLLROutputS1xD(88)(2);
  VNStageIntLLRInputS1xD(241)(1) <= CNStageIntLLROutputS1xD(88)(3);
  VNStageIntLLRInputS1xD(317)(0) <= CNStageIntLLROutputS1xD(88)(4);
  VNStageIntLLRInputS1xD(354)(1) <= CNStageIntLLROutputS1xD(88)(5);
  VNStageIntLLRInputS1xD(5)(1) <= CNStageIntLLROutputS1xD(89)(0);
  VNStageIntLLRInputS1xD(118)(1) <= CNStageIntLLROutputS1xD(89)(1);
  VNStageIntLLRInputS1xD(176)(1) <= CNStageIntLLROutputS1xD(89)(2);
  VNStageIntLLRInputS1xD(252)(0) <= CNStageIntLLROutputS1xD(89)(3);
  VNStageIntLLRInputS1xD(289)(1) <= CNStageIntLLROutputS1xD(89)(4);
  VNStageIntLLRInputS1xD(346)(1) <= CNStageIntLLROutputS1xD(89)(5);
  VNStageIntLLRInputS1xD(4)(1) <= CNStageIntLLROutputS1xD(90)(0);
  VNStageIntLLRInputS1xD(111)(1) <= CNStageIntLLROutputS1xD(90)(1);
  VNStageIntLLRInputS1xD(187)(0) <= CNStageIntLLROutputS1xD(90)(2);
  VNStageIntLLRInputS1xD(224)(1) <= CNStageIntLLROutputS1xD(90)(3);
  VNStageIntLLRInputS1xD(281)(1) <= CNStageIntLLROutputS1xD(90)(4);
  VNStageIntLLRInputS1xD(363)(0) <= CNStageIntLLROutputS1xD(90)(5);
  VNStageIntLLRInputS1xD(3)(0) <= CNStageIntLLROutputS1xD(91)(0);
  VNStageIntLLRInputS1xD(122)(0) <= CNStageIntLLROutputS1xD(91)(1);
  VNStageIntLLRInputS1xD(159)(1) <= CNStageIntLLROutputS1xD(91)(2);
  VNStageIntLLRInputS1xD(216)(1) <= CNStageIntLLROutputS1xD(91)(3);
  VNStageIntLLRInputS1xD(298)(1) <= CNStageIntLLROutputS1xD(91)(4);
  VNStageIntLLRInputS1xD(360)(1) <= CNStageIntLLROutputS1xD(91)(5);
  VNStageIntLLRInputS1xD(2)(1) <= CNStageIntLLROutputS1xD(92)(0);
  VNStageIntLLRInputS1xD(94)(1) <= CNStageIntLLROutputS1xD(92)(1);
  VNStageIntLLRInputS1xD(151)(1) <= CNStageIntLLROutputS1xD(92)(2);
  VNStageIntLLRInputS1xD(233)(1) <= CNStageIntLLROutputS1xD(92)(3);
  VNStageIntLLRInputS1xD(295)(1) <= CNStageIntLLROutputS1xD(92)(4);
  VNStageIntLLRInputS1xD(331)(1) <= CNStageIntLLROutputS1xD(92)(5);
  VNStageIntLLRInputS1xD(63)(1) <= CNStageIntLLROutputS1xD(93)(0);
  VNStageIntLLRInputS1xD(103)(1) <= CNStageIntLLROutputS1xD(93)(1);
  VNStageIntLLRInputS1xD(165)(1) <= CNStageIntLLROutputS1xD(93)(2);
  VNStageIntLLRInputS1xD(201)(1) <= CNStageIntLLROutputS1xD(93)(3);
  VNStageIntLLRInputS1xD(286)(1) <= CNStageIntLLROutputS1xD(93)(4);
  VNStageIntLLRInputS1xD(337)(1) <= CNStageIntLLROutputS1xD(93)(5);
  VNStageIntLLRInputS1xD(62)(0) <= CNStageIntLLROutputS1xD(94)(0);
  VNStageIntLLRInputS1xD(100)(1) <= CNStageIntLLROutputS1xD(94)(1);
  VNStageIntLLRInputS1xD(136)(1) <= CNStageIntLLROutputS1xD(94)(2);
  VNStageIntLLRInputS1xD(221)(1) <= CNStageIntLLROutputS1xD(94)(3);
  VNStageIntLLRInputS1xD(272)(1) <= CNStageIntLLROutputS1xD(94)(4);
  VNStageIntLLRInputS1xD(327)(1) <= CNStageIntLLROutputS1xD(94)(5);
  VNStageIntLLRInputS1xD(61)(0) <= CNStageIntLLROutputS1xD(95)(0);
  VNStageIntLLRInputS1xD(71)(1) <= CNStageIntLLROutputS1xD(95)(1);
  VNStageIntLLRInputS1xD(156)(1) <= CNStageIntLLROutputS1xD(95)(2);
  VNStageIntLLRInputS1xD(207)(1) <= CNStageIntLLROutputS1xD(95)(3);
  VNStageIntLLRInputS1xD(262)(1) <= CNStageIntLLROutputS1xD(95)(4);
  VNStageIntLLRInputS1xD(356)(1) <= CNStageIntLLROutputS1xD(95)(5);
  VNStageIntLLRInputS1xD(60)(0) <= CNStageIntLLROutputS1xD(96)(0);
  VNStageIntLLRInputS1xD(91)(1) <= CNStageIntLLROutputS1xD(96)(1);
  VNStageIntLLRInputS1xD(142)(1) <= CNStageIntLLROutputS1xD(96)(2);
  VNStageIntLLRInputS1xD(197)(1) <= CNStageIntLLROutputS1xD(96)(3);
  VNStageIntLLRInputS1xD(291)(1) <= CNStageIntLLROutputS1xD(96)(4);
  VNStageIntLLRInputS1xD(339)(1) <= CNStageIntLLROutputS1xD(96)(5);
  VNStageIntLLRInputS1xD(58)(0) <= CNStageIntLLROutputS1xD(97)(0);
  VNStageIntLLRInputS1xD(67)(0) <= CNStageIntLLROutputS1xD(97)(1);
  VNStageIntLLRInputS1xD(161)(1) <= CNStageIntLLROutputS1xD(97)(2);
  VNStageIntLLRInputS1xD(209)(1) <= CNStageIntLLROutputS1xD(97)(3);
  VNStageIntLLRInputS1xD(304)(1) <= CNStageIntLLROutputS1xD(97)(4);
  VNStageIntLLRInputS1xD(329)(1) <= CNStageIntLLROutputS1xD(97)(5);
  VNStageIntLLRInputS1xD(57)(0) <= CNStageIntLLROutputS1xD(98)(0);
  VNStageIntLLRInputS1xD(96)(1) <= CNStageIntLLROutputS1xD(98)(1);
  VNStageIntLLRInputS1xD(144)(1) <= CNStageIntLLROutputS1xD(98)(2);
  VNStageIntLLRInputS1xD(239)(1) <= CNStageIntLLROutputS1xD(98)(3);
  VNStageIntLLRInputS1xD(264)(1) <= CNStageIntLLROutputS1xD(98)(4);
  VNStageIntLLRInputS1xD(365)(1) <= CNStageIntLLROutputS1xD(98)(5);
  VNStageIntLLRInputS1xD(56)(1) <= CNStageIntLLROutputS1xD(99)(0);
  VNStageIntLLRInputS1xD(79)(1) <= CNStageIntLLROutputS1xD(99)(1);
  VNStageIntLLRInputS1xD(174)(1) <= CNStageIntLLROutputS1xD(99)(2);
  VNStageIntLLRInputS1xD(199)(1) <= CNStageIntLLROutputS1xD(99)(3);
  VNStageIntLLRInputS1xD(300)(1) <= CNStageIntLLROutputS1xD(99)(4);
  VNStageIntLLRInputS1xD(349)(1) <= CNStageIntLLROutputS1xD(99)(5);
  VNStageIntLLRInputS1xD(55)(1) <= CNStageIntLLROutputS1xD(100)(0);
  VNStageIntLLRInputS1xD(109)(1) <= CNStageIntLLROutputS1xD(100)(1);
  VNStageIntLLRInputS1xD(134)(1) <= CNStageIntLLROutputS1xD(100)(2);
  VNStageIntLLRInputS1xD(235)(0) <= CNStageIntLLROutputS1xD(100)(3);
  VNStageIntLLRInputS1xD(284)(1) <= CNStageIntLLROutputS1xD(100)(4);
  VNStageIntLLRInputS1xD(352)(1) <= CNStageIntLLROutputS1xD(100)(5);
  VNStageIntLLRInputS1xD(54)(1) <= CNStageIntLLROutputS1xD(101)(0);
  VNStageIntLLRInputS1xD(69)(1) <= CNStageIntLLROutputS1xD(101)(1);
  VNStageIntLLRInputS1xD(170)(1) <= CNStageIntLLROutputS1xD(101)(2);
  VNStageIntLLRInputS1xD(219)(1) <= CNStageIntLLROutputS1xD(101)(3);
  VNStageIntLLRInputS1xD(287)(1) <= CNStageIntLLROutputS1xD(101)(4);
  VNStageIntLLRInputS1xD(330)(1) <= CNStageIntLLROutputS1xD(101)(5);
  VNStageIntLLRInputS1xD(52)(0) <= CNStageIntLLROutputS1xD(102)(0);
  VNStageIntLLRInputS1xD(89)(1) <= CNStageIntLLROutputS1xD(102)(1);
  VNStageIntLLRInputS1xD(157)(1) <= CNStageIntLLROutputS1xD(102)(2);
  VNStageIntLLRInputS1xD(200)(1) <= CNStageIntLLROutputS1xD(102)(3);
  VNStageIntLLRInputS1xD(303)(1) <= CNStageIntLLROutputS1xD(102)(4);
  VNStageIntLLRInputS1xD(366)(1) <= CNStageIntLLROutputS1xD(102)(5);
  VNStageIntLLRInputS1xD(51)(1) <= CNStageIntLLROutputS1xD(103)(0);
  VNStageIntLLRInputS1xD(92)(1) <= CNStageIntLLROutputS1xD(103)(1);
  VNStageIntLLRInputS1xD(135)(1) <= CNStageIntLLROutputS1xD(103)(2);
  VNStageIntLLRInputS1xD(238)(1) <= CNStageIntLLROutputS1xD(103)(3);
  VNStageIntLLRInputS1xD(301)(1) <= CNStageIntLLROutputS1xD(103)(4);
  VNStageIntLLRInputS1xD(328)(1) <= CNStageIntLLROutputS1xD(103)(5);
  VNStageIntLLRInputS1xD(50)(1) <= CNStageIntLLROutputS1xD(104)(0);
  VNStageIntLLRInputS1xD(70)(1) <= CNStageIntLLROutputS1xD(104)(1);
  VNStageIntLLRInputS1xD(173)(1) <= CNStageIntLLROutputS1xD(104)(2);
  VNStageIntLLRInputS1xD(236)(1) <= CNStageIntLLROutputS1xD(104)(3);
  VNStageIntLLRInputS1xD(263)(1) <= CNStageIntLLROutputS1xD(104)(4);
  VNStageIntLLRInputS1xD(336)(1) <= CNStageIntLLROutputS1xD(104)(5);
  VNStageIntLLRInputS1xD(49)(1) <= CNStageIntLLROutputS1xD(105)(0);
  VNStageIntLLRInputS1xD(108)(1) <= CNStageIntLLROutputS1xD(105)(1);
  VNStageIntLLRInputS1xD(171)(0) <= CNStageIntLLROutputS1xD(105)(2);
  VNStageIntLLRInputS1xD(198)(1) <= CNStageIntLLROutputS1xD(105)(3);
  VNStageIntLLRInputS1xD(271)(1) <= CNStageIntLLROutputS1xD(105)(4);
  VNStageIntLLRInputS1xD(379)(0) <= CNStageIntLLROutputS1xD(105)(5);
  VNStageIntLLRInputS1xD(46)(1) <= CNStageIntLLROutputS1xD(106)(0);
  VNStageIntLLRInputS1xD(76)(1) <= CNStageIntLLROutputS1xD(106)(1);
  VNStageIntLLRInputS1xD(184)(1) <= CNStageIntLLROutputS1xD(106)(2);
  VNStageIntLLRInputS1xD(243)(1) <= CNStageIntLLROutputS1xD(106)(3);
  VNStageIntLLRInputS1xD(256)(1) <= CNStageIntLLROutputS1xD(106)(4);
  VNStageIntLLRInputS1xD(372)(0) <= CNStageIntLLROutputS1xD(106)(5);
  VNStageIntLLRInputS1xD(45)(1) <= CNStageIntLLROutputS1xD(107)(0);
  VNStageIntLLRInputS1xD(119)(1) <= CNStageIntLLROutputS1xD(107)(1);
  VNStageIntLLRInputS1xD(178)(1) <= CNStageIntLLROutputS1xD(107)(2);
  VNStageIntLLRInputS1xD(192)(1) <= CNStageIntLLROutputS1xD(107)(3);
  VNStageIntLLRInputS1xD(307)(1) <= CNStageIntLLROutputS1xD(107)(4);
  VNStageIntLLRInputS1xD(377)(0) <= CNStageIntLLROutputS1xD(107)(5);
  VNStageIntLLRInputS1xD(44)(1) <= CNStageIntLLROutputS1xD(108)(0);
  VNStageIntLLRInputS1xD(113)(1) <= CNStageIntLLROutputS1xD(108)(1);
  VNStageIntLLRInputS1xD(128)(1) <= CNStageIntLLROutputS1xD(108)(2);
  VNStageIntLLRInputS1xD(242)(1) <= CNStageIntLLROutputS1xD(108)(3);
  VNStageIntLLRInputS1xD(312)(1) <= CNStageIntLLROutputS1xD(108)(4);
  VNStageIntLLRInputS1xD(333)(0) <= CNStageIntLLROutputS1xD(108)(5);
  VNStageIntLLRInputS1xD(43)(0) <= CNStageIntLLROutputS1xD(109)(0);
  VNStageIntLLRInputS1xD(64)(1) <= CNStageIntLLROutputS1xD(109)(1);
  VNStageIntLLRInputS1xD(177)(1) <= CNStageIntLLROutputS1xD(109)(2);
  VNStageIntLLRInputS1xD(247)(1) <= CNStageIntLLROutputS1xD(109)(3);
  VNStageIntLLRInputS1xD(268)(1) <= CNStageIntLLROutputS1xD(109)(4);
  VNStageIntLLRInputS1xD(324)(1) <= CNStageIntLLROutputS1xD(109)(5);
  VNStageIntLLRInputS1xD(0)(1) <= CNStageIntLLROutputS1xD(110)(0);
  VNStageIntLLRInputS1xD(107)(0) <= CNStageIntLLROutputS1xD(110)(1);
  VNStageIntLLRInputS1xD(172)(1) <= CNStageIntLLROutputS1xD(110)(2);
  VNStageIntLLRInputS1xD(237)(1) <= CNStageIntLLROutputS1xD(110)(3);
  VNStageIntLLRInputS1xD(302)(1) <= CNStageIntLLROutputS1xD(110)(4);
  VNStageIntLLRInputS1xD(367)(1) <= CNStageIntLLROutputS1xD(110)(5);
  VNStageIntLLRInputS1xD(32)(2) <= CNStageIntLLROutputS1xD(111)(0);
  VNStageIntLLRInputS1xD(117)(2) <= CNStageIntLLROutputS1xD(111)(1);
  VNStageIntLLRInputS1xD(136)(2) <= CNStageIntLLROutputS1xD(111)(2);
  VNStageIntLLRInputS1xD(198)(2) <= CNStageIntLLROutputS1xD(111)(3);
  VNStageIntLLRInputS1xD(297)(2) <= CNStageIntLLROutputS1xD(111)(4);
  VNStageIntLLRInputS1xD(382)(1) <= CNStageIntLLROutputS1xD(111)(5);
  VNStageIntLLRInputS1xD(30)(2) <= CNStageIntLLROutputS1xD(112)(0);
  VNStageIntLLRInputS1xD(68)(1) <= CNStageIntLLROutputS1xD(112)(1);
  VNStageIntLLRInputS1xD(167)(2) <= CNStageIntLLROutputS1xD(112)(2);
  VNStageIntLLRInputS1xD(252)(1) <= CNStageIntLLROutputS1xD(112)(3);
  VNStageIntLLRInputS1xD(303)(2) <= CNStageIntLLROutputS1xD(112)(4);
  VNStageIntLLRInputS1xD(358)(2) <= CNStageIntLLROutputS1xD(112)(5);
  VNStageIntLLRInputS1xD(29)(2) <= CNStageIntLLROutputS1xD(113)(0);
  VNStageIntLLRInputS1xD(102)(2) <= CNStageIntLLROutputS1xD(113)(1);
  VNStageIntLLRInputS1xD(187)(1) <= CNStageIntLLROutputS1xD(113)(2);
  VNStageIntLLRInputS1xD(238)(2) <= CNStageIntLLROutputS1xD(113)(3);
  VNStageIntLLRInputS1xD(293)(2) <= CNStageIntLLROutputS1xD(113)(4);
  VNStageIntLLRInputS1xD(324)(2) <= CNStageIntLLROutputS1xD(113)(5);
  VNStageIntLLRInputS1xD(28)(2) <= CNStageIntLLROutputS1xD(114)(0);
  VNStageIntLLRInputS1xD(122)(1) <= CNStageIntLLROutputS1xD(114)(1);
  VNStageIntLLRInputS1xD(173)(2) <= CNStageIntLLROutputS1xD(114)(2);
  VNStageIntLLRInputS1xD(228)(2) <= CNStageIntLLROutputS1xD(114)(3);
  VNStageIntLLRInputS1xD(259)(1) <= CNStageIntLLROutputS1xD(114)(4);
  VNStageIntLLRInputS1xD(370)(1) <= CNStageIntLLROutputS1xD(114)(5);
  VNStageIntLLRInputS1xD(27)(2) <= CNStageIntLLROutputS1xD(115)(0);
  VNStageIntLLRInputS1xD(108)(2) <= CNStageIntLLROutputS1xD(115)(1);
  VNStageIntLLRInputS1xD(163)(2) <= CNStageIntLLROutputS1xD(115)(2);
  VNStageIntLLRInputS1xD(194)(2) <= CNStageIntLLROutputS1xD(115)(3);
  VNStageIntLLRInputS1xD(305)(2) <= CNStageIntLLROutputS1xD(115)(4);
  VNStageIntLLRInputS1xD(337)(2) <= CNStageIntLLROutputS1xD(115)(5);
  VNStageIntLLRInputS1xD(26)(2) <= CNStageIntLLROutputS1xD(116)(0);
  VNStageIntLLRInputS1xD(98)(1) <= CNStageIntLLROutputS1xD(116)(1);
  VNStageIntLLRInputS1xD(129)(2) <= CNStageIntLLROutputS1xD(116)(2);
  VNStageIntLLRInputS1xD(240)(2) <= CNStageIntLLROutputS1xD(116)(3);
  VNStageIntLLRInputS1xD(272)(2) <= CNStageIntLLROutputS1xD(116)(4);
  VNStageIntLLRInputS1xD(360)(2) <= CNStageIntLLROutputS1xD(116)(5);
  VNStageIntLLRInputS1xD(25)(2) <= CNStageIntLLROutputS1xD(117)(0);
  VNStageIntLLRInputS1xD(127)(2) <= CNStageIntLLROutputS1xD(117)(1);
  VNStageIntLLRInputS1xD(175)(2) <= CNStageIntLLROutputS1xD(117)(2);
  VNStageIntLLRInputS1xD(207)(2) <= CNStageIntLLROutputS1xD(117)(3);
  VNStageIntLLRInputS1xD(295)(2) <= CNStageIntLLROutputS1xD(117)(4);
  VNStageIntLLRInputS1xD(333)(1) <= CNStageIntLLROutputS1xD(117)(5);
  VNStageIntLLRInputS1xD(24)(2) <= CNStageIntLLROutputS1xD(118)(0);
  VNStageIntLLRInputS1xD(110)(2) <= CNStageIntLLROutputS1xD(118)(1);
  VNStageIntLLRInputS1xD(142)(2) <= CNStageIntLLROutputS1xD(118)(2);
  VNStageIntLLRInputS1xD(230)(1) <= CNStageIntLLROutputS1xD(118)(3);
  VNStageIntLLRInputS1xD(268)(2) <= CNStageIntLLROutputS1xD(118)(4);
  VNStageIntLLRInputS1xD(380)(1) <= CNStageIntLLROutputS1xD(118)(5);
  VNStageIntLLRInputS1xD(23)(2) <= CNStageIntLLROutputS1xD(119)(0);
  VNStageIntLLRInputS1xD(77)(0) <= CNStageIntLLROutputS1xD(119)(1);
  VNStageIntLLRInputS1xD(165)(2) <= CNStageIntLLROutputS1xD(119)(2);
  VNStageIntLLRInputS1xD(203)(2) <= CNStageIntLLROutputS1xD(119)(3);
  VNStageIntLLRInputS1xD(315)(1) <= CNStageIntLLROutputS1xD(119)(4);
  VNStageIntLLRInputS1xD(383)(2) <= CNStageIntLLROutputS1xD(119)(5);
  VNStageIntLLRInputS1xD(22)(2) <= CNStageIntLLROutputS1xD(120)(0);
  VNStageIntLLRInputS1xD(100)(2) <= CNStageIntLLROutputS1xD(120)(1);
  VNStageIntLLRInputS1xD(138)(2) <= CNStageIntLLROutputS1xD(120)(2);
  VNStageIntLLRInputS1xD(250)(1) <= CNStageIntLLROutputS1xD(120)(3);
  VNStageIntLLRInputS1xD(318)(0) <= CNStageIntLLROutputS1xD(120)(4);
  VNStageIntLLRInputS1xD(361)(2) <= CNStageIntLLROutputS1xD(120)(5);
  VNStageIntLLRInputS1xD(21)(2) <= CNStageIntLLROutputS1xD(121)(0);
  VNStageIntLLRInputS1xD(73)(2) <= CNStageIntLLROutputS1xD(121)(1);
  VNStageIntLLRInputS1xD(185)(0) <= CNStageIntLLROutputS1xD(121)(2);
  VNStageIntLLRInputS1xD(253)(1) <= CNStageIntLLROutputS1xD(121)(3);
  VNStageIntLLRInputS1xD(296)(2) <= CNStageIntLLROutputS1xD(121)(4);
  VNStageIntLLRInputS1xD(336)(2) <= CNStageIntLLROutputS1xD(121)(5);
  VNStageIntLLRInputS1xD(19)(2) <= CNStageIntLLROutputS1xD(122)(0);
  VNStageIntLLRInputS1xD(123)(1) <= CNStageIntLLROutputS1xD(122)(1);
  VNStageIntLLRInputS1xD(166)(2) <= CNStageIntLLROutputS1xD(122)(2);
  VNStageIntLLRInputS1xD(206)(1) <= CNStageIntLLROutputS1xD(122)(3);
  VNStageIntLLRInputS1xD(269)(1) <= CNStageIntLLROutputS1xD(122)(4);
  VNStageIntLLRInputS1xD(359)(2) <= CNStageIntLLROutputS1xD(122)(5);
  VNStageIntLLRInputS1xD(18)(2) <= CNStageIntLLROutputS1xD(123)(0);
  VNStageIntLLRInputS1xD(101)(2) <= CNStageIntLLROutputS1xD(123)(1);
  VNStageIntLLRInputS1xD(141)(0) <= CNStageIntLLROutputS1xD(123)(2);
  VNStageIntLLRInputS1xD(204)(2) <= CNStageIntLLROutputS1xD(123)(3);
  VNStageIntLLRInputS1xD(294)(2) <= CNStageIntLLROutputS1xD(123)(4);
  VNStageIntLLRInputS1xD(367)(2) <= CNStageIntLLROutputS1xD(123)(5);
  VNStageIntLLRInputS1xD(17)(2) <= CNStageIntLLROutputS1xD(124)(0);
  VNStageIntLLRInputS1xD(76)(2) <= CNStageIntLLROutputS1xD(124)(1);
  VNStageIntLLRInputS1xD(139)(2) <= CNStageIntLLROutputS1xD(124)(2);
  VNStageIntLLRInputS1xD(229)(2) <= CNStageIntLLROutputS1xD(124)(3);
  VNStageIntLLRInputS1xD(302)(2) <= CNStageIntLLROutputS1xD(124)(4);
  VNStageIntLLRInputS1xD(347)(2) <= CNStageIntLLROutputS1xD(124)(5);
  VNStageIntLLRInputS1xD(16)(1) <= CNStageIntLLROutputS1xD(125)(0);
  VNStageIntLLRInputS1xD(74)(2) <= CNStageIntLLROutputS1xD(125)(1);
  VNStageIntLLRInputS1xD(164)(2) <= CNStageIntLLROutputS1xD(125)(2);
  VNStageIntLLRInputS1xD(237)(2) <= CNStageIntLLROutputS1xD(125)(3);
  VNStageIntLLRInputS1xD(282)(2) <= CNStageIntLLROutputS1xD(125)(4);
  VNStageIntLLRInputS1xD(341)(2) <= CNStageIntLLROutputS1xD(125)(5);
  VNStageIntLLRInputS1xD(15)(2) <= CNStageIntLLROutputS1xD(126)(0);
  VNStageIntLLRInputS1xD(99)(2) <= CNStageIntLLROutputS1xD(126)(1);
  VNStageIntLLRInputS1xD(172)(2) <= CNStageIntLLROutputS1xD(126)(2);
  VNStageIntLLRInputS1xD(217)(2) <= CNStageIntLLROutputS1xD(126)(3);
  VNStageIntLLRInputS1xD(276)(2) <= CNStageIntLLROutputS1xD(126)(4);
  VNStageIntLLRInputS1xD(320)(1) <= CNStageIntLLROutputS1xD(126)(5);
  VNStageIntLLRInputS1xD(14)(2) <= CNStageIntLLROutputS1xD(127)(0);
  VNStageIntLLRInputS1xD(107)(1) <= CNStageIntLLROutputS1xD(127)(1);
  VNStageIntLLRInputS1xD(152)(2) <= CNStageIntLLROutputS1xD(127)(2);
  VNStageIntLLRInputS1xD(211)(2) <= CNStageIntLLROutputS1xD(127)(3);
  VNStageIntLLRInputS1xD(256)(2) <= CNStageIntLLROutputS1xD(127)(4);
  VNStageIntLLRInputS1xD(340)(2) <= CNStageIntLLROutputS1xD(127)(5);
  VNStageIntLLRInputS1xD(13)(1) <= CNStageIntLLROutputS1xD(128)(0);
  VNStageIntLLRInputS1xD(87)(2) <= CNStageIntLLROutputS1xD(128)(1);
  VNStageIntLLRInputS1xD(146)(2) <= CNStageIntLLROutputS1xD(128)(2);
  VNStageIntLLRInputS1xD(192)(2) <= CNStageIntLLROutputS1xD(128)(3);
  VNStageIntLLRInputS1xD(275)(2) <= CNStageIntLLROutputS1xD(128)(4);
  VNStageIntLLRInputS1xD(345)(2) <= CNStageIntLLROutputS1xD(128)(5);
  VNStageIntLLRInputS1xD(12)(2) <= CNStageIntLLROutputS1xD(129)(0);
  VNStageIntLLRInputS1xD(81)(2) <= CNStageIntLLROutputS1xD(129)(1);
  VNStageIntLLRInputS1xD(128)(2) <= CNStageIntLLROutputS1xD(129)(2);
  VNStageIntLLRInputS1xD(210)(2) <= CNStageIntLLROutputS1xD(129)(3);
  VNStageIntLLRInputS1xD(280)(2) <= CNStageIntLLROutputS1xD(129)(4);
  VNStageIntLLRInputS1xD(364)(2) <= CNStageIntLLROutputS1xD(129)(5);
  VNStageIntLLRInputS1xD(11)(2) <= CNStageIntLLROutputS1xD(130)(0);
  VNStageIntLLRInputS1xD(64)(2) <= CNStageIntLLROutputS1xD(130)(1);
  VNStageIntLLRInputS1xD(145)(2) <= CNStageIntLLROutputS1xD(130)(2);
  VNStageIntLLRInputS1xD(215)(2) <= CNStageIntLLROutputS1xD(130)(3);
  VNStageIntLLRInputS1xD(299)(1) <= CNStageIntLLROutputS1xD(130)(4);
  VNStageIntLLRInputS1xD(355)(2) <= CNStageIntLLROutputS1xD(130)(5);
  VNStageIntLLRInputS1xD(10)(2) <= CNStageIntLLROutputS1xD(131)(0);
  VNStageIntLLRInputS1xD(80)(2) <= CNStageIntLLROutputS1xD(131)(1);
  VNStageIntLLRInputS1xD(150)(2) <= CNStageIntLLROutputS1xD(131)(2);
  VNStageIntLLRInputS1xD(234)(2) <= CNStageIntLLROutputS1xD(131)(3);
  VNStageIntLLRInputS1xD(290)(2) <= CNStageIntLLROutputS1xD(131)(4);
  VNStageIntLLRInputS1xD(329)(2) <= CNStageIntLLROutputS1xD(131)(5);
  VNStageIntLLRInputS1xD(9)(2) <= CNStageIntLLROutputS1xD(132)(0);
  VNStageIntLLRInputS1xD(85)(1) <= CNStageIntLLROutputS1xD(132)(1);
  VNStageIntLLRInputS1xD(169)(2) <= CNStageIntLLROutputS1xD(132)(2);
  VNStageIntLLRInputS1xD(225)(2) <= CNStageIntLLROutputS1xD(132)(3);
  VNStageIntLLRInputS1xD(264)(2) <= CNStageIntLLROutputS1xD(132)(4);
  VNStageIntLLRInputS1xD(330)(2) <= CNStageIntLLROutputS1xD(132)(5);
  VNStageIntLLRInputS1xD(8)(1) <= CNStageIntLLROutputS1xD(133)(0);
  VNStageIntLLRInputS1xD(104)(2) <= CNStageIntLLROutputS1xD(133)(1);
  VNStageIntLLRInputS1xD(160)(2) <= CNStageIntLLROutputS1xD(133)(2);
  VNStageIntLLRInputS1xD(199)(2) <= CNStageIntLLROutputS1xD(133)(3);
  VNStageIntLLRInputS1xD(265)(1) <= CNStageIntLLROutputS1xD(133)(4);
  VNStageIntLLRInputS1xD(354)(2) <= CNStageIntLLROutputS1xD(133)(5);
  VNStageIntLLRInputS1xD(7)(2) <= CNStageIntLLROutputS1xD(134)(0);
  VNStageIntLLRInputS1xD(95)(2) <= CNStageIntLLROutputS1xD(134)(1);
  VNStageIntLLRInputS1xD(134)(2) <= CNStageIntLLROutputS1xD(134)(2);
  VNStageIntLLRInputS1xD(200)(2) <= CNStageIntLLROutputS1xD(134)(3);
  VNStageIntLLRInputS1xD(289)(2) <= CNStageIntLLROutputS1xD(134)(4);
  VNStageIntLLRInputS1xD(375)(2) <= CNStageIntLLROutputS1xD(134)(5);
  VNStageIntLLRInputS1xD(6)(2) <= CNStageIntLLROutputS1xD(135)(0);
  VNStageIntLLRInputS1xD(69)(2) <= CNStageIntLLROutputS1xD(135)(1);
  VNStageIntLLRInputS1xD(135)(2) <= CNStageIntLLROutputS1xD(135)(2);
  VNStageIntLLRInputS1xD(224)(2) <= CNStageIntLLROutputS1xD(135)(3);
  VNStageIntLLRInputS1xD(310)(2) <= CNStageIntLLROutputS1xD(135)(4);
  VNStageIntLLRInputS1xD(371)(1) <= CNStageIntLLROutputS1xD(135)(5);
  VNStageIntLLRInputS1xD(5)(2) <= CNStageIntLLROutputS1xD(136)(0);
  VNStageIntLLRInputS1xD(70)(2) <= CNStageIntLLROutputS1xD(136)(1);
  VNStageIntLLRInputS1xD(159)(2) <= CNStageIntLLROutputS1xD(136)(2);
  VNStageIntLLRInputS1xD(245)(2) <= CNStageIntLLROutputS1xD(136)(3);
  VNStageIntLLRInputS1xD(306)(2) <= CNStageIntLLROutputS1xD(136)(4);
  VNStageIntLLRInputS1xD(323)(1) <= CNStageIntLLROutputS1xD(136)(5);
  VNStageIntLLRInputS1xD(3)(1) <= CNStageIntLLROutputS1xD(137)(0);
  VNStageIntLLRInputS1xD(115)(2) <= CNStageIntLLROutputS1xD(137)(1);
  VNStageIntLLRInputS1xD(176)(2) <= CNStageIntLLROutputS1xD(137)(2);
  VNStageIntLLRInputS1xD(193)(2) <= CNStageIntLLROutputS1xD(137)(3);
  VNStageIntLLRInputS1xD(284)(2) <= CNStageIntLLROutputS1xD(137)(4);
  VNStageIntLLRInputS1xD(325)(2) <= CNStageIntLLROutputS1xD(137)(5);
  VNStageIntLLRInputS1xD(2)(2) <= CNStageIntLLROutputS1xD(138)(0);
  VNStageIntLLRInputS1xD(111)(2) <= CNStageIntLLROutputS1xD(138)(1);
  VNStageIntLLRInputS1xD(191)(2) <= CNStageIntLLROutputS1xD(138)(2);
  VNStageIntLLRInputS1xD(219)(2) <= CNStageIntLLROutputS1xD(138)(3);
  VNStageIntLLRInputS1xD(260)(2) <= CNStageIntLLROutputS1xD(138)(4);
  VNStageIntLLRInputS1xD(357)(2) <= CNStageIntLLROutputS1xD(138)(5);
  VNStageIntLLRInputS1xD(1)(1) <= CNStageIntLLROutputS1xD(139)(0);
  VNStageIntLLRInputS1xD(126)(1) <= CNStageIntLLROutputS1xD(139)(1);
  VNStageIntLLRInputS1xD(154)(1) <= CNStageIntLLROutputS1xD(139)(2);
  VNStageIntLLRInputS1xD(195)(1) <= CNStageIntLLROutputS1xD(139)(3);
  VNStageIntLLRInputS1xD(292)(2) <= CNStageIntLLROutputS1xD(139)(4);
  VNStageIntLLRInputS1xD(373)(1) <= CNStageIntLLROutputS1xD(139)(5);
  VNStageIntLLRInputS1xD(63)(2) <= CNStageIntLLROutputS1xD(140)(0);
  VNStageIntLLRInputS1xD(89)(2) <= CNStageIntLLROutputS1xD(140)(1);
  VNStageIntLLRInputS1xD(130)(2) <= CNStageIntLLROutputS1xD(140)(2);
  VNStageIntLLRInputS1xD(227)(2) <= CNStageIntLLROutputS1xD(140)(3);
  VNStageIntLLRInputS1xD(308)(0) <= CNStageIntLLROutputS1xD(140)(4);
  VNStageIntLLRInputS1xD(343)(2) <= CNStageIntLLROutputS1xD(140)(5);
  VNStageIntLLRInputS1xD(62)(1) <= CNStageIntLLROutputS1xD(141)(0);
  VNStageIntLLRInputS1xD(65)(2) <= CNStageIntLLROutputS1xD(141)(1);
  VNStageIntLLRInputS1xD(162)(2) <= CNStageIntLLROutputS1xD(141)(2);
  VNStageIntLLRInputS1xD(243)(2) <= CNStageIntLLROutputS1xD(141)(3);
  VNStageIntLLRInputS1xD(278)(2) <= CNStageIntLLROutputS1xD(141)(4);
  VNStageIntLLRInputS1xD(352)(2) <= CNStageIntLLROutputS1xD(141)(5);
  VNStageIntLLRInputS1xD(61)(1) <= CNStageIntLLROutputS1xD(142)(0);
  VNStageIntLLRInputS1xD(97)(2) <= CNStageIntLLROutputS1xD(142)(1);
  VNStageIntLLRInputS1xD(178)(2) <= CNStageIntLLROutputS1xD(142)(2);
  VNStageIntLLRInputS1xD(213)(2) <= CNStageIntLLROutputS1xD(142)(3);
  VNStageIntLLRInputS1xD(287)(2) <= CNStageIntLLROutputS1xD(142)(4);
  VNStageIntLLRInputS1xD(365)(2) <= CNStageIntLLROutputS1xD(142)(5);
  VNStageIntLLRInputS1xD(60)(1) <= CNStageIntLLROutputS1xD(143)(0);
  VNStageIntLLRInputS1xD(113)(2) <= CNStageIntLLROutputS1xD(143)(1);
  VNStageIntLLRInputS1xD(148)(2) <= CNStageIntLLROutputS1xD(143)(2);
  VNStageIntLLRInputS1xD(222)(1) <= CNStageIntLLROutputS1xD(143)(3);
  VNStageIntLLRInputS1xD(300)(2) <= CNStageIntLLROutputS1xD(143)(4);
  VNStageIntLLRInputS1xD(344)(2) <= CNStageIntLLROutputS1xD(143)(5);
  VNStageIntLLRInputS1xD(59)(0) <= CNStageIntLLROutputS1xD(144)(0);
  VNStageIntLLRInputS1xD(83)(2) <= CNStageIntLLROutputS1xD(144)(1);
  VNStageIntLLRInputS1xD(157)(2) <= CNStageIntLLROutputS1xD(144)(2);
  VNStageIntLLRInputS1xD(235)(1) <= CNStageIntLLROutputS1xD(144)(3);
  VNStageIntLLRInputS1xD(279)(2) <= CNStageIntLLROutputS1xD(144)(4);
  VNStageIntLLRInputS1xD(372)(1) <= CNStageIntLLROutputS1xD(144)(5);
  VNStageIntLLRInputS1xD(58)(1) <= CNStageIntLLROutputS1xD(145)(0);
  VNStageIntLLRInputS1xD(92)(2) <= CNStageIntLLROutputS1xD(145)(1);
  VNStageIntLLRInputS1xD(170)(2) <= CNStageIntLLROutputS1xD(145)(2);
  VNStageIntLLRInputS1xD(214)(2) <= CNStageIntLLROutputS1xD(145)(3);
  VNStageIntLLRInputS1xD(307)(2) <= CNStageIntLLROutputS1xD(145)(4);
  VNStageIntLLRInputS1xD(374)(2) <= CNStageIntLLROutputS1xD(145)(5);
  VNStageIntLLRInputS1xD(57)(1) <= CNStageIntLLROutputS1xD(146)(0);
  VNStageIntLLRInputS1xD(105)(1) <= CNStageIntLLROutputS1xD(146)(1);
  VNStageIntLLRInputS1xD(149)(2) <= CNStageIntLLROutputS1xD(146)(2);
  VNStageIntLLRInputS1xD(242)(2) <= CNStageIntLLROutputS1xD(146)(3);
  VNStageIntLLRInputS1xD(309)(2) <= CNStageIntLLROutputS1xD(146)(4);
  VNStageIntLLRInputS1xD(356)(2) <= CNStageIntLLROutputS1xD(146)(5);
  VNStageIntLLRInputS1xD(56)(2) <= CNStageIntLLROutputS1xD(147)(0);
  VNStageIntLLRInputS1xD(84)(2) <= CNStageIntLLROutputS1xD(147)(1);
  VNStageIntLLRInputS1xD(177)(2) <= CNStageIntLLROutputS1xD(147)(2);
  VNStageIntLLRInputS1xD(244)(0) <= CNStageIntLLROutputS1xD(147)(3);
  VNStageIntLLRInputS1xD(291)(2) <= CNStageIntLLROutputS1xD(147)(4);
  VNStageIntLLRInputS1xD(363)(1) <= CNStageIntLLROutputS1xD(147)(5);
  VNStageIntLLRInputS1xD(55)(2) <= CNStageIntLLROutputS1xD(148)(0);
  VNStageIntLLRInputS1xD(112)(2) <= CNStageIntLLROutputS1xD(148)(1);
  VNStageIntLLRInputS1xD(179)(2) <= CNStageIntLLROutputS1xD(148)(2);
  VNStageIntLLRInputS1xD(226)(1) <= CNStageIntLLROutputS1xD(148)(3);
  VNStageIntLLRInputS1xD(298)(2) <= CNStageIntLLROutputS1xD(148)(4);
  VNStageIntLLRInputS1xD(327)(2) <= CNStageIntLLROutputS1xD(148)(5);
  VNStageIntLLRInputS1xD(54)(2) <= CNStageIntLLROutputS1xD(149)(0);
  VNStageIntLLRInputS1xD(114)(2) <= CNStageIntLLROutputS1xD(149)(1);
  VNStageIntLLRInputS1xD(161)(2) <= CNStageIntLLROutputS1xD(149)(2);
  VNStageIntLLRInputS1xD(233)(2) <= CNStageIntLLROutputS1xD(149)(3);
  VNStageIntLLRInputS1xD(262)(2) <= CNStageIntLLROutputS1xD(149)(4);
  VNStageIntLLRInputS1xD(378)(1) <= CNStageIntLLROutputS1xD(149)(5);
  VNStageIntLLRInputS1xD(53)(1) <= CNStageIntLLROutputS1xD(150)(0);
  VNStageIntLLRInputS1xD(96)(2) <= CNStageIntLLROutputS1xD(150)(1);
  VNStageIntLLRInputS1xD(168)(1) <= CNStageIntLLROutputS1xD(150)(2);
  VNStageIntLLRInputS1xD(197)(2) <= CNStageIntLLROutputS1xD(150)(3);
  VNStageIntLLRInputS1xD(313)(0) <= CNStageIntLLROutputS1xD(150)(4);
  VNStageIntLLRInputS1xD(321)(2) <= CNStageIntLLROutputS1xD(150)(5);
  VNStageIntLLRInputS1xD(52)(1) <= CNStageIntLLROutputS1xD(151)(0);
  VNStageIntLLRInputS1xD(103)(2) <= CNStageIntLLROutputS1xD(151)(1);
  VNStageIntLLRInputS1xD(132)(1) <= CNStageIntLLROutputS1xD(151)(2);
  VNStageIntLLRInputS1xD(248)(2) <= CNStageIntLLROutputS1xD(151)(3);
  VNStageIntLLRInputS1xD(319)(2) <= CNStageIntLLROutputS1xD(151)(4);
  VNStageIntLLRInputS1xD(379)(1) <= CNStageIntLLROutputS1xD(151)(5);
  VNStageIntLLRInputS1xD(50)(2) <= CNStageIntLLROutputS1xD(152)(0);
  VNStageIntLLRInputS1xD(118)(2) <= CNStageIntLLROutputS1xD(152)(1);
  VNStageIntLLRInputS1xD(189)(1) <= CNStageIntLLROutputS1xD(152)(2);
  VNStageIntLLRInputS1xD(249)(0) <= CNStageIntLLROutputS1xD(152)(3);
  VNStageIntLLRInputS1xD(261)(2) <= CNStageIntLLROutputS1xD(152)(4);
  VNStageIntLLRInputS1xD(348)(2) <= CNStageIntLLROutputS1xD(152)(5);
  VNStageIntLLRInputS1xD(49)(2) <= CNStageIntLLROutputS1xD(153)(0);
  VNStageIntLLRInputS1xD(124)(1) <= CNStageIntLLROutputS1xD(153)(1);
  VNStageIntLLRInputS1xD(184)(2) <= CNStageIntLLROutputS1xD(153)(2);
  VNStageIntLLRInputS1xD(196)(2) <= CNStageIntLLROutputS1xD(153)(3);
  VNStageIntLLRInputS1xD(283)(2) <= CNStageIntLLROutputS1xD(153)(4);
  VNStageIntLLRInputS1xD(366)(2) <= CNStageIntLLROutputS1xD(153)(5);
  VNStageIntLLRInputS1xD(48)(1) <= CNStageIntLLROutputS1xD(154)(0);
  VNStageIntLLRInputS1xD(119)(2) <= CNStageIntLLROutputS1xD(154)(1);
  VNStageIntLLRInputS1xD(131)(1) <= CNStageIntLLROutputS1xD(154)(2);
  VNStageIntLLRInputS1xD(218)(2) <= CNStageIntLLROutputS1xD(154)(3);
  VNStageIntLLRInputS1xD(301)(2) <= CNStageIntLLROutputS1xD(154)(4);
  VNStageIntLLRInputS1xD(351)(1) <= CNStageIntLLROutputS1xD(154)(5);
  VNStageIntLLRInputS1xD(47)(1) <= CNStageIntLLROutputS1xD(155)(0);
  VNStageIntLLRInputS1xD(66)(2) <= CNStageIntLLROutputS1xD(155)(1);
  VNStageIntLLRInputS1xD(153)(2) <= CNStageIntLLROutputS1xD(155)(2);
  VNStageIntLLRInputS1xD(236)(2) <= CNStageIntLLROutputS1xD(155)(3);
  VNStageIntLLRInputS1xD(286)(2) <= CNStageIntLLROutputS1xD(155)(4);
  VNStageIntLLRInputS1xD(338)(2) <= CNStageIntLLROutputS1xD(155)(5);
  VNStageIntLLRInputS1xD(46)(2) <= CNStageIntLLROutputS1xD(156)(0);
  VNStageIntLLRInputS1xD(88)(2) <= CNStageIntLLROutputS1xD(156)(1);
  VNStageIntLLRInputS1xD(171)(1) <= CNStageIntLLROutputS1xD(156)(2);
  VNStageIntLLRInputS1xD(221)(2) <= CNStageIntLLROutputS1xD(156)(3);
  VNStageIntLLRInputS1xD(273)(2) <= CNStageIntLLROutputS1xD(156)(4);
  VNStageIntLLRInputS1xD(369)(1) <= CNStageIntLLROutputS1xD(156)(5);
  VNStageIntLLRInputS1xD(45)(2) <= CNStageIntLLROutputS1xD(157)(0);
  VNStageIntLLRInputS1xD(106)(1) <= CNStageIntLLROutputS1xD(157)(1);
  VNStageIntLLRInputS1xD(156)(2) <= CNStageIntLLROutputS1xD(157)(2);
  VNStageIntLLRInputS1xD(208)(2) <= CNStageIntLLROutputS1xD(157)(3);
  VNStageIntLLRInputS1xD(304)(2) <= CNStageIntLLROutputS1xD(157)(4);
  VNStageIntLLRInputS1xD(381)(1) <= CNStageIntLLROutputS1xD(157)(5);
  VNStageIntLLRInputS1xD(44)(2) <= CNStageIntLLROutputS1xD(158)(0);
  VNStageIntLLRInputS1xD(91)(2) <= CNStageIntLLROutputS1xD(158)(1);
  VNStageIntLLRInputS1xD(143)(2) <= CNStageIntLLROutputS1xD(158)(2);
  VNStageIntLLRInputS1xD(239)(2) <= CNStageIntLLROutputS1xD(158)(3);
  VNStageIntLLRInputS1xD(316)(1) <= CNStageIntLLROutputS1xD(158)(4);
  VNStageIntLLRInputS1xD(332)(2) <= CNStageIntLLROutputS1xD(158)(5);
  VNStageIntLLRInputS1xD(43)(1) <= CNStageIntLLROutputS1xD(159)(0);
  VNStageIntLLRInputS1xD(78)(2) <= CNStageIntLLROutputS1xD(159)(1);
  VNStageIntLLRInputS1xD(174)(2) <= CNStageIntLLROutputS1xD(159)(2);
  VNStageIntLLRInputS1xD(251)(1) <= CNStageIntLLROutputS1xD(159)(3);
  VNStageIntLLRInputS1xD(267)(2) <= CNStageIntLLROutputS1xD(159)(4);
  VNStageIntLLRInputS1xD(376)(2) <= CNStageIntLLROutputS1xD(159)(5);
  VNStageIntLLRInputS1xD(42)(2) <= CNStageIntLLROutputS1xD(160)(0);
  VNStageIntLLRInputS1xD(109)(2) <= CNStageIntLLROutputS1xD(160)(1);
  VNStageIntLLRInputS1xD(186)(1) <= CNStageIntLLROutputS1xD(160)(2);
  VNStageIntLLRInputS1xD(202)(2) <= CNStageIntLLROutputS1xD(160)(3);
  VNStageIntLLRInputS1xD(311)(2) <= CNStageIntLLROutputS1xD(160)(4);
  VNStageIntLLRInputS1xD(353)(2) <= CNStageIntLLROutputS1xD(160)(5);
  VNStageIntLLRInputS1xD(41)(2) <= CNStageIntLLROutputS1xD(161)(0);
  VNStageIntLLRInputS1xD(121)(1) <= CNStageIntLLROutputS1xD(161)(1);
  VNStageIntLLRInputS1xD(137)(2) <= CNStageIntLLROutputS1xD(161)(2);
  VNStageIntLLRInputS1xD(246)(2) <= CNStageIntLLROutputS1xD(161)(3);
  VNStageIntLLRInputS1xD(288)(2) <= CNStageIntLLROutputS1xD(161)(4);
  VNStageIntLLRInputS1xD(342)(2) <= CNStageIntLLROutputS1xD(161)(5);
  VNStageIntLLRInputS1xD(40)(2) <= CNStageIntLLROutputS1xD(162)(0);
  VNStageIntLLRInputS1xD(72)(2) <= CNStageIntLLROutputS1xD(162)(1);
  VNStageIntLLRInputS1xD(181)(2) <= CNStageIntLLROutputS1xD(162)(2);
  VNStageIntLLRInputS1xD(223)(2) <= CNStageIntLLROutputS1xD(162)(3);
  VNStageIntLLRInputS1xD(277)(2) <= CNStageIntLLROutputS1xD(162)(4);
  VNStageIntLLRInputS1xD(346)(2) <= CNStageIntLLROutputS1xD(162)(5);
  VNStageIntLLRInputS1xD(39)(2) <= CNStageIntLLROutputS1xD(163)(0);
  VNStageIntLLRInputS1xD(116)(1) <= CNStageIntLLROutputS1xD(163)(1);
  VNStageIntLLRInputS1xD(158)(2) <= CNStageIntLLROutputS1xD(163)(2);
  VNStageIntLLRInputS1xD(212)(2) <= CNStageIntLLROutputS1xD(163)(3);
  VNStageIntLLRInputS1xD(281)(2) <= CNStageIntLLROutputS1xD(163)(4);
  VNStageIntLLRInputS1xD(339)(2) <= CNStageIntLLROutputS1xD(163)(5);
  VNStageIntLLRInputS1xD(38)(2) <= CNStageIntLLROutputS1xD(164)(0);
  VNStageIntLLRInputS1xD(93)(2) <= CNStageIntLLROutputS1xD(164)(1);
  VNStageIntLLRInputS1xD(147)(2) <= CNStageIntLLROutputS1xD(164)(2);
  VNStageIntLLRInputS1xD(216)(2) <= CNStageIntLLROutputS1xD(164)(3);
  VNStageIntLLRInputS1xD(274)(1) <= CNStageIntLLROutputS1xD(164)(4);
  VNStageIntLLRInputS1xD(350)(2) <= CNStageIntLLROutputS1xD(164)(5);
  VNStageIntLLRInputS1xD(37)(2) <= CNStageIntLLROutputS1xD(165)(0);
  VNStageIntLLRInputS1xD(82)(2) <= CNStageIntLLROutputS1xD(165)(1);
  VNStageIntLLRInputS1xD(151)(2) <= CNStageIntLLROutputS1xD(165)(2);
  VNStageIntLLRInputS1xD(209)(2) <= CNStageIntLLROutputS1xD(165)(3);
  VNStageIntLLRInputS1xD(285)(2) <= CNStageIntLLROutputS1xD(165)(4);
  VNStageIntLLRInputS1xD(322)(2) <= CNStageIntLLROutputS1xD(165)(5);
  VNStageIntLLRInputS1xD(36)(2) <= CNStageIntLLROutputS1xD(166)(0);
  VNStageIntLLRInputS1xD(86)(1) <= CNStageIntLLROutputS1xD(166)(1);
  VNStageIntLLRInputS1xD(144)(2) <= CNStageIntLLROutputS1xD(166)(2);
  VNStageIntLLRInputS1xD(220)(2) <= CNStageIntLLROutputS1xD(166)(3);
  VNStageIntLLRInputS1xD(257)(2) <= CNStageIntLLROutputS1xD(166)(4);
  VNStageIntLLRInputS1xD(377)(1) <= CNStageIntLLROutputS1xD(166)(5);
  VNStageIntLLRInputS1xD(35)(2) <= CNStageIntLLROutputS1xD(167)(0);
  VNStageIntLLRInputS1xD(79)(2) <= CNStageIntLLROutputS1xD(167)(1);
  VNStageIntLLRInputS1xD(155)(2) <= CNStageIntLLROutputS1xD(167)(2);
  VNStageIntLLRInputS1xD(255)(2) <= CNStageIntLLROutputS1xD(167)(3);
  VNStageIntLLRInputS1xD(312)(2) <= CNStageIntLLROutputS1xD(167)(4);
  VNStageIntLLRInputS1xD(331)(2) <= CNStageIntLLROutputS1xD(167)(5);
  VNStageIntLLRInputS1xD(34)(2) <= CNStageIntLLROutputS1xD(168)(0);
  VNStageIntLLRInputS1xD(90)(2) <= CNStageIntLLROutputS1xD(168)(1);
  VNStageIntLLRInputS1xD(190)(0) <= CNStageIntLLROutputS1xD(168)(2);
  VNStageIntLLRInputS1xD(247)(2) <= CNStageIntLLROutputS1xD(168)(3);
  VNStageIntLLRInputS1xD(266)(1) <= CNStageIntLLROutputS1xD(168)(4);
  VNStageIntLLRInputS1xD(328)(2) <= CNStageIntLLROutputS1xD(168)(5);
  VNStageIntLLRInputS1xD(33)(2) <= CNStageIntLLROutputS1xD(169)(0);
  VNStageIntLLRInputS1xD(125)(1) <= CNStageIntLLROutputS1xD(169)(1);
  VNStageIntLLRInputS1xD(182)(2) <= CNStageIntLLROutputS1xD(169)(2);
  VNStageIntLLRInputS1xD(201)(2) <= CNStageIntLLROutputS1xD(169)(3);
  VNStageIntLLRInputS1xD(263)(2) <= CNStageIntLLROutputS1xD(169)(4);
  VNStageIntLLRInputS1xD(362)(2) <= CNStageIntLLROutputS1xD(169)(5);
  VNStageIntLLRInputS1xD(0)(2) <= CNStageIntLLROutputS1xD(170)(0);
  VNStageIntLLRInputS1xD(75)(2) <= CNStageIntLLROutputS1xD(170)(1);
  VNStageIntLLRInputS1xD(140)(2) <= CNStageIntLLROutputS1xD(170)(2);
  VNStageIntLLRInputS1xD(205)(0) <= CNStageIntLLROutputS1xD(170)(3);
  VNStageIntLLRInputS1xD(270)(2) <= CNStageIntLLROutputS1xD(170)(4);
  VNStageIntLLRInputS1xD(335)(2) <= CNStageIntLLROutputS1xD(170)(5);
  VNStageIntLLRInputS1xD(62)(2) <= CNStageIntLLROutputS1xD(171)(0);
  VNStageIntLLRInputS1xD(109)(3) <= CNStageIntLLROutputS1xD(171)(1);
  VNStageIntLLRInputS1xD(161)(3) <= CNStageIntLLROutputS1xD(171)(2);
  VNStageIntLLRInputS1xD(194)(3) <= CNStageIntLLROutputS1xD(171)(3);
  VNStageIntLLRInputS1xD(271)(2) <= CNStageIntLLROutputS1xD(171)(4);
  VNStageIntLLRInputS1xD(350)(3) <= CNStageIntLLROutputS1xD(171)(5);
  VNStageIntLLRInputS1xD(61)(2) <= CNStageIntLLROutputS1xD(172)(0);
  VNStageIntLLRInputS1xD(96)(3) <= CNStageIntLLROutputS1xD(172)(1);
  VNStageIntLLRInputS1xD(129)(3) <= CNStageIntLLROutputS1xD(172)(2);
  VNStageIntLLRInputS1xD(206)(2) <= CNStageIntLLROutputS1xD(172)(3);
  VNStageIntLLRInputS1xD(285)(3) <= CNStageIntLLROutputS1xD(172)(4);
  VNStageIntLLRInputS1xD(331)(3) <= CNStageIntLLROutputS1xD(172)(5);
  VNStageIntLLRInputS1xD(60)(2) <= CNStageIntLLROutputS1xD(173)(0);
  VNStageIntLLRInputS1xD(127)(3) <= CNStageIntLLROutputS1xD(173)(1);
  VNStageIntLLRInputS1xD(141)(1) <= CNStageIntLLROutputS1xD(173)(2);
  VNStageIntLLRInputS1xD(220)(3) <= CNStageIntLLROutputS1xD(173)(3);
  VNStageIntLLRInputS1xD(266)(2) <= CNStageIntLLROutputS1xD(173)(4);
  VNStageIntLLRInputS1xD(371)(2) <= CNStageIntLLROutputS1xD(173)(5);
  VNStageIntLLRInputS1xD(59)(1) <= CNStageIntLLROutputS1xD(174)(0);
  VNStageIntLLRInputS1xD(76)(3) <= CNStageIntLLROutputS1xD(174)(1);
  VNStageIntLLRInputS1xD(155)(3) <= CNStageIntLLROutputS1xD(174)(2);
  VNStageIntLLRInputS1xD(201)(3) <= CNStageIntLLROutputS1xD(174)(3);
  VNStageIntLLRInputS1xD(306)(3) <= CNStageIntLLROutputS1xD(174)(4);
  VNStageIntLLRInputS1xD(360)(3) <= CNStageIntLLROutputS1xD(174)(5);
  VNStageIntLLRInputS1xD(58)(2) <= CNStageIntLLROutputS1xD(175)(0);
  VNStageIntLLRInputS1xD(90)(3) <= CNStageIntLLROutputS1xD(175)(1);
  VNStageIntLLRInputS1xD(136)(3) <= CNStageIntLLROutputS1xD(175)(2);
  VNStageIntLLRInputS1xD(241)(2) <= CNStageIntLLROutputS1xD(175)(3);
  VNStageIntLLRInputS1xD(295)(3) <= CNStageIntLLROutputS1xD(175)(4);
  VNStageIntLLRInputS1xD(364)(3) <= CNStageIntLLROutputS1xD(175)(5);
  VNStageIntLLRInputS1xD(57)(2) <= CNStageIntLLROutputS1xD(176)(0);
  VNStageIntLLRInputS1xD(71)(2) <= CNStageIntLLROutputS1xD(176)(1);
  VNStageIntLLRInputS1xD(176)(3) <= CNStageIntLLROutputS1xD(176)(2);
  VNStageIntLLRInputS1xD(230)(2) <= CNStageIntLLROutputS1xD(176)(3);
  VNStageIntLLRInputS1xD(299)(2) <= CNStageIntLLROutputS1xD(176)(4);
  VNStageIntLLRInputS1xD(357)(3) <= CNStageIntLLROutputS1xD(176)(5);
  VNStageIntLLRInputS1xD(56)(3) <= CNStageIntLLROutputS1xD(177)(0);
  VNStageIntLLRInputS1xD(111)(3) <= CNStageIntLLROutputS1xD(177)(1);
  VNStageIntLLRInputS1xD(165)(3) <= CNStageIntLLROutputS1xD(177)(2);
  VNStageIntLLRInputS1xD(234)(3) <= CNStageIntLLROutputS1xD(177)(3);
  VNStageIntLLRInputS1xD(292)(3) <= CNStageIntLLROutputS1xD(177)(4);
  VNStageIntLLRInputS1xD(368)(1) <= CNStageIntLLROutputS1xD(177)(5);
  VNStageIntLLRInputS1xD(55)(3) <= CNStageIntLLROutputS1xD(178)(0);
  VNStageIntLLRInputS1xD(100)(3) <= CNStageIntLLROutputS1xD(178)(1);
  VNStageIntLLRInputS1xD(169)(3) <= CNStageIntLLROutputS1xD(178)(2);
  VNStageIntLLRInputS1xD(227)(3) <= CNStageIntLLROutputS1xD(178)(3);
  VNStageIntLLRInputS1xD(303)(3) <= CNStageIntLLROutputS1xD(178)(4);
  VNStageIntLLRInputS1xD(340)(3) <= CNStageIntLLROutputS1xD(178)(5);
  VNStageIntLLRInputS1xD(54)(3) <= CNStageIntLLROutputS1xD(179)(0);
  VNStageIntLLRInputS1xD(104)(3) <= CNStageIntLLROutputS1xD(179)(1);
  VNStageIntLLRInputS1xD(162)(3) <= CNStageIntLLROutputS1xD(179)(2);
  VNStageIntLLRInputS1xD(238)(3) <= CNStageIntLLROutputS1xD(179)(3);
  VNStageIntLLRInputS1xD(275)(3) <= CNStageIntLLROutputS1xD(179)(4);
  VNStageIntLLRInputS1xD(332)(3) <= CNStageIntLLROutputS1xD(179)(5);
  VNStageIntLLRInputS1xD(53)(2) <= CNStageIntLLROutputS1xD(180)(0);
  VNStageIntLLRInputS1xD(97)(3) <= CNStageIntLLROutputS1xD(180)(1);
  VNStageIntLLRInputS1xD(173)(3) <= CNStageIntLLROutputS1xD(180)(2);
  VNStageIntLLRInputS1xD(210)(3) <= CNStageIntLLROutputS1xD(180)(3);
  VNStageIntLLRInputS1xD(267)(3) <= CNStageIntLLROutputS1xD(180)(4);
  VNStageIntLLRInputS1xD(349)(2) <= CNStageIntLLROutputS1xD(180)(5);
  VNStageIntLLRInputS1xD(52)(2) <= CNStageIntLLROutputS1xD(181)(0);
  VNStageIntLLRInputS1xD(108)(3) <= CNStageIntLLROutputS1xD(181)(1);
  VNStageIntLLRInputS1xD(145)(3) <= CNStageIntLLROutputS1xD(181)(2);
  VNStageIntLLRInputS1xD(202)(3) <= CNStageIntLLROutputS1xD(181)(3);
  VNStageIntLLRInputS1xD(284)(3) <= CNStageIntLLROutputS1xD(181)(4);
  VNStageIntLLRInputS1xD(346)(3) <= CNStageIntLLROutputS1xD(181)(5);
  VNStageIntLLRInputS1xD(51)(2) <= CNStageIntLLROutputS1xD(182)(0);
  VNStageIntLLRInputS1xD(80)(3) <= CNStageIntLLROutputS1xD(182)(1);
  VNStageIntLLRInputS1xD(137)(3) <= CNStageIntLLROutputS1xD(182)(2);
  VNStageIntLLRInputS1xD(219)(3) <= CNStageIntLLROutputS1xD(182)(3);
  VNStageIntLLRInputS1xD(281)(3) <= CNStageIntLLROutputS1xD(182)(4);
  VNStageIntLLRInputS1xD(380)(2) <= CNStageIntLLROutputS1xD(182)(5);
  VNStageIntLLRInputS1xD(50)(3) <= CNStageIntLLROutputS1xD(183)(0);
  VNStageIntLLRInputS1xD(72)(3) <= CNStageIntLLROutputS1xD(183)(1);
  VNStageIntLLRInputS1xD(154)(2) <= CNStageIntLLROutputS1xD(183)(2);
  VNStageIntLLRInputS1xD(216)(3) <= CNStageIntLLROutputS1xD(183)(3);
  VNStageIntLLRInputS1xD(315)(2) <= CNStageIntLLROutputS1xD(183)(4);
  VNStageIntLLRInputS1xD(337)(3) <= CNStageIntLLROutputS1xD(183)(5);
  VNStageIntLLRInputS1xD(49)(3) <= CNStageIntLLROutputS1xD(184)(0);
  VNStageIntLLRInputS1xD(89)(3) <= CNStageIntLLROutputS1xD(184)(1);
  VNStageIntLLRInputS1xD(151)(3) <= CNStageIntLLROutputS1xD(184)(2);
  VNStageIntLLRInputS1xD(250)(2) <= CNStageIntLLROutputS1xD(184)(3);
  VNStageIntLLRInputS1xD(272)(3) <= CNStageIntLLROutputS1xD(184)(4);
  VNStageIntLLRInputS1xD(323)(2) <= CNStageIntLLROutputS1xD(184)(5);
  VNStageIntLLRInputS1xD(46)(3) <= CNStageIntLLROutputS1xD(185)(0);
  VNStageIntLLRInputS1xD(77)(1) <= CNStageIntLLROutputS1xD(185)(1);
  VNStageIntLLRInputS1xD(191)(3) <= CNStageIntLLROutputS1xD(185)(2);
  VNStageIntLLRInputS1xD(246)(3) <= CNStageIntLLROutputS1xD(185)(3);
  VNStageIntLLRInputS1xD(277)(3) <= CNStageIntLLROutputS1xD(185)(4);
  VNStageIntLLRInputS1xD(325)(3) <= CNStageIntLLROutputS1xD(185)(5);
  VNStageIntLLRInputS1xD(45)(3) <= CNStageIntLLROutputS1xD(186)(0);
  VNStageIntLLRInputS1xD(126)(2) <= CNStageIntLLROutputS1xD(186)(1);
  VNStageIntLLRInputS1xD(181)(3) <= CNStageIntLLROutputS1xD(186)(2);
  VNStageIntLLRInputS1xD(212)(3) <= CNStageIntLLROutputS1xD(186)(3);
  VNStageIntLLRInputS1xD(260)(3) <= CNStageIntLLROutputS1xD(186)(4);
  VNStageIntLLRInputS1xD(355)(3) <= CNStageIntLLROutputS1xD(186)(5);
  VNStageIntLLRInputS1xD(44)(3) <= CNStageIntLLROutputS1xD(187)(0);
  VNStageIntLLRInputS1xD(116)(2) <= CNStageIntLLROutputS1xD(187)(1);
  VNStageIntLLRInputS1xD(147)(3) <= CNStageIntLLROutputS1xD(187)(2);
  VNStageIntLLRInputS1xD(195)(2) <= CNStageIntLLROutputS1xD(187)(3);
  VNStageIntLLRInputS1xD(290)(3) <= CNStageIntLLROutputS1xD(187)(4);
  VNStageIntLLRInputS1xD(378)(2) <= CNStageIntLLROutputS1xD(187)(5);
  VNStageIntLLRInputS1xD(43)(2) <= CNStageIntLLROutputS1xD(188)(0);
  VNStageIntLLRInputS1xD(82)(3) <= CNStageIntLLROutputS1xD(188)(1);
  VNStageIntLLRInputS1xD(130)(3) <= CNStageIntLLROutputS1xD(188)(2);
  VNStageIntLLRInputS1xD(225)(3) <= CNStageIntLLROutputS1xD(188)(3);
  VNStageIntLLRInputS1xD(313)(1) <= CNStageIntLLROutputS1xD(188)(4);
  VNStageIntLLRInputS1xD(351)(2) <= CNStageIntLLROutputS1xD(188)(5);
  VNStageIntLLRInputS1xD(42)(3) <= CNStageIntLLROutputS1xD(189)(0);
  VNStageIntLLRInputS1xD(65)(3) <= CNStageIntLLROutputS1xD(189)(1);
  VNStageIntLLRInputS1xD(160)(3) <= CNStageIntLLROutputS1xD(189)(2);
  VNStageIntLLRInputS1xD(248)(3) <= CNStageIntLLROutputS1xD(189)(3);
  VNStageIntLLRInputS1xD(286)(3) <= CNStageIntLLROutputS1xD(189)(4);
  VNStageIntLLRInputS1xD(335)(3) <= CNStageIntLLROutputS1xD(189)(5);
  VNStageIntLLRInputS1xD(41)(3) <= CNStageIntLLROutputS1xD(190)(0);
  VNStageIntLLRInputS1xD(95)(3) <= CNStageIntLLROutputS1xD(190)(1);
  VNStageIntLLRInputS1xD(183)(2) <= CNStageIntLLROutputS1xD(190)(2);
  VNStageIntLLRInputS1xD(221)(3) <= CNStageIntLLROutputS1xD(190)(3);
  VNStageIntLLRInputS1xD(270)(3) <= CNStageIntLLROutputS1xD(190)(4);
  VNStageIntLLRInputS1xD(338)(3) <= CNStageIntLLROutputS1xD(190)(5);
  VNStageIntLLRInputS1xD(39)(3) <= CNStageIntLLROutputS1xD(191)(0);
  VNStageIntLLRInputS1xD(91)(3) <= CNStageIntLLROutputS1xD(191)(1);
  VNStageIntLLRInputS1xD(140)(3) <= CNStageIntLLROutputS1xD(191)(2);
  VNStageIntLLRInputS1xD(208)(3) <= CNStageIntLLROutputS1xD(191)(3);
  VNStageIntLLRInputS1xD(314)(0) <= CNStageIntLLROutputS1xD(191)(4);
  VNStageIntLLRInputS1xD(354)(3) <= CNStageIntLLROutputS1xD(191)(5);
  VNStageIntLLRInputS1xD(38)(3) <= CNStageIntLLROutputS1xD(192)(0);
  VNStageIntLLRInputS1xD(75)(3) <= CNStageIntLLROutputS1xD(192)(1);
  VNStageIntLLRInputS1xD(143)(3) <= CNStageIntLLROutputS1xD(192)(2);
  VNStageIntLLRInputS1xD(249)(1) <= CNStageIntLLROutputS1xD(192)(3);
  VNStageIntLLRInputS1xD(289)(3) <= CNStageIntLLROutputS1xD(192)(4);
  VNStageIntLLRInputS1xD(352)(3) <= CNStageIntLLROutputS1xD(192)(5);
  VNStageIntLLRInputS1xD(37)(3) <= CNStageIntLLROutputS1xD(193)(0);
  VNStageIntLLRInputS1xD(78)(3) <= CNStageIntLLROutputS1xD(193)(1);
  VNStageIntLLRInputS1xD(184)(3) <= CNStageIntLLROutputS1xD(193)(2);
  VNStageIntLLRInputS1xD(224)(3) <= CNStageIntLLROutputS1xD(193)(3);
  VNStageIntLLRInputS1xD(287)(3) <= CNStageIntLLROutputS1xD(193)(4);
  VNStageIntLLRInputS1xD(377)(2) <= CNStageIntLLROutputS1xD(193)(5);
  VNStageIntLLRInputS1xD(35)(3) <= CNStageIntLLROutputS1xD(194)(0);
  VNStageIntLLRInputS1xD(94)(2) <= CNStageIntLLROutputS1xD(194)(1);
  VNStageIntLLRInputS1xD(157)(3) <= CNStageIntLLROutputS1xD(194)(2);
  VNStageIntLLRInputS1xD(247)(3) <= CNStageIntLLROutputS1xD(194)(3);
  VNStageIntLLRInputS1xD(257)(3) <= CNStageIntLLROutputS1xD(194)(4);
  VNStageIntLLRInputS1xD(365)(3) <= CNStageIntLLROutputS1xD(194)(5);
  VNStageIntLLRInputS1xD(34)(3) <= CNStageIntLLROutputS1xD(195)(0);
  VNStageIntLLRInputS1xD(92)(3) <= CNStageIntLLROutputS1xD(195)(1);
  VNStageIntLLRInputS1xD(182)(3) <= CNStageIntLLROutputS1xD(195)(2);
  VNStageIntLLRInputS1xD(255)(3) <= CNStageIntLLROutputS1xD(195)(3);
  VNStageIntLLRInputS1xD(300)(3) <= CNStageIntLLROutputS1xD(195)(4);
  VNStageIntLLRInputS1xD(359)(3) <= CNStageIntLLROutputS1xD(195)(5);
  VNStageIntLLRInputS1xD(33)(3) <= CNStageIntLLROutputS1xD(196)(0);
  VNStageIntLLRInputS1xD(117)(3) <= CNStageIntLLROutputS1xD(196)(1);
  VNStageIntLLRInputS1xD(190)(1) <= CNStageIntLLROutputS1xD(196)(2);
  VNStageIntLLRInputS1xD(235)(2) <= CNStageIntLLROutputS1xD(196)(3);
  VNStageIntLLRInputS1xD(294)(3) <= CNStageIntLLROutputS1xD(196)(4);
  VNStageIntLLRInputS1xD(320)(2) <= CNStageIntLLROutputS1xD(196)(5);
  VNStageIntLLRInputS1xD(31)(2) <= CNStageIntLLROutputS1xD(197)(0);
  VNStageIntLLRInputS1xD(105)(2) <= CNStageIntLLROutputS1xD(197)(1);
  VNStageIntLLRInputS1xD(164)(3) <= CNStageIntLLROutputS1xD(197)(2);
  VNStageIntLLRInputS1xD(192)(3) <= CNStageIntLLROutputS1xD(197)(3);
  VNStageIntLLRInputS1xD(293)(3) <= CNStageIntLLROutputS1xD(197)(4);
  VNStageIntLLRInputS1xD(363)(2) <= CNStageIntLLROutputS1xD(197)(5);
  VNStageIntLLRInputS1xD(30)(3) <= CNStageIntLLROutputS1xD(198)(0);
  VNStageIntLLRInputS1xD(99)(3) <= CNStageIntLLROutputS1xD(198)(1);
  VNStageIntLLRInputS1xD(128)(3) <= CNStageIntLLROutputS1xD(198)(2);
  VNStageIntLLRInputS1xD(228)(3) <= CNStageIntLLROutputS1xD(198)(3);
  VNStageIntLLRInputS1xD(298)(3) <= CNStageIntLLROutputS1xD(198)(4);
  VNStageIntLLRInputS1xD(382)(2) <= CNStageIntLLROutputS1xD(198)(5);
  VNStageIntLLRInputS1xD(28)(3) <= CNStageIntLLROutputS1xD(199)(0);
  VNStageIntLLRInputS1xD(98)(2) <= CNStageIntLLROutputS1xD(199)(1);
  VNStageIntLLRInputS1xD(168)(2) <= CNStageIntLLROutputS1xD(199)(2);
  VNStageIntLLRInputS1xD(252)(2) <= CNStageIntLLROutputS1xD(199)(3);
  VNStageIntLLRInputS1xD(308)(1) <= CNStageIntLLROutputS1xD(199)(4);
  VNStageIntLLRInputS1xD(347)(3) <= CNStageIntLLROutputS1xD(199)(5);
  VNStageIntLLRInputS1xD(27)(3) <= CNStageIntLLROutputS1xD(200)(0);
  VNStageIntLLRInputS1xD(103)(3) <= CNStageIntLLROutputS1xD(200)(1);
  VNStageIntLLRInputS1xD(187)(2) <= CNStageIntLLROutputS1xD(200)(2);
  VNStageIntLLRInputS1xD(243)(3) <= CNStageIntLLROutputS1xD(200)(3);
  VNStageIntLLRInputS1xD(282)(3) <= CNStageIntLLROutputS1xD(200)(4);
  VNStageIntLLRInputS1xD(348)(3) <= CNStageIntLLROutputS1xD(200)(5);
  VNStageIntLLRInputS1xD(26)(3) <= CNStageIntLLROutputS1xD(201)(0);
  VNStageIntLLRInputS1xD(122)(2) <= CNStageIntLLROutputS1xD(201)(1);
  VNStageIntLLRInputS1xD(178)(3) <= CNStageIntLLROutputS1xD(201)(2);
  VNStageIntLLRInputS1xD(217)(3) <= CNStageIntLLROutputS1xD(201)(3);
  VNStageIntLLRInputS1xD(283)(3) <= CNStageIntLLROutputS1xD(201)(4);
  VNStageIntLLRInputS1xD(372)(2) <= CNStageIntLLROutputS1xD(201)(5);
  VNStageIntLLRInputS1xD(25)(3) <= CNStageIntLLROutputS1xD(202)(0);
  VNStageIntLLRInputS1xD(113)(3) <= CNStageIntLLROutputS1xD(202)(1);
  VNStageIntLLRInputS1xD(152)(3) <= CNStageIntLLROutputS1xD(202)(2);
  VNStageIntLLRInputS1xD(218)(3) <= CNStageIntLLROutputS1xD(202)(3);
  VNStageIntLLRInputS1xD(307)(3) <= CNStageIntLLROutputS1xD(202)(4);
  VNStageIntLLRInputS1xD(330)(3) <= CNStageIntLLROutputS1xD(202)(5);
  VNStageIntLLRInputS1xD(24)(3) <= CNStageIntLLROutputS1xD(203)(0);
  VNStageIntLLRInputS1xD(87)(3) <= CNStageIntLLROutputS1xD(203)(1);
  VNStageIntLLRInputS1xD(153)(3) <= CNStageIntLLROutputS1xD(203)(2);
  VNStageIntLLRInputS1xD(242)(3) <= CNStageIntLLROutputS1xD(203)(3);
  VNStageIntLLRInputS1xD(265)(2) <= CNStageIntLLROutputS1xD(203)(4);
  VNStageIntLLRInputS1xD(326)(2) <= CNStageIntLLROutputS1xD(203)(5);
  VNStageIntLLRInputS1xD(23)(3) <= CNStageIntLLROutputS1xD(204)(0);
  VNStageIntLLRInputS1xD(88)(3) <= CNStageIntLLROutputS1xD(204)(1);
  VNStageIntLLRInputS1xD(177)(3) <= CNStageIntLLROutputS1xD(204)(2);
  VNStageIntLLRInputS1xD(200)(3) <= CNStageIntLLROutputS1xD(204)(3);
  VNStageIntLLRInputS1xD(261)(3) <= CNStageIntLLROutputS1xD(204)(4);
  VNStageIntLLRInputS1xD(341)(3) <= CNStageIntLLROutputS1xD(204)(5);
  VNStageIntLLRInputS1xD(22)(3) <= CNStageIntLLROutputS1xD(205)(0);
  VNStageIntLLRInputS1xD(112)(3) <= CNStageIntLLROutputS1xD(205)(1);
  VNStageIntLLRInputS1xD(135)(3) <= CNStageIntLLROutputS1xD(205)(2);
  VNStageIntLLRInputS1xD(196)(3) <= CNStageIntLLROutputS1xD(205)(3);
  VNStageIntLLRInputS1xD(276)(3) <= CNStageIntLLROutputS1xD(205)(4);
  VNStageIntLLRInputS1xD(367)(3) <= CNStageIntLLROutputS1xD(205)(5);
  VNStageIntLLRInputS1xD(21)(3) <= CNStageIntLLROutputS1xD(206)(0);
  VNStageIntLLRInputS1xD(70)(3) <= CNStageIntLLROutputS1xD(206)(1);
  VNStageIntLLRInputS1xD(131)(2) <= CNStageIntLLROutputS1xD(206)(2);
  VNStageIntLLRInputS1xD(211)(3) <= CNStageIntLLROutputS1xD(206)(3);
  VNStageIntLLRInputS1xD(302)(3) <= CNStageIntLLROutputS1xD(206)(4);
  VNStageIntLLRInputS1xD(343)(3) <= CNStageIntLLROutputS1xD(206)(5);
  VNStageIntLLRInputS1xD(18)(3) <= CNStageIntLLROutputS1xD(207)(0);
  VNStageIntLLRInputS1xD(107)(2) <= CNStageIntLLROutputS1xD(207)(1);
  VNStageIntLLRInputS1xD(148)(3) <= CNStageIntLLROutputS1xD(207)(2);
  VNStageIntLLRInputS1xD(245)(3) <= CNStageIntLLROutputS1xD(207)(3);
  VNStageIntLLRInputS1xD(263)(3) <= CNStageIntLLROutputS1xD(207)(4);
  VNStageIntLLRInputS1xD(361)(3) <= CNStageIntLLROutputS1xD(207)(5);
  VNStageIntLLRInputS1xD(17)(3) <= CNStageIntLLROutputS1xD(208)(0);
  VNStageIntLLRInputS1xD(83)(3) <= CNStageIntLLROutputS1xD(208)(1);
  VNStageIntLLRInputS1xD(180)(1) <= CNStageIntLLROutputS1xD(208)(2);
  VNStageIntLLRInputS1xD(198)(3) <= CNStageIntLLROutputS1xD(208)(3);
  VNStageIntLLRInputS1xD(296)(3) <= CNStageIntLLROutputS1xD(208)(4);
  VNStageIntLLRInputS1xD(370)(2) <= CNStageIntLLROutputS1xD(208)(5);
  VNStageIntLLRInputS1xD(16)(2) <= CNStageIntLLROutputS1xD(209)(0);
  VNStageIntLLRInputS1xD(115)(3) <= CNStageIntLLROutputS1xD(209)(1);
  VNStageIntLLRInputS1xD(133)(1) <= CNStageIntLLROutputS1xD(209)(2);
  VNStageIntLLRInputS1xD(231)(2) <= CNStageIntLLROutputS1xD(209)(3);
  VNStageIntLLRInputS1xD(305)(3) <= CNStageIntLLROutputS1xD(209)(4);
  VNStageIntLLRInputS1xD(383)(3) <= CNStageIntLLROutputS1xD(209)(5);
  VNStageIntLLRInputS1xD(15)(3) <= CNStageIntLLROutputS1xD(210)(0);
  VNStageIntLLRInputS1xD(68)(2) <= CNStageIntLLROutputS1xD(210)(1);
  VNStageIntLLRInputS1xD(166)(3) <= CNStageIntLLROutputS1xD(210)(2);
  VNStageIntLLRInputS1xD(240)(3) <= CNStageIntLLROutputS1xD(210)(3);
  VNStageIntLLRInputS1xD(318)(1) <= CNStageIntLLROutputS1xD(210)(4);
  VNStageIntLLRInputS1xD(362)(3) <= CNStageIntLLROutputS1xD(210)(5);
  VNStageIntLLRInputS1xD(14)(3) <= CNStageIntLLROutputS1xD(211)(0);
  VNStageIntLLRInputS1xD(101)(3) <= CNStageIntLLROutputS1xD(211)(1);
  VNStageIntLLRInputS1xD(175)(3) <= CNStageIntLLROutputS1xD(211)(2);
  VNStageIntLLRInputS1xD(253)(2) <= CNStageIntLLROutputS1xD(211)(3);
  VNStageIntLLRInputS1xD(297)(3) <= CNStageIntLLROutputS1xD(211)(4);
  VNStageIntLLRInputS1xD(327)(3) <= CNStageIntLLROutputS1xD(211)(5);
  VNStageIntLLRInputS1xD(13)(2) <= CNStageIntLLROutputS1xD(212)(0);
  VNStageIntLLRInputS1xD(110)(3) <= CNStageIntLLROutputS1xD(212)(1);
  VNStageIntLLRInputS1xD(188)(1) <= CNStageIntLLROutputS1xD(212)(2);
  VNStageIntLLRInputS1xD(232)(2) <= CNStageIntLLROutputS1xD(212)(3);
  VNStageIntLLRInputS1xD(262)(3) <= CNStageIntLLROutputS1xD(212)(4);
  VNStageIntLLRInputS1xD(329)(3) <= CNStageIntLLROutputS1xD(212)(5);
  VNStageIntLLRInputS1xD(12)(3) <= CNStageIntLLROutputS1xD(213)(0);
  VNStageIntLLRInputS1xD(123)(2) <= CNStageIntLLROutputS1xD(213)(1);
  VNStageIntLLRInputS1xD(167)(3) <= CNStageIntLLROutputS1xD(213)(2);
  VNStageIntLLRInputS1xD(197)(3) <= CNStageIntLLROutputS1xD(213)(3);
  VNStageIntLLRInputS1xD(264)(3) <= CNStageIntLLROutputS1xD(213)(4);
  VNStageIntLLRInputS1xD(374)(3) <= CNStageIntLLROutputS1xD(213)(5);
  VNStageIntLLRInputS1xD(11)(3) <= CNStageIntLLROutputS1xD(214)(0);
  VNStageIntLLRInputS1xD(102)(3) <= CNStageIntLLROutputS1xD(214)(1);
  VNStageIntLLRInputS1xD(132)(2) <= CNStageIntLLROutputS1xD(214)(2);
  VNStageIntLLRInputS1xD(199)(3) <= CNStageIntLLROutputS1xD(214)(3);
  VNStageIntLLRInputS1xD(309)(3) <= CNStageIntLLROutputS1xD(214)(4);
  VNStageIntLLRInputS1xD(381)(2) <= CNStageIntLLROutputS1xD(214)(5);
  VNStageIntLLRInputS1xD(9)(3) <= CNStageIntLLROutputS1xD(215)(0);
  VNStageIntLLRInputS1xD(69)(3) <= CNStageIntLLROutputS1xD(215)(1);
  VNStageIntLLRInputS1xD(179)(3) <= CNStageIntLLROutputS1xD(215)(2);
  VNStageIntLLRInputS1xD(251)(2) <= CNStageIntLLROutputS1xD(215)(3);
  VNStageIntLLRInputS1xD(280)(3) <= CNStageIntLLROutputS1xD(215)(4);
  VNStageIntLLRInputS1xD(333)(2) <= CNStageIntLLROutputS1xD(215)(5);
  VNStageIntLLRInputS1xD(8)(2) <= CNStageIntLLROutputS1xD(216)(0);
  VNStageIntLLRInputS1xD(114)(3) <= CNStageIntLLROutputS1xD(216)(1);
  VNStageIntLLRInputS1xD(186)(2) <= CNStageIntLLROutputS1xD(216)(2);
  VNStageIntLLRInputS1xD(215)(3) <= CNStageIntLLROutputS1xD(216)(3);
  VNStageIntLLRInputS1xD(268)(3) <= CNStageIntLLROutputS1xD(216)(4);
  VNStageIntLLRInputS1xD(339)(3) <= CNStageIntLLROutputS1xD(216)(5);
  VNStageIntLLRInputS1xD(7)(3) <= CNStageIntLLROutputS1xD(217)(0);
  VNStageIntLLRInputS1xD(121)(2) <= CNStageIntLLROutputS1xD(217)(1);
  VNStageIntLLRInputS1xD(150)(3) <= CNStageIntLLROutputS1xD(217)(2);
  VNStageIntLLRInputS1xD(203)(3) <= CNStageIntLLROutputS1xD(217)(3);
  VNStageIntLLRInputS1xD(274)(2) <= CNStageIntLLROutputS1xD(217)(4);
  VNStageIntLLRInputS1xD(334)(2) <= CNStageIntLLROutputS1xD(217)(5);
  VNStageIntLLRInputS1xD(6)(3) <= CNStageIntLLROutputS1xD(218)(0);
  VNStageIntLLRInputS1xD(85)(2) <= CNStageIntLLROutputS1xD(218)(1);
  VNStageIntLLRInputS1xD(138)(3) <= CNStageIntLLROutputS1xD(218)(2);
  VNStageIntLLRInputS1xD(209)(3) <= CNStageIntLLROutputS1xD(218)(3);
  VNStageIntLLRInputS1xD(269)(2) <= CNStageIntLLROutputS1xD(218)(4);
  VNStageIntLLRInputS1xD(344)(3) <= CNStageIntLLROutputS1xD(218)(5);
  VNStageIntLLRInputS1xD(5)(3) <= CNStageIntLLROutputS1xD(219)(0);
  VNStageIntLLRInputS1xD(73)(3) <= CNStageIntLLROutputS1xD(219)(1);
  VNStageIntLLRInputS1xD(144)(3) <= CNStageIntLLROutputS1xD(219)(2);
  VNStageIntLLRInputS1xD(204)(3) <= CNStageIntLLROutputS1xD(219)(3);
  VNStageIntLLRInputS1xD(279)(3) <= CNStageIntLLROutputS1xD(219)(4);
  VNStageIntLLRInputS1xD(366)(3) <= CNStageIntLLROutputS1xD(219)(5);
  VNStageIntLLRInputS1xD(4)(2) <= CNStageIntLLROutputS1xD(220)(0);
  VNStageIntLLRInputS1xD(79)(3) <= CNStageIntLLROutputS1xD(220)(1);
  VNStageIntLLRInputS1xD(139)(3) <= CNStageIntLLROutputS1xD(220)(2);
  VNStageIntLLRInputS1xD(214)(3) <= CNStageIntLLROutputS1xD(220)(3);
  VNStageIntLLRInputS1xD(301)(3) <= CNStageIntLLROutputS1xD(220)(4);
  VNStageIntLLRInputS1xD(321)(3) <= CNStageIntLLROutputS1xD(220)(5);
  VNStageIntLLRInputS1xD(3)(2) <= CNStageIntLLROutputS1xD(221)(0);
  VNStageIntLLRInputS1xD(74)(3) <= CNStageIntLLROutputS1xD(221)(1);
  VNStageIntLLRInputS1xD(149)(3) <= CNStageIntLLROutputS1xD(221)(2);
  VNStageIntLLRInputS1xD(236)(3) <= CNStageIntLLROutputS1xD(221)(3);
  VNStageIntLLRInputS1xD(319)(3) <= CNStageIntLLROutputS1xD(221)(4);
  VNStageIntLLRInputS1xD(369)(2) <= CNStageIntLLROutputS1xD(221)(5);
  VNStageIntLLRInputS1xD(2)(3) <= CNStageIntLLROutputS1xD(222)(0);
  VNStageIntLLRInputS1xD(84)(3) <= CNStageIntLLROutputS1xD(222)(1);
  VNStageIntLLRInputS1xD(171)(2) <= CNStageIntLLROutputS1xD(222)(2);
  VNStageIntLLRInputS1xD(254)(1) <= CNStageIntLLROutputS1xD(222)(3);
  VNStageIntLLRInputS1xD(304)(3) <= CNStageIntLLROutputS1xD(222)(4);
  VNStageIntLLRInputS1xD(356)(3) <= CNStageIntLLROutputS1xD(222)(5);
  VNStageIntLLRInputS1xD(1)(2) <= CNStageIntLLROutputS1xD(223)(0);
  VNStageIntLLRInputS1xD(106)(2) <= CNStageIntLLROutputS1xD(223)(1);
  VNStageIntLLRInputS1xD(189)(2) <= CNStageIntLLROutputS1xD(223)(2);
  VNStageIntLLRInputS1xD(239)(3) <= CNStageIntLLROutputS1xD(223)(3);
  VNStageIntLLRInputS1xD(291)(3) <= CNStageIntLLROutputS1xD(223)(4);
  VNStageIntLLRInputS1xD(324)(3) <= CNStageIntLLROutputS1xD(223)(5);
  VNStageIntLLRInputS1xD(0)(3) <= CNStageIntLLROutputS1xD(224)(0);
  VNStageIntLLRInputS1xD(93)(3) <= CNStageIntLLROutputS1xD(224)(1);
  VNStageIntLLRInputS1xD(158)(3) <= CNStageIntLLROutputS1xD(224)(2);
  VNStageIntLLRInputS1xD(223)(3) <= CNStageIntLLROutputS1xD(224)(3);
  VNStageIntLLRInputS1xD(288)(3) <= CNStageIntLLROutputS1xD(224)(4);
  VNStageIntLLRInputS1xD(353)(3) <= CNStageIntLLROutputS1xD(224)(5);
  VNStageIntLLRInputS1xD(18)(4) <= CNStageIntLLROutputS1xD(225)(0);
  VNStageIntLLRInputS1xD(110)(4) <= CNStageIntLLROutputS1xD(225)(1);
  VNStageIntLLRInputS1xD(167)(4) <= CNStageIntLLROutputS1xD(225)(2);
  VNStageIntLLRInputS1xD(249)(2) <= CNStageIntLLROutputS1xD(225)(3);
  VNStageIntLLRInputS1xD(311)(3) <= CNStageIntLLROutputS1xD(225)(4);
  VNStageIntLLRInputS1xD(347)(4) <= CNStageIntLLROutputS1xD(225)(5);
  VNStageIntLLRInputS1xD(17)(4) <= CNStageIntLLROutputS1xD(226)(0);
  VNStageIntLLRInputS1xD(102)(4) <= CNStageIntLLROutputS1xD(226)(1);
  VNStageIntLLRInputS1xD(184)(4) <= CNStageIntLLROutputS1xD(226)(2);
  VNStageIntLLRInputS1xD(246)(4) <= CNStageIntLLROutputS1xD(226)(3);
  VNStageIntLLRInputS1xD(282)(4) <= CNStageIntLLROutputS1xD(226)(4);
  VNStageIntLLRInputS1xD(367)(4) <= CNStageIntLLROutputS1xD(226)(5);
  VNStageIntLLRInputS1xD(16)(3) <= CNStageIntLLROutputS1xD(227)(0);
  VNStageIntLLRInputS1xD(119)(3) <= CNStageIntLLROutputS1xD(227)(1);
  VNStageIntLLRInputS1xD(181)(4) <= CNStageIntLLROutputS1xD(227)(2);
  VNStageIntLLRInputS1xD(217)(4) <= CNStageIntLLROutputS1xD(227)(3);
  VNStageIntLLRInputS1xD(302)(4) <= CNStageIntLLROutputS1xD(227)(4);
  VNStageIntLLRInputS1xD(353)(4) <= CNStageIntLLROutputS1xD(227)(5);
  VNStageIntLLRInputS1xD(15)(4) <= CNStageIntLLROutputS1xD(228)(0);
  VNStageIntLLRInputS1xD(116)(3) <= CNStageIntLLROutputS1xD(228)(1);
  VNStageIntLLRInputS1xD(152)(4) <= CNStageIntLLROutputS1xD(228)(2);
  VNStageIntLLRInputS1xD(237)(3) <= CNStageIntLLROutputS1xD(228)(3);
  VNStageIntLLRInputS1xD(288)(4) <= CNStageIntLLROutputS1xD(228)(4);
  VNStageIntLLRInputS1xD(343)(4) <= CNStageIntLLROutputS1xD(228)(5);
  VNStageIntLLRInputS1xD(14)(4) <= CNStageIntLLROutputS1xD(229)(0);
  VNStageIntLLRInputS1xD(87)(4) <= CNStageIntLLROutputS1xD(229)(1);
  VNStageIntLLRInputS1xD(172)(3) <= CNStageIntLLROutputS1xD(229)(2);
  VNStageIntLLRInputS1xD(223)(4) <= CNStageIntLLROutputS1xD(229)(3);
  VNStageIntLLRInputS1xD(278)(3) <= CNStageIntLLROutputS1xD(229)(4);
  VNStageIntLLRInputS1xD(372)(3) <= CNStageIntLLROutputS1xD(229)(5);
  VNStageIntLLRInputS1xD(13)(3) <= CNStageIntLLROutputS1xD(230)(0);
  VNStageIntLLRInputS1xD(107)(3) <= CNStageIntLLROutputS1xD(230)(1);
  VNStageIntLLRInputS1xD(158)(4) <= CNStageIntLLROutputS1xD(230)(2);
  VNStageIntLLRInputS1xD(213)(3) <= CNStageIntLLROutputS1xD(230)(3);
  VNStageIntLLRInputS1xD(307)(4) <= CNStageIntLLROutputS1xD(230)(4);
  VNStageIntLLRInputS1xD(355)(4) <= CNStageIntLLROutputS1xD(230)(5);
  VNStageIntLLRInputS1xD(12)(4) <= CNStageIntLLROutputS1xD(231)(0);
  VNStageIntLLRInputS1xD(93)(4) <= CNStageIntLLROutputS1xD(231)(1);
  VNStageIntLLRInputS1xD(148)(4) <= CNStageIntLLROutputS1xD(231)(2);
  VNStageIntLLRInputS1xD(242)(4) <= CNStageIntLLROutputS1xD(231)(3);
  VNStageIntLLRInputS1xD(290)(4) <= CNStageIntLLROutputS1xD(231)(4);
  VNStageIntLLRInputS1xD(322)(3) <= CNStageIntLLROutputS1xD(231)(5);
  VNStageIntLLRInputS1xD(11)(4) <= CNStageIntLLROutputS1xD(232)(0);
  VNStageIntLLRInputS1xD(83)(4) <= CNStageIntLLROutputS1xD(232)(1);
  VNStageIntLLRInputS1xD(177)(4) <= CNStageIntLLROutputS1xD(232)(2);
  VNStageIntLLRInputS1xD(225)(4) <= CNStageIntLLROutputS1xD(232)(3);
  VNStageIntLLRInputS1xD(257)(4) <= CNStageIntLLROutputS1xD(232)(4);
  VNStageIntLLRInputS1xD(345)(3) <= CNStageIntLLROutputS1xD(232)(5);
  VNStageIntLLRInputS1xD(10)(3) <= CNStageIntLLROutputS1xD(233)(0);
  VNStageIntLLRInputS1xD(112)(4) <= CNStageIntLLROutputS1xD(233)(1);
  VNStageIntLLRInputS1xD(160)(4) <= CNStageIntLLROutputS1xD(233)(2);
  VNStageIntLLRInputS1xD(255)(4) <= CNStageIntLLROutputS1xD(233)(3);
  VNStageIntLLRInputS1xD(280)(4) <= CNStageIntLLROutputS1xD(233)(4);
  VNStageIntLLRInputS1xD(381)(3) <= CNStageIntLLROutputS1xD(233)(5);
  VNStageIntLLRInputS1xD(9)(4) <= CNStageIntLLROutputS1xD(234)(0);
  VNStageIntLLRInputS1xD(95)(4) <= CNStageIntLLROutputS1xD(234)(1);
  VNStageIntLLRInputS1xD(190)(2) <= CNStageIntLLROutputS1xD(234)(2);
  VNStageIntLLRInputS1xD(215)(4) <= CNStageIntLLROutputS1xD(234)(3);
  VNStageIntLLRInputS1xD(316)(2) <= CNStageIntLLROutputS1xD(234)(4);
  VNStageIntLLRInputS1xD(365)(4) <= CNStageIntLLROutputS1xD(234)(5);
  VNStageIntLLRInputS1xD(7)(4) <= CNStageIntLLROutputS1xD(235)(0);
  VNStageIntLLRInputS1xD(85)(3) <= CNStageIntLLROutputS1xD(235)(1);
  VNStageIntLLRInputS1xD(186)(3) <= CNStageIntLLROutputS1xD(235)(2);
  VNStageIntLLRInputS1xD(235)(3) <= CNStageIntLLROutputS1xD(235)(3);
  VNStageIntLLRInputS1xD(303)(4) <= CNStageIntLLROutputS1xD(235)(4);
  VNStageIntLLRInputS1xD(346)(4) <= CNStageIntLLROutputS1xD(235)(5);
  VNStageIntLLRInputS1xD(6)(4) <= CNStageIntLLROutputS1xD(236)(0);
  VNStageIntLLRInputS1xD(121)(3) <= CNStageIntLLROutputS1xD(236)(1);
  VNStageIntLLRInputS1xD(170)(3) <= CNStageIntLLROutputS1xD(236)(2);
  VNStageIntLLRInputS1xD(238)(4) <= CNStageIntLLROutputS1xD(236)(3);
  VNStageIntLLRInputS1xD(281)(4) <= CNStageIntLLROutputS1xD(236)(4);
  VNStageIntLLRInputS1xD(321)(4) <= CNStageIntLLROutputS1xD(236)(5);
  VNStageIntLLRInputS1xD(5)(4) <= CNStageIntLLROutputS1xD(237)(0);
  VNStageIntLLRInputS1xD(105)(3) <= CNStageIntLLROutputS1xD(237)(1);
  VNStageIntLLRInputS1xD(173)(4) <= CNStageIntLLROutputS1xD(237)(2);
  VNStageIntLLRInputS1xD(216)(4) <= CNStageIntLLROutputS1xD(237)(3);
  VNStageIntLLRInputS1xD(319)(4) <= CNStageIntLLROutputS1xD(237)(4);
  VNStageIntLLRInputS1xD(382)(3) <= CNStageIntLLROutputS1xD(237)(5);
  VNStageIntLLRInputS1xD(4)(3) <= CNStageIntLLROutputS1xD(238)(0);
  VNStageIntLLRInputS1xD(108)(4) <= CNStageIntLLROutputS1xD(238)(1);
  VNStageIntLLRInputS1xD(151)(4) <= CNStageIntLLROutputS1xD(238)(2);
  VNStageIntLLRInputS1xD(254)(2) <= CNStageIntLLROutputS1xD(238)(3);
  VNStageIntLLRInputS1xD(317)(1) <= CNStageIntLLROutputS1xD(238)(4);
  VNStageIntLLRInputS1xD(344)(4) <= CNStageIntLLROutputS1xD(238)(5);
  VNStageIntLLRInputS1xD(3)(3) <= CNStageIntLLROutputS1xD(239)(0);
  VNStageIntLLRInputS1xD(86)(2) <= CNStageIntLLROutputS1xD(239)(1);
  VNStageIntLLRInputS1xD(189)(3) <= CNStageIntLLROutputS1xD(239)(2);
  VNStageIntLLRInputS1xD(252)(3) <= CNStageIntLLROutputS1xD(239)(3);
  VNStageIntLLRInputS1xD(279)(4) <= CNStageIntLLROutputS1xD(239)(4);
  VNStageIntLLRInputS1xD(352)(4) <= CNStageIntLLROutputS1xD(239)(5);
  VNStageIntLLRInputS1xD(2)(4) <= CNStageIntLLROutputS1xD(240)(0);
  VNStageIntLLRInputS1xD(124)(2) <= CNStageIntLLROutputS1xD(240)(1);
  VNStageIntLLRInputS1xD(187)(3) <= CNStageIntLLROutputS1xD(240)(2);
  VNStageIntLLRInputS1xD(214)(4) <= CNStageIntLLROutputS1xD(240)(3);
  VNStageIntLLRInputS1xD(287)(4) <= CNStageIntLLROutputS1xD(240)(4);
  VNStageIntLLRInputS1xD(332)(4) <= CNStageIntLLROutputS1xD(240)(5);
  VNStageIntLLRInputS1xD(1)(3) <= CNStageIntLLROutputS1xD(241)(0);
  VNStageIntLLRInputS1xD(122)(3) <= CNStageIntLLROutputS1xD(241)(1);
  VNStageIntLLRInputS1xD(149)(4) <= CNStageIntLLROutputS1xD(241)(2);
  VNStageIntLLRInputS1xD(222)(2) <= CNStageIntLLROutputS1xD(241)(3);
  VNStageIntLLRInputS1xD(267)(4) <= CNStageIntLLROutputS1xD(241)(4);
  VNStageIntLLRInputS1xD(326)(3) <= CNStageIntLLROutputS1xD(241)(5);
  VNStageIntLLRInputS1xD(62)(3) <= CNStageIntLLROutputS1xD(242)(0);
  VNStageIntLLRInputS1xD(92)(4) <= CNStageIntLLROutputS1xD(242)(1);
  VNStageIntLLRInputS1xD(137)(4) <= CNStageIntLLROutputS1xD(242)(2);
  VNStageIntLLRInputS1xD(196)(4) <= CNStageIntLLROutputS1xD(242)(3);
  VNStageIntLLRInputS1xD(256)(3) <= CNStageIntLLROutputS1xD(242)(4);
  VNStageIntLLRInputS1xD(325)(4) <= CNStageIntLLROutputS1xD(242)(5);
  VNStageIntLLRInputS1xD(61)(3) <= CNStageIntLLROutputS1xD(243)(0);
  VNStageIntLLRInputS1xD(72)(4) <= CNStageIntLLROutputS1xD(243)(1);
  VNStageIntLLRInputS1xD(131)(3) <= CNStageIntLLROutputS1xD(243)(2);
  VNStageIntLLRInputS1xD(192)(4) <= CNStageIntLLROutputS1xD(243)(3);
  VNStageIntLLRInputS1xD(260)(4) <= CNStageIntLLROutputS1xD(243)(4);
  VNStageIntLLRInputS1xD(330)(4) <= CNStageIntLLROutputS1xD(243)(5);
  VNStageIntLLRInputS1xD(60)(3) <= CNStageIntLLROutputS1xD(244)(0);
  VNStageIntLLRInputS1xD(66)(3) <= CNStageIntLLROutputS1xD(244)(1);
  VNStageIntLLRInputS1xD(128)(4) <= CNStageIntLLROutputS1xD(244)(2);
  VNStageIntLLRInputS1xD(195)(3) <= CNStageIntLLROutputS1xD(244)(3);
  VNStageIntLLRInputS1xD(265)(3) <= CNStageIntLLROutputS1xD(244)(4);
  VNStageIntLLRInputS1xD(349)(3) <= CNStageIntLLROutputS1xD(244)(5);
  VNStageIntLLRInputS1xD(59)(2) <= CNStageIntLLROutputS1xD(245)(0);
  VNStageIntLLRInputS1xD(64)(3) <= CNStageIntLLROutputS1xD(245)(1);
  VNStageIntLLRInputS1xD(130)(4) <= CNStageIntLLROutputS1xD(245)(2);
  VNStageIntLLRInputS1xD(200)(4) <= CNStageIntLLROutputS1xD(245)(3);
  VNStageIntLLRInputS1xD(284)(4) <= CNStageIntLLROutputS1xD(245)(4);
  VNStageIntLLRInputS1xD(340)(4) <= CNStageIntLLROutputS1xD(245)(5);
  VNStageIntLLRInputS1xD(57)(3) <= CNStageIntLLROutputS1xD(246)(0);
  VNStageIntLLRInputS1xD(70)(4) <= CNStageIntLLROutputS1xD(246)(1);
  VNStageIntLLRInputS1xD(154)(3) <= CNStageIntLLROutputS1xD(246)(2);
  VNStageIntLLRInputS1xD(210)(4) <= CNStageIntLLROutputS1xD(246)(3);
  VNStageIntLLRInputS1xD(312)(3) <= CNStageIntLLROutputS1xD(246)(4);
  VNStageIntLLRInputS1xD(378)(3) <= CNStageIntLLROutputS1xD(246)(5);
  VNStageIntLLRInputS1xD(56)(4) <= CNStageIntLLROutputS1xD(247)(0);
  VNStageIntLLRInputS1xD(89)(4) <= CNStageIntLLROutputS1xD(247)(1);
  VNStageIntLLRInputS1xD(145)(4) <= CNStageIntLLROutputS1xD(247)(2);
  VNStageIntLLRInputS1xD(247)(4) <= CNStageIntLLROutputS1xD(247)(3);
  VNStageIntLLRInputS1xD(313)(2) <= CNStageIntLLROutputS1xD(247)(4);
  VNStageIntLLRInputS1xD(339)(4) <= CNStageIntLLROutputS1xD(247)(5);
  VNStageIntLLRInputS1xD(55)(4) <= CNStageIntLLROutputS1xD(248)(0);
  VNStageIntLLRInputS1xD(80)(4) <= CNStageIntLLROutputS1xD(248)(1);
  VNStageIntLLRInputS1xD(182)(4) <= CNStageIntLLROutputS1xD(248)(2);
  VNStageIntLLRInputS1xD(248)(4) <= CNStageIntLLROutputS1xD(248)(3);
  VNStageIntLLRInputS1xD(274)(3) <= CNStageIntLLROutputS1xD(248)(4);
  VNStageIntLLRInputS1xD(360)(4) <= CNStageIntLLROutputS1xD(248)(5);
  VNStageIntLLRInputS1xD(53)(3) <= CNStageIntLLROutputS1xD(249)(0);
  VNStageIntLLRInputS1xD(118)(3) <= CNStageIntLLROutputS1xD(249)(1);
  VNStageIntLLRInputS1xD(144)(4) <= CNStageIntLLROutputS1xD(249)(2);
  VNStageIntLLRInputS1xD(230)(3) <= CNStageIntLLROutputS1xD(249)(3);
  VNStageIntLLRInputS1xD(291)(4) <= CNStageIntLLROutputS1xD(249)(4);
  VNStageIntLLRInputS1xD(371)(3) <= CNStageIntLLROutputS1xD(249)(5);
  VNStageIntLLRInputS1xD(51)(3) <= CNStageIntLLROutputS1xD(250)(0);
  VNStageIntLLRInputS1xD(100)(4) <= CNStageIntLLROutputS1xD(250)(1);
  VNStageIntLLRInputS1xD(161)(4) <= CNStageIntLLROutputS1xD(250)(2);
  VNStageIntLLRInputS1xD(241)(3) <= CNStageIntLLROutputS1xD(250)(3);
  VNStageIntLLRInputS1xD(269)(3) <= CNStageIntLLROutputS1xD(250)(4);
  VNStageIntLLRInputS1xD(373)(2) <= CNStageIntLLROutputS1xD(250)(5);
  VNStageIntLLRInputS1xD(50)(4) <= CNStageIntLLROutputS1xD(251)(0);
  VNStageIntLLRInputS1xD(96)(4) <= CNStageIntLLROutputS1xD(251)(1);
  VNStageIntLLRInputS1xD(176)(4) <= CNStageIntLLROutputS1xD(251)(2);
  VNStageIntLLRInputS1xD(204)(4) <= CNStageIntLLROutputS1xD(251)(3);
  VNStageIntLLRInputS1xD(308)(2) <= CNStageIntLLROutputS1xD(251)(4);
  VNStageIntLLRInputS1xD(342)(3) <= CNStageIntLLROutputS1xD(251)(5);
  VNStageIntLLRInputS1xD(49)(4) <= CNStageIntLLROutputS1xD(252)(0);
  VNStageIntLLRInputS1xD(111)(4) <= CNStageIntLLROutputS1xD(252)(1);
  VNStageIntLLRInputS1xD(139)(4) <= CNStageIntLLROutputS1xD(252)(2);
  VNStageIntLLRInputS1xD(243)(4) <= CNStageIntLLROutputS1xD(252)(3);
  VNStageIntLLRInputS1xD(277)(4) <= CNStageIntLLROutputS1xD(252)(4);
  VNStageIntLLRInputS1xD(358)(3) <= CNStageIntLLROutputS1xD(252)(5);
  VNStageIntLLRInputS1xD(47)(2) <= CNStageIntLLROutputS1xD(253)(0);
  VNStageIntLLRInputS1xD(113)(4) <= CNStageIntLLROutputS1xD(253)(1);
  VNStageIntLLRInputS1xD(147)(4) <= CNStageIntLLROutputS1xD(253)(2);
  VNStageIntLLRInputS1xD(228)(4) <= CNStageIntLLROutputS1xD(253)(3);
  VNStageIntLLRInputS1xD(263)(4) <= CNStageIntLLROutputS1xD(253)(4);
  VNStageIntLLRInputS1xD(337)(4) <= CNStageIntLLROutputS1xD(253)(5);
  VNStageIntLLRInputS1xD(46)(4) <= CNStageIntLLROutputS1xD(254)(0);
  VNStageIntLLRInputS1xD(82)(4) <= CNStageIntLLROutputS1xD(254)(1);
  VNStageIntLLRInputS1xD(163)(3) <= CNStageIntLLROutputS1xD(254)(2);
  VNStageIntLLRInputS1xD(198)(4) <= CNStageIntLLROutputS1xD(254)(3);
  VNStageIntLLRInputS1xD(272)(4) <= CNStageIntLLROutputS1xD(254)(4);
  VNStageIntLLRInputS1xD(350)(4) <= CNStageIntLLROutputS1xD(254)(5);
  VNStageIntLLRInputS1xD(45)(4) <= CNStageIntLLROutputS1xD(255)(0);
  VNStageIntLLRInputS1xD(98)(3) <= CNStageIntLLROutputS1xD(255)(1);
  VNStageIntLLRInputS1xD(133)(2) <= CNStageIntLLROutputS1xD(255)(2);
  VNStageIntLLRInputS1xD(207)(3) <= CNStageIntLLROutputS1xD(255)(3);
  VNStageIntLLRInputS1xD(285)(4) <= CNStageIntLLROutputS1xD(255)(4);
  VNStageIntLLRInputS1xD(329)(4) <= CNStageIntLLROutputS1xD(255)(5);
  VNStageIntLLRInputS1xD(44)(4) <= CNStageIntLLROutputS1xD(256)(0);
  VNStageIntLLRInputS1xD(68)(3) <= CNStageIntLLROutputS1xD(256)(1);
  VNStageIntLLRInputS1xD(142)(3) <= CNStageIntLLROutputS1xD(256)(2);
  VNStageIntLLRInputS1xD(220)(4) <= CNStageIntLLROutputS1xD(256)(3);
  VNStageIntLLRInputS1xD(264)(4) <= CNStageIntLLROutputS1xD(256)(4);
  VNStageIntLLRInputS1xD(357)(4) <= CNStageIntLLROutputS1xD(256)(5);
  VNStageIntLLRInputS1xD(43)(3) <= CNStageIntLLROutputS1xD(257)(0);
  VNStageIntLLRInputS1xD(77)(2) <= CNStageIntLLROutputS1xD(257)(1);
  VNStageIntLLRInputS1xD(155)(4) <= CNStageIntLLROutputS1xD(257)(2);
  VNStageIntLLRInputS1xD(199)(4) <= CNStageIntLLROutputS1xD(257)(3);
  VNStageIntLLRInputS1xD(292)(4) <= CNStageIntLLROutputS1xD(257)(4);
  VNStageIntLLRInputS1xD(359)(4) <= CNStageIntLLROutputS1xD(257)(5);
  VNStageIntLLRInputS1xD(42)(4) <= CNStageIntLLROutputS1xD(258)(0);
  VNStageIntLLRInputS1xD(90)(4) <= CNStageIntLLROutputS1xD(258)(1);
  VNStageIntLLRInputS1xD(134)(3) <= CNStageIntLLROutputS1xD(258)(2);
  VNStageIntLLRInputS1xD(227)(4) <= CNStageIntLLROutputS1xD(258)(3);
  VNStageIntLLRInputS1xD(294)(4) <= CNStageIntLLROutputS1xD(258)(4);
  VNStageIntLLRInputS1xD(341)(4) <= CNStageIntLLROutputS1xD(258)(5);
  VNStageIntLLRInputS1xD(41)(4) <= CNStageIntLLROutputS1xD(259)(0);
  VNStageIntLLRInputS1xD(69)(4) <= CNStageIntLLROutputS1xD(259)(1);
  VNStageIntLLRInputS1xD(162)(4) <= CNStageIntLLROutputS1xD(259)(2);
  VNStageIntLLRInputS1xD(229)(3) <= CNStageIntLLROutputS1xD(259)(3);
  VNStageIntLLRInputS1xD(276)(4) <= CNStageIntLLROutputS1xD(259)(4);
  VNStageIntLLRInputS1xD(348)(4) <= CNStageIntLLROutputS1xD(259)(5);
  VNStageIntLLRInputS1xD(40)(3) <= CNStageIntLLROutputS1xD(260)(0);
  VNStageIntLLRInputS1xD(97)(4) <= CNStageIntLLROutputS1xD(260)(1);
  VNStageIntLLRInputS1xD(164)(4) <= CNStageIntLLROutputS1xD(260)(2);
  VNStageIntLLRInputS1xD(211)(4) <= CNStageIntLLROutputS1xD(260)(3);
  VNStageIntLLRInputS1xD(283)(4) <= CNStageIntLLROutputS1xD(260)(4);
  VNStageIntLLRInputS1xD(375)(3) <= CNStageIntLLROutputS1xD(260)(5);
  VNStageIntLLRInputS1xD(39)(4) <= CNStageIntLLROutputS1xD(261)(0);
  VNStageIntLLRInputS1xD(99)(4) <= CNStageIntLLROutputS1xD(261)(1);
  VNStageIntLLRInputS1xD(146)(3) <= CNStageIntLLROutputS1xD(261)(2);
  VNStageIntLLRInputS1xD(218)(4) <= CNStageIntLLROutputS1xD(261)(3);
  VNStageIntLLRInputS1xD(310)(3) <= CNStageIntLLROutputS1xD(261)(4);
  VNStageIntLLRInputS1xD(363)(3) <= CNStageIntLLROutputS1xD(261)(5);
  VNStageIntLLRInputS1xD(38)(4) <= CNStageIntLLROutputS1xD(262)(0);
  VNStageIntLLRInputS1xD(81)(3) <= CNStageIntLLROutputS1xD(262)(1);
  VNStageIntLLRInputS1xD(153)(4) <= CNStageIntLLROutputS1xD(262)(2);
  VNStageIntLLRInputS1xD(245)(4) <= CNStageIntLLROutputS1xD(262)(3);
  VNStageIntLLRInputS1xD(298)(4) <= CNStageIntLLROutputS1xD(262)(4);
  VNStageIntLLRInputS1xD(369)(3) <= CNStageIntLLROutputS1xD(262)(5);
  VNStageIntLLRInputS1xD(37)(4) <= CNStageIntLLROutputS1xD(263)(0);
  VNStageIntLLRInputS1xD(88)(4) <= CNStageIntLLROutputS1xD(263)(1);
  VNStageIntLLRInputS1xD(180)(2) <= CNStageIntLLROutputS1xD(263)(2);
  VNStageIntLLRInputS1xD(233)(3) <= CNStageIntLLROutputS1xD(263)(3);
  VNStageIntLLRInputS1xD(304)(4) <= CNStageIntLLROutputS1xD(263)(4);
  VNStageIntLLRInputS1xD(364)(4) <= CNStageIntLLROutputS1xD(263)(5);
  VNStageIntLLRInputS1xD(36)(3) <= CNStageIntLLROutputS1xD(264)(0);
  VNStageIntLLRInputS1xD(115)(4) <= CNStageIntLLROutputS1xD(264)(1);
  VNStageIntLLRInputS1xD(168)(3) <= CNStageIntLLROutputS1xD(264)(2);
  VNStageIntLLRInputS1xD(239)(4) <= CNStageIntLLROutputS1xD(264)(3);
  VNStageIntLLRInputS1xD(299)(3) <= CNStageIntLLROutputS1xD(264)(4);
  VNStageIntLLRInputS1xD(374)(4) <= CNStageIntLLROutputS1xD(264)(5);
  VNStageIntLLRInputS1xD(35)(4) <= CNStageIntLLROutputS1xD(265)(0);
  VNStageIntLLRInputS1xD(103)(4) <= CNStageIntLLROutputS1xD(265)(1);
  VNStageIntLLRInputS1xD(174)(3) <= CNStageIntLLROutputS1xD(265)(2);
  VNStageIntLLRInputS1xD(234)(4) <= CNStageIntLLROutputS1xD(265)(3);
  VNStageIntLLRInputS1xD(309)(4) <= CNStageIntLLROutputS1xD(265)(4);
  VNStageIntLLRInputS1xD(333)(3) <= CNStageIntLLROutputS1xD(265)(5);
  VNStageIntLLRInputS1xD(34)(4) <= CNStageIntLLROutputS1xD(266)(0);
  VNStageIntLLRInputS1xD(109)(4) <= CNStageIntLLROutputS1xD(266)(1);
  VNStageIntLLRInputS1xD(169)(4) <= CNStageIntLLROutputS1xD(266)(2);
  VNStageIntLLRInputS1xD(244)(1) <= CNStageIntLLROutputS1xD(266)(3);
  VNStageIntLLRInputS1xD(268)(4) <= CNStageIntLLROutputS1xD(266)(4);
  VNStageIntLLRInputS1xD(351)(3) <= CNStageIntLLROutputS1xD(266)(5);
  VNStageIntLLRInputS1xD(33)(4) <= CNStageIntLLROutputS1xD(267)(0);
  VNStageIntLLRInputS1xD(104)(4) <= CNStageIntLLROutputS1xD(267)(1);
  VNStageIntLLRInputS1xD(179)(4) <= CNStageIntLLROutputS1xD(267)(2);
  VNStageIntLLRInputS1xD(203)(4) <= CNStageIntLLROutputS1xD(267)(3);
  VNStageIntLLRInputS1xD(286)(4) <= CNStageIntLLROutputS1xD(267)(4);
  VNStageIntLLRInputS1xD(336)(3) <= CNStageIntLLROutputS1xD(267)(5);
  VNStageIntLLRInputS1xD(32)(3) <= CNStageIntLLROutputS1xD(268)(0);
  VNStageIntLLRInputS1xD(114)(4) <= CNStageIntLLROutputS1xD(268)(1);
  VNStageIntLLRInputS1xD(138)(4) <= CNStageIntLLROutputS1xD(268)(2);
  VNStageIntLLRInputS1xD(221)(4) <= CNStageIntLLROutputS1xD(268)(3);
  VNStageIntLLRInputS1xD(271)(3) <= CNStageIntLLROutputS1xD(268)(4);
  VNStageIntLLRInputS1xD(323)(3) <= CNStageIntLLROutputS1xD(268)(5);
  VNStageIntLLRInputS1xD(30)(4) <= CNStageIntLLROutputS1xD(269)(0);
  VNStageIntLLRInputS1xD(91)(4) <= CNStageIntLLROutputS1xD(269)(1);
  VNStageIntLLRInputS1xD(141)(2) <= CNStageIntLLROutputS1xD(269)(2);
  VNStageIntLLRInputS1xD(193)(3) <= CNStageIntLLROutputS1xD(269)(3);
  VNStageIntLLRInputS1xD(289)(4) <= CNStageIntLLROutputS1xD(269)(4);
  VNStageIntLLRInputS1xD(366)(4) <= CNStageIntLLROutputS1xD(269)(5);
  VNStageIntLLRInputS1xD(29)(3) <= CNStageIntLLROutputS1xD(270)(0);
  VNStageIntLLRInputS1xD(76)(4) <= CNStageIntLLROutputS1xD(270)(1);
  VNStageIntLLRInputS1xD(191)(4) <= CNStageIntLLROutputS1xD(270)(2);
  VNStageIntLLRInputS1xD(224)(4) <= CNStageIntLLROutputS1xD(270)(3);
  VNStageIntLLRInputS1xD(301)(4) <= CNStageIntLLROutputS1xD(270)(4);
  VNStageIntLLRInputS1xD(380)(3) <= CNStageIntLLROutputS1xD(270)(5);
  VNStageIntLLRInputS1xD(28)(4) <= CNStageIntLLROutputS1xD(271)(0);
  VNStageIntLLRInputS1xD(126)(3) <= CNStageIntLLROutputS1xD(271)(1);
  VNStageIntLLRInputS1xD(159)(3) <= CNStageIntLLROutputS1xD(271)(2);
  VNStageIntLLRInputS1xD(236)(4) <= CNStageIntLLROutputS1xD(271)(3);
  VNStageIntLLRInputS1xD(315)(3) <= CNStageIntLLROutputS1xD(271)(4);
  VNStageIntLLRInputS1xD(361)(4) <= CNStageIntLLROutputS1xD(271)(5);
  VNStageIntLLRInputS1xD(26)(4) <= CNStageIntLLROutputS1xD(272)(0);
  VNStageIntLLRInputS1xD(106)(3) <= CNStageIntLLROutputS1xD(272)(1);
  VNStageIntLLRInputS1xD(185)(1) <= CNStageIntLLROutputS1xD(272)(2);
  VNStageIntLLRInputS1xD(231)(3) <= CNStageIntLLROutputS1xD(272)(3);
  VNStageIntLLRInputS1xD(273)(3) <= CNStageIntLLROutputS1xD(272)(4);
  VNStageIntLLRInputS1xD(327)(4) <= CNStageIntLLROutputS1xD(272)(5);
  VNStageIntLLRInputS1xD(24)(4) <= CNStageIntLLROutputS1xD(273)(0);
  VNStageIntLLRInputS1xD(101)(4) <= CNStageIntLLROutputS1xD(273)(1);
  VNStageIntLLRInputS1xD(143)(4) <= CNStageIntLLROutputS1xD(273)(2);
  VNStageIntLLRInputS1xD(197)(4) <= CNStageIntLLROutputS1xD(273)(3);
  VNStageIntLLRInputS1xD(266)(3) <= CNStageIntLLROutputS1xD(273)(4);
  VNStageIntLLRInputS1xD(324)(4) <= CNStageIntLLROutputS1xD(273)(5);
  VNStageIntLLRInputS1xD(23)(4) <= CNStageIntLLROutputS1xD(274)(0);
  VNStageIntLLRInputS1xD(78)(4) <= CNStageIntLLROutputS1xD(274)(1);
  VNStageIntLLRInputS1xD(132)(3) <= CNStageIntLLROutputS1xD(274)(2);
  VNStageIntLLRInputS1xD(201)(4) <= CNStageIntLLROutputS1xD(274)(3);
  VNStageIntLLRInputS1xD(259)(2) <= CNStageIntLLROutputS1xD(274)(4);
  VNStageIntLLRInputS1xD(335)(4) <= CNStageIntLLROutputS1xD(274)(5);
  VNStageIntLLRInputS1xD(22)(4) <= CNStageIntLLROutputS1xD(275)(0);
  VNStageIntLLRInputS1xD(67)(1) <= CNStageIntLLROutputS1xD(275)(1);
  VNStageIntLLRInputS1xD(136)(4) <= CNStageIntLLROutputS1xD(275)(2);
  VNStageIntLLRInputS1xD(194)(4) <= CNStageIntLLROutputS1xD(275)(3);
  VNStageIntLLRInputS1xD(270)(4) <= CNStageIntLLROutputS1xD(275)(4);
  VNStageIntLLRInputS1xD(370)(3) <= CNStageIntLLROutputS1xD(275)(5);
  VNStageIntLLRInputS1xD(21)(4) <= CNStageIntLLROutputS1xD(276)(0);
  VNStageIntLLRInputS1xD(71)(3) <= CNStageIntLLROutputS1xD(276)(1);
  VNStageIntLLRInputS1xD(129)(4) <= CNStageIntLLROutputS1xD(276)(2);
  VNStageIntLLRInputS1xD(205)(1) <= CNStageIntLLROutputS1xD(276)(3);
  VNStageIntLLRInputS1xD(305)(4) <= CNStageIntLLROutputS1xD(276)(4);
  VNStageIntLLRInputS1xD(362)(4) <= CNStageIntLLROutputS1xD(276)(5);
  VNStageIntLLRInputS1xD(20)(2) <= CNStageIntLLROutputS1xD(277)(0);
  VNStageIntLLRInputS1xD(127)(4) <= CNStageIntLLROutputS1xD(277)(1);
  VNStageIntLLRInputS1xD(140)(4) <= CNStageIntLLROutputS1xD(277)(2);
  VNStageIntLLRInputS1xD(240)(4) <= CNStageIntLLROutputS1xD(277)(3);
  VNStageIntLLRInputS1xD(297)(4) <= CNStageIntLLROutputS1xD(277)(4);
  VNStageIntLLRInputS1xD(379)(2) <= CNStageIntLLROutputS1xD(277)(5);
  VNStageIntLLRInputS1xD(19)(3) <= CNStageIntLLROutputS1xD(278)(0);
  VNStageIntLLRInputS1xD(75)(4) <= CNStageIntLLROutputS1xD(278)(1);
  VNStageIntLLRInputS1xD(175)(4) <= CNStageIntLLROutputS1xD(278)(2);
  VNStageIntLLRInputS1xD(232)(3) <= CNStageIntLLROutputS1xD(278)(3);
  VNStageIntLLRInputS1xD(314)(1) <= CNStageIntLLROutputS1xD(278)(4);
  VNStageIntLLRInputS1xD(376)(3) <= CNStageIntLLROutputS1xD(278)(5);
  VNStageIntLLRInputS1xD(0)(4) <= CNStageIntLLROutputS1xD(279)(0);
  VNStageIntLLRInputS1xD(123)(3) <= CNStageIntLLROutputS1xD(279)(1);
  VNStageIntLLRInputS1xD(188)(2) <= CNStageIntLLROutputS1xD(279)(2);
  VNStageIntLLRInputS1xD(253)(3) <= CNStageIntLLROutputS1xD(279)(3);
  VNStageIntLLRInputS1xD(318)(2) <= CNStageIntLLROutputS1xD(279)(4);
  VNStageIntLLRInputS1xD(383)(4) <= CNStageIntLLROutputS1xD(279)(5);
  VNStageIntLLRInputS1xD(35)(5) <= CNStageIntLLROutputS1xD(280)(0);
  VNStageIntLLRInputS1xD(91)(5) <= CNStageIntLLROutputS1xD(280)(1);
  VNStageIntLLRInputS1xD(191)(5) <= CNStageIntLLROutputS1xD(280)(2);
  VNStageIntLLRInputS1xD(248)(5) <= CNStageIntLLROutputS1xD(280)(3);
  VNStageIntLLRInputS1xD(267)(5) <= CNStageIntLLROutputS1xD(280)(4);
  VNStageIntLLRInputS1xD(329)(5) <= CNStageIntLLROutputS1xD(280)(5);
  VNStageIntLLRInputS1xD(34)(5) <= CNStageIntLLROutputS1xD(281)(0);
  VNStageIntLLRInputS1xD(126)(4) <= CNStageIntLLROutputS1xD(281)(1);
  VNStageIntLLRInputS1xD(183)(3) <= CNStageIntLLROutputS1xD(281)(2);
  VNStageIntLLRInputS1xD(202)(4) <= CNStageIntLLROutputS1xD(281)(3);
  VNStageIntLLRInputS1xD(264)(5) <= CNStageIntLLROutputS1xD(281)(4);
  VNStageIntLLRInputS1xD(363)(4) <= CNStageIntLLROutputS1xD(281)(5);
  VNStageIntLLRInputS1xD(33)(5) <= CNStageIntLLROutputS1xD(282)(0);
  VNStageIntLLRInputS1xD(118)(4) <= CNStageIntLLROutputS1xD(282)(1);
  VNStageIntLLRInputS1xD(137)(5) <= CNStageIntLLROutputS1xD(282)(2);
  VNStageIntLLRInputS1xD(199)(5) <= CNStageIntLLROutputS1xD(282)(3);
  VNStageIntLLRInputS1xD(298)(5) <= CNStageIntLLROutputS1xD(282)(4);
  VNStageIntLLRInputS1xD(383)(5) <= CNStageIntLLROutputS1xD(282)(5);
  VNStageIntLLRInputS1xD(31)(3) <= CNStageIntLLROutputS1xD(283)(0);
  VNStageIntLLRInputS1xD(69)(5) <= CNStageIntLLROutputS1xD(283)(1);
  VNStageIntLLRInputS1xD(168)(4) <= CNStageIntLLROutputS1xD(283)(2);
  VNStageIntLLRInputS1xD(253)(4) <= CNStageIntLLROutputS1xD(283)(3);
  VNStageIntLLRInputS1xD(304)(5) <= CNStageIntLLROutputS1xD(283)(4);
  VNStageIntLLRInputS1xD(359)(5) <= CNStageIntLLROutputS1xD(283)(5);
  VNStageIntLLRInputS1xD(30)(5) <= CNStageIntLLROutputS1xD(284)(0);
  VNStageIntLLRInputS1xD(103)(5) <= CNStageIntLLROutputS1xD(284)(1);
  VNStageIntLLRInputS1xD(188)(3) <= CNStageIntLLROutputS1xD(284)(2);
  VNStageIntLLRInputS1xD(239)(5) <= CNStageIntLLROutputS1xD(284)(3);
  VNStageIntLLRInputS1xD(294)(5) <= CNStageIntLLROutputS1xD(284)(4);
  VNStageIntLLRInputS1xD(325)(5) <= CNStageIntLLROutputS1xD(284)(5);
  VNStageIntLLRInputS1xD(27)(4) <= CNStageIntLLROutputS1xD(285)(0);
  VNStageIntLLRInputS1xD(99)(5) <= CNStageIntLLROutputS1xD(285)(1);
  VNStageIntLLRInputS1xD(130)(5) <= CNStageIntLLROutputS1xD(285)(2);
  VNStageIntLLRInputS1xD(241)(4) <= CNStageIntLLROutputS1xD(285)(3);
  VNStageIntLLRInputS1xD(273)(4) <= CNStageIntLLROutputS1xD(285)(4);
  VNStageIntLLRInputS1xD(361)(5) <= CNStageIntLLROutputS1xD(285)(5);
  VNStageIntLLRInputS1xD(26)(5) <= CNStageIntLLROutputS1xD(286)(0);
  VNStageIntLLRInputS1xD(65)(4) <= CNStageIntLLROutputS1xD(286)(1);
  VNStageIntLLRInputS1xD(176)(5) <= CNStageIntLLROutputS1xD(286)(2);
  VNStageIntLLRInputS1xD(208)(4) <= CNStageIntLLROutputS1xD(286)(3);
  VNStageIntLLRInputS1xD(296)(4) <= CNStageIntLLROutputS1xD(286)(4);
  VNStageIntLLRInputS1xD(334)(3) <= CNStageIntLLROutputS1xD(286)(5);
  VNStageIntLLRInputS1xD(25)(4) <= CNStageIntLLROutputS1xD(287)(0);
  VNStageIntLLRInputS1xD(111)(5) <= CNStageIntLLROutputS1xD(287)(1);
  VNStageIntLLRInputS1xD(143)(5) <= CNStageIntLLROutputS1xD(287)(2);
  VNStageIntLLRInputS1xD(231)(4) <= CNStageIntLLROutputS1xD(287)(3);
  VNStageIntLLRInputS1xD(269)(4) <= CNStageIntLLROutputS1xD(287)(4);
  VNStageIntLLRInputS1xD(381)(4) <= CNStageIntLLROutputS1xD(287)(5);
  VNStageIntLLRInputS1xD(24)(5) <= CNStageIntLLROutputS1xD(288)(0);
  VNStageIntLLRInputS1xD(78)(5) <= CNStageIntLLROutputS1xD(288)(1);
  VNStageIntLLRInputS1xD(166)(4) <= CNStageIntLLROutputS1xD(288)(2);
  VNStageIntLLRInputS1xD(204)(5) <= CNStageIntLLROutputS1xD(288)(3);
  VNStageIntLLRInputS1xD(316)(3) <= CNStageIntLLROutputS1xD(288)(4);
  VNStageIntLLRInputS1xD(321)(5) <= CNStageIntLLROutputS1xD(288)(5);
  VNStageIntLLRInputS1xD(23)(5) <= CNStageIntLLROutputS1xD(289)(0);
  VNStageIntLLRInputS1xD(101)(5) <= CNStageIntLLROutputS1xD(289)(1);
  VNStageIntLLRInputS1xD(139)(5) <= CNStageIntLLROutputS1xD(289)(2);
  VNStageIntLLRInputS1xD(251)(3) <= CNStageIntLLROutputS1xD(289)(3);
  VNStageIntLLRInputS1xD(319)(5) <= CNStageIntLLROutputS1xD(289)(4);
  VNStageIntLLRInputS1xD(362)(5) <= CNStageIntLLROutputS1xD(289)(5);
  VNStageIntLLRInputS1xD(22)(5) <= CNStageIntLLROutputS1xD(290)(0);
  VNStageIntLLRInputS1xD(74)(4) <= CNStageIntLLROutputS1xD(290)(1);
  VNStageIntLLRInputS1xD(186)(4) <= CNStageIntLLROutputS1xD(290)(2);
  VNStageIntLLRInputS1xD(254)(3) <= CNStageIntLLROutputS1xD(290)(3);
  VNStageIntLLRInputS1xD(297)(5) <= CNStageIntLLROutputS1xD(290)(4);
  VNStageIntLLRInputS1xD(337)(5) <= CNStageIntLLROutputS1xD(290)(5);
  VNStageIntLLRInputS1xD(21)(5) <= CNStageIntLLROutputS1xD(291)(0);
  VNStageIntLLRInputS1xD(121)(4) <= CNStageIntLLROutputS1xD(291)(1);
  VNStageIntLLRInputS1xD(189)(4) <= CNStageIntLLROutputS1xD(291)(2);
  VNStageIntLLRInputS1xD(232)(4) <= CNStageIntLLROutputS1xD(291)(3);
  VNStageIntLLRInputS1xD(272)(5) <= CNStageIntLLROutputS1xD(291)(4);
  VNStageIntLLRInputS1xD(335)(5) <= CNStageIntLLROutputS1xD(291)(5);
  VNStageIntLLRInputS1xD(20)(3) <= CNStageIntLLROutputS1xD(292)(0);
  VNStageIntLLRInputS1xD(124)(3) <= CNStageIntLLROutputS1xD(292)(1);
  VNStageIntLLRInputS1xD(167)(5) <= CNStageIntLLROutputS1xD(292)(2);
  VNStageIntLLRInputS1xD(207)(4) <= CNStageIntLLROutputS1xD(292)(3);
  VNStageIntLLRInputS1xD(270)(5) <= CNStageIntLLROutputS1xD(292)(4);
  VNStageIntLLRInputS1xD(360)(5) <= CNStageIntLLROutputS1xD(292)(5);
  VNStageIntLLRInputS1xD(18)(5) <= CNStageIntLLROutputS1xD(293)(0);
  VNStageIntLLRInputS1xD(77)(3) <= CNStageIntLLROutputS1xD(293)(1);
  VNStageIntLLRInputS1xD(140)(5) <= CNStageIntLLROutputS1xD(293)(2);
  VNStageIntLLRInputS1xD(230)(4) <= CNStageIntLLROutputS1xD(293)(3);
  VNStageIntLLRInputS1xD(303)(5) <= CNStageIntLLROutputS1xD(293)(4);
  VNStageIntLLRInputS1xD(348)(5) <= CNStageIntLLROutputS1xD(293)(5);
  VNStageIntLLRInputS1xD(17)(5) <= CNStageIntLLROutputS1xD(294)(0);
  VNStageIntLLRInputS1xD(75)(5) <= CNStageIntLLROutputS1xD(294)(1);
  VNStageIntLLRInputS1xD(165)(4) <= CNStageIntLLROutputS1xD(294)(2);
  VNStageIntLLRInputS1xD(238)(5) <= CNStageIntLLROutputS1xD(294)(3);
  VNStageIntLLRInputS1xD(283)(5) <= CNStageIntLLROutputS1xD(294)(4);
  VNStageIntLLRInputS1xD(342)(4) <= CNStageIntLLROutputS1xD(294)(5);
  VNStageIntLLRInputS1xD(16)(4) <= CNStageIntLLROutputS1xD(295)(0);
  VNStageIntLLRInputS1xD(100)(5) <= CNStageIntLLROutputS1xD(295)(1);
  VNStageIntLLRInputS1xD(173)(5) <= CNStageIntLLROutputS1xD(295)(2);
  VNStageIntLLRInputS1xD(218)(5) <= CNStageIntLLROutputS1xD(295)(3);
  VNStageIntLLRInputS1xD(277)(5) <= CNStageIntLLROutputS1xD(295)(4);
  VNStageIntLLRInputS1xD(320)(3) <= CNStageIntLLROutputS1xD(295)(5);
  VNStageIntLLRInputS1xD(15)(5) <= CNStageIntLLROutputS1xD(296)(0);
  VNStageIntLLRInputS1xD(108)(5) <= CNStageIntLLROutputS1xD(296)(1);
  VNStageIntLLRInputS1xD(153)(5) <= CNStageIntLLROutputS1xD(296)(2);
  VNStageIntLLRInputS1xD(212)(4) <= CNStageIntLLROutputS1xD(296)(3);
  VNStageIntLLRInputS1xD(256)(4) <= CNStageIntLLROutputS1xD(296)(4);
  VNStageIntLLRInputS1xD(341)(5) <= CNStageIntLLROutputS1xD(296)(5);
  VNStageIntLLRInputS1xD(14)(5) <= CNStageIntLLROutputS1xD(297)(0);
  VNStageIntLLRInputS1xD(88)(5) <= CNStageIntLLROutputS1xD(297)(1);
  VNStageIntLLRInputS1xD(147)(5) <= CNStageIntLLROutputS1xD(297)(2);
  VNStageIntLLRInputS1xD(192)(5) <= CNStageIntLLROutputS1xD(297)(3);
  VNStageIntLLRInputS1xD(276)(5) <= CNStageIntLLROutputS1xD(297)(4);
  VNStageIntLLRInputS1xD(346)(5) <= CNStageIntLLROutputS1xD(297)(5);
  VNStageIntLLRInputS1xD(13)(4) <= CNStageIntLLROutputS1xD(298)(0);
  VNStageIntLLRInputS1xD(82)(5) <= CNStageIntLLROutputS1xD(298)(1);
  VNStageIntLLRInputS1xD(128)(5) <= CNStageIntLLROutputS1xD(298)(2);
  VNStageIntLLRInputS1xD(211)(5) <= CNStageIntLLROutputS1xD(298)(3);
  VNStageIntLLRInputS1xD(281)(5) <= CNStageIntLLROutputS1xD(298)(4);
  VNStageIntLLRInputS1xD(365)(5) <= CNStageIntLLROutputS1xD(298)(5);
  VNStageIntLLRInputS1xD(12)(5) <= CNStageIntLLROutputS1xD(299)(0);
  VNStageIntLLRInputS1xD(64)(4) <= CNStageIntLLROutputS1xD(299)(1);
  VNStageIntLLRInputS1xD(146)(4) <= CNStageIntLLROutputS1xD(299)(2);
  VNStageIntLLRInputS1xD(216)(5) <= CNStageIntLLROutputS1xD(299)(3);
  VNStageIntLLRInputS1xD(300)(4) <= CNStageIntLLROutputS1xD(299)(4);
  VNStageIntLLRInputS1xD(356)(4) <= CNStageIntLLROutputS1xD(299)(5);
  VNStageIntLLRInputS1xD(9)(5) <= CNStageIntLLROutputS1xD(300)(0);
  VNStageIntLLRInputS1xD(105)(4) <= CNStageIntLLROutputS1xD(300)(1);
  VNStageIntLLRInputS1xD(161)(5) <= CNStageIntLLROutputS1xD(300)(2);
  VNStageIntLLRInputS1xD(200)(5) <= CNStageIntLLROutputS1xD(300)(3);
  VNStageIntLLRInputS1xD(266)(4) <= CNStageIntLLROutputS1xD(300)(4);
  VNStageIntLLRInputS1xD(355)(5) <= CNStageIntLLROutputS1xD(300)(5);
  VNStageIntLLRInputS1xD(7)(5) <= CNStageIntLLROutputS1xD(301)(0);
  VNStageIntLLRInputS1xD(70)(5) <= CNStageIntLLROutputS1xD(301)(1);
  VNStageIntLLRInputS1xD(136)(5) <= CNStageIntLLROutputS1xD(301)(2);
  VNStageIntLLRInputS1xD(225)(5) <= CNStageIntLLROutputS1xD(301)(3);
  VNStageIntLLRInputS1xD(311)(4) <= CNStageIntLLROutputS1xD(301)(4);
  VNStageIntLLRInputS1xD(372)(4) <= CNStageIntLLROutputS1xD(301)(5);
  VNStageIntLLRInputS1xD(6)(5) <= CNStageIntLLROutputS1xD(302)(0);
  VNStageIntLLRInputS1xD(71)(4) <= CNStageIntLLROutputS1xD(302)(1);
  VNStageIntLLRInputS1xD(160)(5) <= CNStageIntLLROutputS1xD(302)(2);
  VNStageIntLLRInputS1xD(246)(5) <= CNStageIntLLROutputS1xD(302)(3);
  VNStageIntLLRInputS1xD(307)(5) <= CNStageIntLLROutputS1xD(302)(4);
  VNStageIntLLRInputS1xD(324)(5) <= CNStageIntLLROutputS1xD(302)(5);
  VNStageIntLLRInputS1xD(5)(5) <= CNStageIntLLROutputS1xD(303)(0);
  VNStageIntLLRInputS1xD(95)(5) <= CNStageIntLLROutputS1xD(303)(1);
  VNStageIntLLRInputS1xD(181)(5) <= CNStageIntLLROutputS1xD(303)(2);
  VNStageIntLLRInputS1xD(242)(5) <= CNStageIntLLROutputS1xD(303)(3);
  VNStageIntLLRInputS1xD(259)(3) <= CNStageIntLLROutputS1xD(303)(4);
  VNStageIntLLRInputS1xD(350)(5) <= CNStageIntLLROutputS1xD(303)(5);
  VNStageIntLLRInputS1xD(4)(4) <= CNStageIntLLROutputS1xD(304)(0);
  VNStageIntLLRInputS1xD(116)(4) <= CNStageIntLLROutputS1xD(304)(1);
  VNStageIntLLRInputS1xD(177)(5) <= CNStageIntLLROutputS1xD(304)(2);
  VNStageIntLLRInputS1xD(194)(5) <= CNStageIntLLROutputS1xD(304)(3);
  VNStageIntLLRInputS1xD(285)(5) <= CNStageIntLLROutputS1xD(304)(4);
  VNStageIntLLRInputS1xD(326)(4) <= CNStageIntLLROutputS1xD(304)(5);
  VNStageIntLLRInputS1xD(3)(4) <= CNStageIntLLROutputS1xD(305)(0);
  VNStageIntLLRInputS1xD(112)(5) <= CNStageIntLLROutputS1xD(305)(1);
  VNStageIntLLRInputS1xD(129)(5) <= CNStageIntLLROutputS1xD(305)(2);
  VNStageIntLLRInputS1xD(220)(5) <= CNStageIntLLROutputS1xD(305)(3);
  VNStageIntLLRInputS1xD(261)(4) <= CNStageIntLLROutputS1xD(305)(4);
  VNStageIntLLRInputS1xD(358)(4) <= CNStageIntLLROutputS1xD(305)(5);
  VNStageIntLLRInputS1xD(2)(5) <= CNStageIntLLROutputS1xD(306)(0);
  VNStageIntLLRInputS1xD(127)(5) <= CNStageIntLLROutputS1xD(306)(1);
  VNStageIntLLRInputS1xD(155)(5) <= CNStageIntLLROutputS1xD(306)(2);
  VNStageIntLLRInputS1xD(196)(5) <= CNStageIntLLROutputS1xD(306)(3);
  VNStageIntLLRInputS1xD(293)(4) <= CNStageIntLLROutputS1xD(306)(4);
  VNStageIntLLRInputS1xD(374)(5) <= CNStageIntLLROutputS1xD(306)(5);
  VNStageIntLLRInputS1xD(1)(4) <= CNStageIntLLROutputS1xD(307)(0);
  VNStageIntLLRInputS1xD(90)(5) <= CNStageIntLLROutputS1xD(307)(1);
  VNStageIntLLRInputS1xD(131)(4) <= CNStageIntLLROutputS1xD(307)(2);
  VNStageIntLLRInputS1xD(228)(5) <= CNStageIntLLROutputS1xD(307)(3);
  VNStageIntLLRInputS1xD(309)(5) <= CNStageIntLLROutputS1xD(307)(4);
  VNStageIntLLRInputS1xD(344)(5) <= CNStageIntLLROutputS1xD(307)(5);
  VNStageIntLLRInputS1xD(62)(4) <= CNStageIntLLROutputS1xD(308)(0);
  VNStageIntLLRInputS1xD(98)(4) <= CNStageIntLLROutputS1xD(308)(1);
  VNStageIntLLRInputS1xD(179)(5) <= CNStageIntLLROutputS1xD(308)(2);
  VNStageIntLLRInputS1xD(214)(5) <= CNStageIntLLROutputS1xD(308)(3);
  VNStageIntLLRInputS1xD(288)(5) <= CNStageIntLLROutputS1xD(308)(4);
  VNStageIntLLRInputS1xD(366)(5) <= CNStageIntLLROutputS1xD(308)(5);
  VNStageIntLLRInputS1xD(61)(4) <= CNStageIntLLROutputS1xD(309)(0);
  VNStageIntLLRInputS1xD(114)(5) <= CNStageIntLLROutputS1xD(309)(1);
  VNStageIntLLRInputS1xD(149)(5) <= CNStageIntLLROutputS1xD(309)(2);
  VNStageIntLLRInputS1xD(223)(5) <= CNStageIntLLROutputS1xD(309)(3);
  VNStageIntLLRInputS1xD(301)(5) <= CNStageIntLLROutputS1xD(309)(4);
  VNStageIntLLRInputS1xD(345)(4) <= CNStageIntLLROutputS1xD(309)(5);
  VNStageIntLLRInputS1xD(60)(4) <= CNStageIntLLROutputS1xD(310)(0);
  VNStageIntLLRInputS1xD(84)(4) <= CNStageIntLLROutputS1xD(310)(1);
  VNStageIntLLRInputS1xD(158)(5) <= CNStageIntLLROutputS1xD(310)(2);
  VNStageIntLLRInputS1xD(236)(5) <= CNStageIntLLROutputS1xD(310)(3);
  VNStageIntLLRInputS1xD(280)(5) <= CNStageIntLLROutputS1xD(310)(4);
  VNStageIntLLRInputS1xD(373)(3) <= CNStageIntLLROutputS1xD(310)(5);
  VNStageIntLLRInputS1xD(59)(3) <= CNStageIntLLROutputS1xD(311)(0);
  VNStageIntLLRInputS1xD(93)(5) <= CNStageIntLLROutputS1xD(311)(1);
  VNStageIntLLRInputS1xD(171)(3) <= CNStageIntLLROutputS1xD(311)(2);
  VNStageIntLLRInputS1xD(215)(5) <= CNStageIntLLROutputS1xD(311)(3);
  VNStageIntLLRInputS1xD(308)(3) <= CNStageIntLLROutputS1xD(311)(4);
  VNStageIntLLRInputS1xD(375)(4) <= CNStageIntLLROutputS1xD(311)(5);
  VNStageIntLLRInputS1xD(58)(3) <= CNStageIntLLROutputS1xD(312)(0);
  VNStageIntLLRInputS1xD(106)(4) <= CNStageIntLLROutputS1xD(312)(1);
  VNStageIntLLRInputS1xD(150)(4) <= CNStageIntLLROutputS1xD(312)(2);
  VNStageIntLLRInputS1xD(243)(5) <= CNStageIntLLROutputS1xD(312)(3);
  VNStageIntLLRInputS1xD(310)(4) <= CNStageIntLLROutputS1xD(312)(4);
  VNStageIntLLRInputS1xD(357)(5) <= CNStageIntLLROutputS1xD(312)(5);
  VNStageIntLLRInputS1xD(57)(4) <= CNStageIntLLROutputS1xD(313)(0);
  VNStageIntLLRInputS1xD(85)(4) <= CNStageIntLLROutputS1xD(313)(1);
  VNStageIntLLRInputS1xD(178)(4) <= CNStageIntLLROutputS1xD(313)(2);
  VNStageIntLLRInputS1xD(245)(5) <= CNStageIntLLROutputS1xD(313)(3);
  VNStageIntLLRInputS1xD(292)(5) <= CNStageIntLLROutputS1xD(313)(4);
  VNStageIntLLRInputS1xD(364)(5) <= CNStageIntLLROutputS1xD(313)(5);
  VNStageIntLLRInputS1xD(56)(5) <= CNStageIntLLROutputS1xD(314)(0);
  VNStageIntLLRInputS1xD(113)(5) <= CNStageIntLLROutputS1xD(314)(1);
  VNStageIntLLRInputS1xD(180)(3) <= CNStageIntLLROutputS1xD(314)(2);
  VNStageIntLLRInputS1xD(227)(5) <= CNStageIntLLROutputS1xD(314)(3);
  VNStageIntLLRInputS1xD(299)(4) <= CNStageIntLLROutputS1xD(314)(4);
  VNStageIntLLRInputS1xD(328)(3) <= CNStageIntLLROutputS1xD(314)(5);
  VNStageIntLLRInputS1xD(55)(5) <= CNStageIntLLROutputS1xD(315)(0);
  VNStageIntLLRInputS1xD(115)(5) <= CNStageIntLLROutputS1xD(315)(1);
  VNStageIntLLRInputS1xD(162)(5) <= CNStageIntLLROutputS1xD(315)(2);
  VNStageIntLLRInputS1xD(234)(5) <= CNStageIntLLROutputS1xD(315)(3);
  VNStageIntLLRInputS1xD(263)(5) <= CNStageIntLLROutputS1xD(315)(4);
  VNStageIntLLRInputS1xD(379)(3) <= CNStageIntLLROutputS1xD(315)(5);
  VNStageIntLLRInputS1xD(54)(4) <= CNStageIntLLROutputS1xD(316)(0);
  VNStageIntLLRInputS1xD(97)(5) <= CNStageIntLLROutputS1xD(316)(1);
  VNStageIntLLRInputS1xD(169)(5) <= CNStageIntLLROutputS1xD(316)(2);
  VNStageIntLLRInputS1xD(198)(5) <= CNStageIntLLROutputS1xD(316)(3);
  VNStageIntLLRInputS1xD(314)(2) <= CNStageIntLLROutputS1xD(316)(4);
  VNStageIntLLRInputS1xD(322)(4) <= CNStageIntLLROutputS1xD(316)(5);
  VNStageIntLLRInputS1xD(53)(4) <= CNStageIntLLROutputS1xD(317)(0);
  VNStageIntLLRInputS1xD(104)(5) <= CNStageIntLLROutputS1xD(317)(1);
  VNStageIntLLRInputS1xD(133)(3) <= CNStageIntLLROutputS1xD(317)(2);
  VNStageIntLLRInputS1xD(249)(3) <= CNStageIntLLROutputS1xD(317)(3);
  VNStageIntLLRInputS1xD(257)(5) <= CNStageIntLLROutputS1xD(317)(4);
  VNStageIntLLRInputS1xD(380)(4) <= CNStageIntLLROutputS1xD(317)(5);
  VNStageIntLLRInputS1xD(52)(3) <= CNStageIntLLROutputS1xD(318)(0);
  VNStageIntLLRInputS1xD(68)(4) <= CNStageIntLLROutputS1xD(318)(1);
  VNStageIntLLRInputS1xD(184)(5) <= CNStageIntLLROutputS1xD(318)(2);
  VNStageIntLLRInputS1xD(255)(5) <= CNStageIntLLROutputS1xD(318)(3);
  VNStageIntLLRInputS1xD(315)(4) <= CNStageIntLLROutputS1xD(318)(4);
  VNStageIntLLRInputS1xD(327)(5) <= CNStageIntLLROutputS1xD(318)(5);
  VNStageIntLLRInputS1xD(51)(4) <= CNStageIntLLROutputS1xD(319)(0);
  VNStageIntLLRInputS1xD(119)(4) <= CNStageIntLLROutputS1xD(319)(1);
  VNStageIntLLRInputS1xD(190)(3) <= CNStageIntLLROutputS1xD(319)(2);
  VNStageIntLLRInputS1xD(250)(3) <= CNStageIntLLROutputS1xD(319)(3);
  VNStageIntLLRInputS1xD(262)(4) <= CNStageIntLLROutputS1xD(319)(4);
  VNStageIntLLRInputS1xD(349)(4) <= CNStageIntLLROutputS1xD(319)(5);
  VNStageIntLLRInputS1xD(50)(5) <= CNStageIntLLROutputS1xD(320)(0);
  VNStageIntLLRInputS1xD(125)(2) <= CNStageIntLLROutputS1xD(320)(1);
  VNStageIntLLRInputS1xD(185)(2) <= CNStageIntLLROutputS1xD(320)(2);
  VNStageIntLLRInputS1xD(197)(5) <= CNStageIntLLROutputS1xD(320)(3);
  VNStageIntLLRInputS1xD(284)(5) <= CNStageIntLLROutputS1xD(320)(4);
  VNStageIntLLRInputS1xD(367)(5) <= CNStageIntLLROutputS1xD(320)(5);
  VNStageIntLLRInputS1xD(49)(5) <= CNStageIntLLROutputS1xD(321)(0);
  VNStageIntLLRInputS1xD(120)(2) <= CNStageIntLLROutputS1xD(321)(1);
  VNStageIntLLRInputS1xD(132)(4) <= CNStageIntLLROutputS1xD(321)(2);
  VNStageIntLLRInputS1xD(219)(4) <= CNStageIntLLROutputS1xD(321)(3);
  VNStageIntLLRInputS1xD(302)(5) <= CNStageIntLLROutputS1xD(321)(4);
  VNStageIntLLRInputS1xD(352)(5) <= CNStageIntLLROutputS1xD(321)(5);
  VNStageIntLLRInputS1xD(48)(2) <= CNStageIntLLROutputS1xD(322)(0);
  VNStageIntLLRInputS1xD(67)(2) <= CNStageIntLLROutputS1xD(322)(1);
  VNStageIntLLRInputS1xD(154)(4) <= CNStageIntLLROutputS1xD(322)(2);
  VNStageIntLLRInputS1xD(237)(4) <= CNStageIntLLROutputS1xD(322)(3);
  VNStageIntLLRInputS1xD(287)(5) <= CNStageIntLLROutputS1xD(322)(4);
  VNStageIntLLRInputS1xD(339)(5) <= CNStageIntLLROutputS1xD(322)(5);
  VNStageIntLLRInputS1xD(46)(5) <= CNStageIntLLROutputS1xD(323)(0);
  VNStageIntLLRInputS1xD(107)(4) <= CNStageIntLLROutputS1xD(323)(1);
  VNStageIntLLRInputS1xD(157)(4) <= CNStageIntLLROutputS1xD(323)(2);
  VNStageIntLLRInputS1xD(209)(4) <= CNStageIntLLROutputS1xD(323)(3);
  VNStageIntLLRInputS1xD(305)(5) <= CNStageIntLLROutputS1xD(323)(4);
  VNStageIntLLRInputS1xD(382)(4) <= CNStageIntLLROutputS1xD(323)(5);
  VNStageIntLLRInputS1xD(45)(5) <= CNStageIntLLROutputS1xD(324)(0);
  VNStageIntLLRInputS1xD(92)(5) <= CNStageIntLLROutputS1xD(324)(1);
  VNStageIntLLRInputS1xD(144)(5) <= CNStageIntLLROutputS1xD(324)(2);
  VNStageIntLLRInputS1xD(240)(5) <= CNStageIntLLROutputS1xD(324)(3);
  VNStageIntLLRInputS1xD(317)(2) <= CNStageIntLLROutputS1xD(324)(4);
  VNStageIntLLRInputS1xD(333)(4) <= CNStageIntLLROutputS1xD(324)(5);
  VNStageIntLLRInputS1xD(44)(5) <= CNStageIntLLROutputS1xD(325)(0);
  VNStageIntLLRInputS1xD(79)(4) <= CNStageIntLLROutputS1xD(325)(1);
  VNStageIntLLRInputS1xD(175)(5) <= CNStageIntLLROutputS1xD(325)(2);
  VNStageIntLLRInputS1xD(252)(4) <= CNStageIntLLROutputS1xD(325)(3);
  VNStageIntLLRInputS1xD(268)(5) <= CNStageIntLLROutputS1xD(325)(4);
  VNStageIntLLRInputS1xD(377)(3) <= CNStageIntLLROutputS1xD(325)(5);
  VNStageIntLLRInputS1xD(43)(4) <= CNStageIntLLROutputS1xD(326)(0);
  VNStageIntLLRInputS1xD(110)(5) <= CNStageIntLLROutputS1xD(326)(1);
  VNStageIntLLRInputS1xD(187)(4) <= CNStageIntLLROutputS1xD(326)(2);
  VNStageIntLLRInputS1xD(203)(5) <= CNStageIntLLROutputS1xD(326)(3);
  VNStageIntLLRInputS1xD(312)(4) <= CNStageIntLLROutputS1xD(326)(4);
  VNStageIntLLRInputS1xD(354)(4) <= CNStageIntLLROutputS1xD(326)(5);
  VNStageIntLLRInputS1xD(42)(5) <= CNStageIntLLROutputS1xD(327)(0);
  VNStageIntLLRInputS1xD(122)(4) <= CNStageIntLLROutputS1xD(327)(1);
  VNStageIntLLRInputS1xD(138)(5) <= CNStageIntLLROutputS1xD(327)(2);
  VNStageIntLLRInputS1xD(247)(5) <= CNStageIntLLROutputS1xD(327)(3);
  VNStageIntLLRInputS1xD(289)(5) <= CNStageIntLLROutputS1xD(327)(4);
  VNStageIntLLRInputS1xD(343)(5) <= CNStageIntLLROutputS1xD(327)(5);
  VNStageIntLLRInputS1xD(41)(5) <= CNStageIntLLROutputS1xD(328)(0);
  VNStageIntLLRInputS1xD(73)(4) <= CNStageIntLLROutputS1xD(328)(1);
  VNStageIntLLRInputS1xD(182)(5) <= CNStageIntLLROutputS1xD(328)(2);
  VNStageIntLLRInputS1xD(224)(5) <= CNStageIntLLROutputS1xD(328)(3);
  VNStageIntLLRInputS1xD(278)(4) <= CNStageIntLLROutputS1xD(328)(4);
  VNStageIntLLRInputS1xD(347)(5) <= CNStageIntLLROutputS1xD(328)(5);
  VNStageIntLLRInputS1xD(39)(5) <= CNStageIntLLROutputS1xD(329)(0);
  VNStageIntLLRInputS1xD(94)(3) <= CNStageIntLLROutputS1xD(329)(1);
  VNStageIntLLRInputS1xD(148)(5) <= CNStageIntLLROutputS1xD(329)(2);
  VNStageIntLLRInputS1xD(217)(5) <= CNStageIntLLROutputS1xD(329)(3);
  VNStageIntLLRInputS1xD(275)(4) <= CNStageIntLLROutputS1xD(329)(4);
  VNStageIntLLRInputS1xD(351)(4) <= CNStageIntLLROutputS1xD(329)(5);
  VNStageIntLLRInputS1xD(38)(5) <= CNStageIntLLROutputS1xD(330)(0);
  VNStageIntLLRInputS1xD(83)(5) <= CNStageIntLLROutputS1xD(330)(1);
  VNStageIntLLRInputS1xD(152)(5) <= CNStageIntLLROutputS1xD(330)(2);
  VNStageIntLLRInputS1xD(210)(5) <= CNStageIntLLROutputS1xD(330)(3);
  VNStageIntLLRInputS1xD(286)(5) <= CNStageIntLLROutputS1xD(330)(4);
  VNStageIntLLRInputS1xD(323)(4) <= CNStageIntLLROutputS1xD(330)(5);
  VNStageIntLLRInputS1xD(37)(5) <= CNStageIntLLROutputS1xD(331)(0);
  VNStageIntLLRInputS1xD(87)(5) <= CNStageIntLLROutputS1xD(331)(1);
  VNStageIntLLRInputS1xD(145)(5) <= CNStageIntLLROutputS1xD(331)(2);
  VNStageIntLLRInputS1xD(221)(5) <= CNStageIntLLROutputS1xD(331)(3);
  VNStageIntLLRInputS1xD(258)(2) <= CNStageIntLLROutputS1xD(331)(4);
  VNStageIntLLRInputS1xD(378)(4) <= CNStageIntLLROutputS1xD(331)(5);
  VNStageIntLLRInputS1xD(0)(5) <= CNStageIntLLROutputS1xD(332)(0);
  VNStageIntLLRInputS1xD(76)(5) <= CNStageIntLLROutputS1xD(332)(1);
  VNStageIntLLRInputS1xD(141)(3) <= CNStageIntLLROutputS1xD(332)(2);
  VNStageIntLLRInputS1xD(206)(3) <= CNStageIntLLROutputS1xD(332)(3);
  VNStageIntLLRInputS1xD(271)(4) <= CNStageIntLLROutputS1xD(332)(4);
  VNStageIntLLRInputS1xD(336)(4) <= CNStageIntLLROutputS1xD(332)(5);
  VNStageIntLLRInputS1xD(28)(5) <= CNStageIntLLROutputS1xD(333)(0);
  VNStageIntLLRInputS1xD(106)(5) <= CNStageIntLLROutputS1xD(333)(1);
  VNStageIntLLRInputS1xD(144)(6) <= CNStageIntLLROutputS1xD(333)(2);
  VNStageIntLLRInputS1xD(193)(4) <= CNStageIntLLROutputS1xD(333)(3);
  VNStageIntLLRInputS1xD(261)(5) <= CNStageIntLLROutputS1xD(333)(4);
  VNStageIntLLRInputS1xD(367)(6) <= CNStageIntLLROutputS1xD(333)(5);
  VNStageIntLLRInputS1xD(26)(6) <= CNStageIntLLROutputS1xD(334)(0);
  VNStageIntLLRInputS1xD(126)(5) <= CNStageIntLLROutputS1xD(334)(1);
  VNStageIntLLRInputS1xD(131)(5) <= CNStageIntLLROutputS1xD(334)(2);
  VNStageIntLLRInputS1xD(237)(5) <= CNStageIntLLROutputS1xD(334)(3);
  VNStageIntLLRInputS1xD(277)(6) <= CNStageIntLLROutputS1xD(334)(4);
  VNStageIntLLRInputS1xD(340)(5) <= CNStageIntLLROutputS1xD(334)(5);
  VNStageIntLLRInputS1xD(24)(6) <= CNStageIntLLROutputS1xD(335)(0);
  VNStageIntLLRInputS1xD(107)(5) <= CNStageIntLLROutputS1xD(335)(1);
  VNStageIntLLRInputS1xD(147)(6) <= CNStageIntLLROutputS1xD(335)(2);
  VNStageIntLLRInputS1xD(210)(6) <= CNStageIntLLROutputS1xD(335)(3);
  VNStageIntLLRInputS1xD(300)(5) <= CNStageIntLLROutputS1xD(335)(4);
  VNStageIntLLRInputS1xD(373)(4) <= CNStageIntLLROutputS1xD(335)(5);
  VNStageIntLLRInputS1xD(23)(6) <= CNStageIntLLROutputS1xD(336)(0);
  VNStageIntLLRInputS1xD(82)(6) <= CNStageIntLLROutputS1xD(336)(1);
  VNStageIntLLRInputS1xD(145)(6) <= CNStageIntLLROutputS1xD(336)(2);
  VNStageIntLLRInputS1xD(235)(4) <= CNStageIntLLROutputS1xD(336)(3);
  VNStageIntLLRInputS1xD(308)(4) <= CNStageIntLLROutputS1xD(336)(4);
  VNStageIntLLRInputS1xD(353)(5) <= CNStageIntLLROutputS1xD(336)(5);
  VNStageIntLLRInputS1xD(22)(6) <= CNStageIntLLROutputS1xD(337)(0);
  VNStageIntLLRInputS1xD(80)(5) <= CNStageIntLLROutputS1xD(337)(1);
  VNStageIntLLRInputS1xD(170)(4) <= CNStageIntLLROutputS1xD(337)(2);
  VNStageIntLLRInputS1xD(243)(6) <= CNStageIntLLROutputS1xD(337)(3);
  VNStageIntLLRInputS1xD(288)(6) <= CNStageIntLLROutputS1xD(337)(4);
  VNStageIntLLRInputS1xD(347)(6) <= CNStageIntLLROutputS1xD(337)(5);
  VNStageIntLLRInputS1xD(21)(6) <= CNStageIntLLROutputS1xD(338)(0);
  VNStageIntLLRInputS1xD(105)(5) <= CNStageIntLLROutputS1xD(338)(1);
  VNStageIntLLRInputS1xD(178)(5) <= CNStageIntLLROutputS1xD(338)(2);
  VNStageIntLLRInputS1xD(223)(6) <= CNStageIntLLROutputS1xD(338)(3);
  VNStageIntLLRInputS1xD(282)(5) <= CNStageIntLLROutputS1xD(338)(4);
  VNStageIntLLRInputS1xD(320)(4) <= CNStageIntLLROutputS1xD(338)(5);
  VNStageIntLLRInputS1xD(20)(4) <= CNStageIntLLROutputS1xD(339)(0);
  VNStageIntLLRInputS1xD(113)(6) <= CNStageIntLLROutputS1xD(339)(1);
  VNStageIntLLRInputS1xD(158)(6) <= CNStageIntLLROutputS1xD(339)(2);
  VNStageIntLLRInputS1xD(217)(6) <= CNStageIntLLROutputS1xD(339)(3);
  VNStageIntLLRInputS1xD(256)(5) <= CNStageIntLLROutputS1xD(339)(4);
  VNStageIntLLRInputS1xD(346)(6) <= CNStageIntLLROutputS1xD(339)(5);
  VNStageIntLLRInputS1xD(19)(4) <= CNStageIntLLROutputS1xD(340)(0);
  VNStageIntLLRInputS1xD(93)(6) <= CNStageIntLLROutputS1xD(340)(1);
  VNStageIntLLRInputS1xD(152)(6) <= CNStageIntLLROutputS1xD(340)(2);
  VNStageIntLLRInputS1xD(192)(6) <= CNStageIntLLROutputS1xD(340)(3);
  VNStageIntLLRInputS1xD(281)(6) <= CNStageIntLLROutputS1xD(340)(4);
  VNStageIntLLRInputS1xD(351)(5) <= CNStageIntLLROutputS1xD(340)(5);
  VNStageIntLLRInputS1xD(18)(6) <= CNStageIntLLROutputS1xD(341)(0);
  VNStageIntLLRInputS1xD(87)(6) <= CNStageIntLLROutputS1xD(341)(1);
  VNStageIntLLRInputS1xD(128)(6) <= CNStageIntLLROutputS1xD(341)(2);
  VNStageIntLLRInputS1xD(216)(6) <= CNStageIntLLROutputS1xD(341)(3);
  VNStageIntLLRInputS1xD(286)(6) <= CNStageIntLLROutputS1xD(341)(4);
  VNStageIntLLRInputS1xD(370)(4) <= CNStageIntLLROutputS1xD(341)(5);
  VNStageIntLLRInputS1xD(17)(6) <= CNStageIntLLROutputS1xD(342)(0);
  VNStageIntLLRInputS1xD(64)(5) <= CNStageIntLLROutputS1xD(342)(1);
  VNStageIntLLRInputS1xD(151)(5) <= CNStageIntLLROutputS1xD(342)(2);
  VNStageIntLLRInputS1xD(221)(6) <= CNStageIntLLROutputS1xD(342)(3);
  VNStageIntLLRInputS1xD(305)(6) <= CNStageIntLLROutputS1xD(342)(4);
  VNStageIntLLRInputS1xD(361)(6) <= CNStageIntLLROutputS1xD(342)(5);
  VNStageIntLLRInputS1xD(16)(5) <= CNStageIntLLROutputS1xD(343)(0);
  VNStageIntLLRInputS1xD(86)(3) <= CNStageIntLLROutputS1xD(343)(1);
  VNStageIntLLRInputS1xD(156)(3) <= CNStageIntLLROutputS1xD(343)(2);
  VNStageIntLLRInputS1xD(240)(6) <= CNStageIntLLROutputS1xD(343)(3);
  VNStageIntLLRInputS1xD(296)(5) <= CNStageIntLLROutputS1xD(343)(4);
  VNStageIntLLRInputS1xD(335)(6) <= CNStageIntLLROutputS1xD(343)(5);
  VNStageIntLLRInputS1xD(15)(6) <= CNStageIntLLROutputS1xD(344)(0);
  VNStageIntLLRInputS1xD(91)(6) <= CNStageIntLLROutputS1xD(344)(1);
  VNStageIntLLRInputS1xD(175)(6) <= CNStageIntLLROutputS1xD(344)(2);
  VNStageIntLLRInputS1xD(231)(5) <= CNStageIntLLROutputS1xD(344)(3);
  VNStageIntLLRInputS1xD(270)(6) <= CNStageIntLLROutputS1xD(344)(4);
  VNStageIntLLRInputS1xD(336)(5) <= CNStageIntLLROutputS1xD(344)(5);
  VNStageIntLLRInputS1xD(14)(6) <= CNStageIntLLROutputS1xD(345)(0);
  VNStageIntLLRInputS1xD(110)(6) <= CNStageIntLLROutputS1xD(345)(1);
  VNStageIntLLRInputS1xD(166)(5) <= CNStageIntLLROutputS1xD(345)(2);
  VNStageIntLLRInputS1xD(205)(2) <= CNStageIntLLROutputS1xD(345)(3);
  VNStageIntLLRInputS1xD(271)(5) <= CNStageIntLLROutputS1xD(345)(4);
  VNStageIntLLRInputS1xD(360)(6) <= CNStageIntLLROutputS1xD(345)(5);
  VNStageIntLLRInputS1xD(13)(5) <= CNStageIntLLROutputS1xD(346)(0);
  VNStageIntLLRInputS1xD(101)(6) <= CNStageIntLLROutputS1xD(346)(1);
  VNStageIntLLRInputS1xD(140)(6) <= CNStageIntLLROutputS1xD(346)(2);
  VNStageIntLLRInputS1xD(206)(4) <= CNStageIntLLROutputS1xD(346)(3);
  VNStageIntLLRInputS1xD(295)(4) <= CNStageIntLLROutputS1xD(346)(4);
  VNStageIntLLRInputS1xD(381)(5) <= CNStageIntLLROutputS1xD(346)(5);
  VNStageIntLLRInputS1xD(12)(6) <= CNStageIntLLROutputS1xD(347)(0);
  VNStageIntLLRInputS1xD(75)(6) <= CNStageIntLLROutputS1xD(347)(1);
  VNStageIntLLRInputS1xD(141)(4) <= CNStageIntLLROutputS1xD(347)(2);
  VNStageIntLLRInputS1xD(230)(5) <= CNStageIntLLROutputS1xD(347)(3);
  VNStageIntLLRInputS1xD(316)(4) <= CNStageIntLLROutputS1xD(347)(4);
  VNStageIntLLRInputS1xD(377)(4) <= CNStageIntLLROutputS1xD(347)(5);
  VNStageIntLLRInputS1xD(11)(5) <= CNStageIntLLROutputS1xD(348)(0);
  VNStageIntLLRInputS1xD(76)(6) <= CNStageIntLLROutputS1xD(348)(1);
  VNStageIntLLRInputS1xD(165)(5) <= CNStageIntLLROutputS1xD(348)(2);
  VNStageIntLLRInputS1xD(251)(4) <= CNStageIntLLROutputS1xD(348)(3);
  VNStageIntLLRInputS1xD(312)(5) <= CNStageIntLLROutputS1xD(348)(4);
  VNStageIntLLRInputS1xD(329)(6) <= CNStageIntLLROutputS1xD(348)(5);
  VNStageIntLLRInputS1xD(10)(4) <= CNStageIntLLROutputS1xD(349)(0);
  VNStageIntLLRInputS1xD(100)(6) <= CNStageIntLLROutputS1xD(349)(1);
  VNStageIntLLRInputS1xD(186)(5) <= CNStageIntLLROutputS1xD(349)(2);
  VNStageIntLLRInputS1xD(247)(6) <= CNStageIntLLROutputS1xD(349)(3);
  VNStageIntLLRInputS1xD(264)(6) <= CNStageIntLLROutputS1xD(349)(4);
  VNStageIntLLRInputS1xD(355)(6) <= CNStageIntLLROutputS1xD(349)(5);
  VNStageIntLLRInputS1xD(9)(6) <= CNStageIntLLROutputS1xD(350)(0);
  VNStageIntLLRInputS1xD(121)(5) <= CNStageIntLLROutputS1xD(350)(1);
  VNStageIntLLRInputS1xD(182)(6) <= CNStageIntLLROutputS1xD(350)(2);
  VNStageIntLLRInputS1xD(199)(6) <= CNStageIntLLROutputS1xD(350)(3);
  VNStageIntLLRInputS1xD(290)(5) <= CNStageIntLLROutputS1xD(350)(4);
  VNStageIntLLRInputS1xD(331)(4) <= CNStageIntLLROutputS1xD(350)(5);
  VNStageIntLLRInputS1xD(7)(6) <= CNStageIntLLROutputS1xD(351)(0);
  VNStageIntLLRInputS1xD(69)(6) <= CNStageIntLLROutputS1xD(351)(1);
  VNStageIntLLRInputS1xD(160)(6) <= CNStageIntLLROutputS1xD(351)(2);
  VNStageIntLLRInputS1xD(201)(5) <= CNStageIntLLROutputS1xD(351)(3);
  VNStageIntLLRInputS1xD(298)(6) <= CNStageIntLLROutputS1xD(351)(4);
  VNStageIntLLRInputS1xD(379)(4) <= CNStageIntLLROutputS1xD(351)(5);
  VNStageIntLLRInputS1xD(6)(6) <= CNStageIntLLROutputS1xD(352)(0);
  VNStageIntLLRInputS1xD(95)(6) <= CNStageIntLLROutputS1xD(352)(1);
  VNStageIntLLRInputS1xD(136)(6) <= CNStageIntLLROutputS1xD(352)(2);
  VNStageIntLLRInputS1xD(233)(4) <= CNStageIntLLROutputS1xD(352)(3);
  VNStageIntLLRInputS1xD(314)(3) <= CNStageIntLLROutputS1xD(352)(4);
  VNStageIntLLRInputS1xD(349)(5) <= CNStageIntLLROutputS1xD(352)(5);
  VNStageIntLLRInputS1xD(5)(6) <= CNStageIntLLROutputS1xD(353)(0);
  VNStageIntLLRInputS1xD(71)(5) <= CNStageIntLLROutputS1xD(353)(1);
  VNStageIntLLRInputS1xD(168)(5) <= CNStageIntLLROutputS1xD(353)(2);
  VNStageIntLLRInputS1xD(249)(4) <= CNStageIntLLROutputS1xD(353)(3);
  VNStageIntLLRInputS1xD(284)(6) <= CNStageIntLLROutputS1xD(353)(4);
  VNStageIntLLRInputS1xD(358)(5) <= CNStageIntLLROutputS1xD(353)(5);
  VNStageIntLLRInputS1xD(4)(5) <= CNStageIntLLROutputS1xD(354)(0);
  VNStageIntLLRInputS1xD(103)(6) <= CNStageIntLLROutputS1xD(354)(1);
  VNStageIntLLRInputS1xD(184)(6) <= CNStageIntLLROutputS1xD(354)(2);
  VNStageIntLLRInputS1xD(219)(5) <= CNStageIntLLROutputS1xD(354)(3);
  VNStageIntLLRInputS1xD(293)(5) <= CNStageIntLLROutputS1xD(354)(4);
  VNStageIntLLRInputS1xD(371)(4) <= CNStageIntLLROutputS1xD(354)(5);
  VNStageIntLLRInputS1xD(2)(6) <= CNStageIntLLROutputS1xD(355)(0);
  VNStageIntLLRInputS1xD(89)(5) <= CNStageIntLLROutputS1xD(355)(1);
  VNStageIntLLRInputS1xD(163)(4) <= CNStageIntLLROutputS1xD(355)(2);
  VNStageIntLLRInputS1xD(241)(5) <= CNStageIntLLROutputS1xD(355)(3);
  VNStageIntLLRInputS1xD(285)(6) <= CNStageIntLLROutputS1xD(355)(4);
  VNStageIntLLRInputS1xD(378)(5) <= CNStageIntLLROutputS1xD(355)(5);
  VNStageIntLLRInputS1xD(1)(5) <= CNStageIntLLROutputS1xD(356)(0);
  VNStageIntLLRInputS1xD(98)(5) <= CNStageIntLLROutputS1xD(356)(1);
  VNStageIntLLRInputS1xD(176)(6) <= CNStageIntLLROutputS1xD(356)(2);
  VNStageIntLLRInputS1xD(220)(6) <= CNStageIntLLROutputS1xD(356)(3);
  VNStageIntLLRInputS1xD(313)(3) <= CNStageIntLLROutputS1xD(356)(4);
  VNStageIntLLRInputS1xD(380)(5) <= CNStageIntLLROutputS1xD(356)(5);
  VNStageIntLLRInputS1xD(63)(3) <= CNStageIntLLROutputS1xD(357)(0);
  VNStageIntLLRInputS1xD(111)(6) <= CNStageIntLLROutputS1xD(357)(1);
  VNStageIntLLRInputS1xD(155)(6) <= CNStageIntLLROutputS1xD(357)(2);
  VNStageIntLLRInputS1xD(248)(6) <= CNStageIntLLROutputS1xD(357)(3);
  VNStageIntLLRInputS1xD(315)(5) <= CNStageIntLLROutputS1xD(357)(4);
  VNStageIntLLRInputS1xD(362)(6) <= CNStageIntLLROutputS1xD(357)(5);
  VNStageIntLLRInputS1xD(62)(5) <= CNStageIntLLROutputS1xD(358)(0);
  VNStageIntLLRInputS1xD(90)(6) <= CNStageIntLLROutputS1xD(358)(1);
  VNStageIntLLRInputS1xD(183)(4) <= CNStageIntLLROutputS1xD(358)(2);
  VNStageIntLLRInputS1xD(250)(4) <= CNStageIntLLROutputS1xD(358)(3);
  VNStageIntLLRInputS1xD(297)(6) <= CNStageIntLLROutputS1xD(358)(4);
  VNStageIntLLRInputS1xD(369)(4) <= CNStageIntLLROutputS1xD(358)(5);
  VNStageIntLLRInputS1xD(61)(5) <= CNStageIntLLROutputS1xD(359)(0);
  VNStageIntLLRInputS1xD(118)(5) <= CNStageIntLLROutputS1xD(359)(1);
  VNStageIntLLRInputS1xD(185)(3) <= CNStageIntLLROutputS1xD(359)(2);
  VNStageIntLLRInputS1xD(232)(5) <= CNStageIntLLROutputS1xD(359)(3);
  VNStageIntLLRInputS1xD(304)(6) <= CNStageIntLLROutputS1xD(359)(4);
  VNStageIntLLRInputS1xD(333)(5) <= CNStageIntLLROutputS1xD(359)(5);
  VNStageIntLLRInputS1xD(60)(5) <= CNStageIntLLROutputS1xD(360)(0);
  VNStageIntLLRInputS1xD(120)(3) <= CNStageIntLLROutputS1xD(360)(1);
  VNStageIntLLRInputS1xD(167)(6) <= CNStageIntLLROutputS1xD(360)(2);
  VNStageIntLLRInputS1xD(239)(6) <= CNStageIntLLROutputS1xD(360)(3);
  VNStageIntLLRInputS1xD(268)(6) <= CNStageIntLLROutputS1xD(360)(4);
  VNStageIntLLRInputS1xD(321)(6) <= CNStageIntLLROutputS1xD(360)(5);
  VNStageIntLLRInputS1xD(59)(4) <= CNStageIntLLROutputS1xD(361)(0);
  VNStageIntLLRInputS1xD(102)(5) <= CNStageIntLLROutputS1xD(361)(1);
  VNStageIntLLRInputS1xD(174)(4) <= CNStageIntLLROutputS1xD(361)(2);
  VNStageIntLLRInputS1xD(203)(6) <= CNStageIntLLROutputS1xD(361)(3);
  VNStageIntLLRInputS1xD(319)(6) <= CNStageIntLLROutputS1xD(361)(4);
  VNStageIntLLRInputS1xD(327)(6) <= CNStageIntLLROutputS1xD(361)(5);
  VNStageIntLLRInputS1xD(58)(4) <= CNStageIntLLROutputS1xD(362)(0);
  VNStageIntLLRInputS1xD(109)(5) <= CNStageIntLLROutputS1xD(362)(1);
  VNStageIntLLRInputS1xD(138)(6) <= CNStageIntLLROutputS1xD(362)(2);
  VNStageIntLLRInputS1xD(254)(4) <= CNStageIntLLROutputS1xD(362)(3);
  VNStageIntLLRInputS1xD(262)(5) <= CNStageIntLLROutputS1xD(362)(4);
  VNStageIntLLRInputS1xD(322)(5) <= CNStageIntLLROutputS1xD(362)(5);
  VNStageIntLLRInputS1xD(57)(5) <= CNStageIntLLROutputS1xD(363)(0);
  VNStageIntLLRInputS1xD(73)(5) <= CNStageIntLLROutputS1xD(363)(1);
  VNStageIntLLRInputS1xD(189)(5) <= CNStageIntLLROutputS1xD(363)(2);
  VNStageIntLLRInputS1xD(197)(6) <= CNStageIntLLROutputS1xD(363)(3);
  VNStageIntLLRInputS1xD(257)(6) <= CNStageIntLLROutputS1xD(363)(4);
  VNStageIntLLRInputS1xD(332)(5) <= CNStageIntLLROutputS1xD(363)(5);
  VNStageIntLLRInputS1xD(56)(6) <= CNStageIntLLROutputS1xD(364)(0);
  VNStageIntLLRInputS1xD(124)(4) <= CNStageIntLLROutputS1xD(364)(1);
  VNStageIntLLRInputS1xD(132)(5) <= CNStageIntLLROutputS1xD(364)(2);
  VNStageIntLLRInputS1xD(255)(6) <= CNStageIntLLROutputS1xD(364)(3);
  VNStageIntLLRInputS1xD(267)(6) <= CNStageIntLLROutputS1xD(364)(4);
  VNStageIntLLRInputS1xD(354)(5) <= CNStageIntLLROutputS1xD(364)(5);
  VNStageIntLLRInputS1xD(55)(6) <= CNStageIntLLROutputS1xD(365)(0);
  VNStageIntLLRInputS1xD(67)(3) <= CNStageIntLLROutputS1xD(365)(1);
  VNStageIntLLRInputS1xD(190)(4) <= CNStageIntLLROutputS1xD(365)(2);
  VNStageIntLLRInputS1xD(202)(5) <= CNStageIntLLROutputS1xD(365)(3);
  VNStageIntLLRInputS1xD(289)(6) <= CNStageIntLLROutputS1xD(365)(4);
  VNStageIntLLRInputS1xD(372)(5) <= CNStageIntLLROutputS1xD(365)(5);
  VNStageIntLLRInputS1xD(54)(5) <= CNStageIntLLROutputS1xD(366)(0);
  VNStageIntLLRInputS1xD(125)(3) <= CNStageIntLLROutputS1xD(366)(1);
  VNStageIntLLRInputS1xD(137)(6) <= CNStageIntLLROutputS1xD(366)(2);
  VNStageIntLLRInputS1xD(224)(6) <= CNStageIntLLROutputS1xD(366)(3);
  VNStageIntLLRInputS1xD(307)(6) <= CNStageIntLLROutputS1xD(366)(4);
  VNStageIntLLRInputS1xD(357)(6) <= CNStageIntLLROutputS1xD(366)(5);
  VNStageIntLLRInputS1xD(53)(5) <= CNStageIntLLROutputS1xD(367)(0);
  VNStageIntLLRInputS1xD(72)(5) <= CNStageIntLLROutputS1xD(367)(1);
  VNStageIntLLRInputS1xD(159)(4) <= CNStageIntLLROutputS1xD(367)(2);
  VNStageIntLLRInputS1xD(242)(6) <= CNStageIntLLROutputS1xD(367)(3);
  VNStageIntLLRInputS1xD(292)(6) <= CNStageIntLLROutputS1xD(367)(4);
  VNStageIntLLRInputS1xD(344)(6) <= CNStageIntLLROutputS1xD(367)(5);
  VNStageIntLLRInputS1xD(52)(4) <= CNStageIntLLROutputS1xD(368)(0);
  VNStageIntLLRInputS1xD(94)(4) <= CNStageIntLLROutputS1xD(368)(1);
  VNStageIntLLRInputS1xD(177)(6) <= CNStageIntLLROutputS1xD(368)(2);
  VNStageIntLLRInputS1xD(227)(6) <= CNStageIntLLROutputS1xD(368)(3);
  VNStageIntLLRInputS1xD(279)(5) <= CNStageIntLLROutputS1xD(368)(4);
  VNStageIntLLRInputS1xD(375)(5) <= CNStageIntLLROutputS1xD(368)(5);
  VNStageIntLLRInputS1xD(51)(5) <= CNStageIntLLROutputS1xD(369)(0);
  VNStageIntLLRInputS1xD(112)(6) <= CNStageIntLLROutputS1xD(369)(1);
  VNStageIntLLRInputS1xD(162)(6) <= CNStageIntLLROutputS1xD(369)(2);
  VNStageIntLLRInputS1xD(214)(6) <= CNStageIntLLROutputS1xD(369)(3);
  VNStageIntLLRInputS1xD(310)(5) <= CNStageIntLLROutputS1xD(369)(4);
  VNStageIntLLRInputS1xD(324)(6) <= CNStageIntLLROutputS1xD(369)(5);
  VNStageIntLLRInputS1xD(50)(6) <= CNStageIntLLROutputS1xD(370)(0);
  VNStageIntLLRInputS1xD(97)(6) <= CNStageIntLLROutputS1xD(370)(1);
  VNStageIntLLRInputS1xD(149)(6) <= CNStageIntLLROutputS1xD(370)(2);
  VNStageIntLLRInputS1xD(245)(6) <= CNStageIntLLROutputS1xD(370)(3);
  VNStageIntLLRInputS1xD(259)(4) <= CNStageIntLLROutputS1xD(370)(4);
  VNStageIntLLRInputS1xD(338)(4) <= CNStageIntLLROutputS1xD(370)(5);
  VNStageIntLLRInputS1xD(49)(6) <= CNStageIntLLROutputS1xD(371)(0);
  VNStageIntLLRInputS1xD(84)(5) <= CNStageIntLLROutputS1xD(371)(1);
  VNStageIntLLRInputS1xD(180)(4) <= CNStageIntLLROutputS1xD(371)(2);
  VNStageIntLLRInputS1xD(194)(6) <= CNStageIntLLROutputS1xD(371)(3);
  VNStageIntLLRInputS1xD(273)(5) <= CNStageIntLLROutputS1xD(371)(4);
  VNStageIntLLRInputS1xD(382)(5) <= CNStageIntLLROutputS1xD(371)(5);
  VNStageIntLLRInputS1xD(48)(3) <= CNStageIntLLROutputS1xD(372)(0);
  VNStageIntLLRInputS1xD(115)(6) <= CNStageIntLLROutputS1xD(372)(1);
  VNStageIntLLRInputS1xD(129)(6) <= CNStageIntLLROutputS1xD(372)(2);
  VNStageIntLLRInputS1xD(208)(5) <= CNStageIntLLROutputS1xD(372)(3);
  VNStageIntLLRInputS1xD(317)(3) <= CNStageIntLLROutputS1xD(372)(4);
  VNStageIntLLRInputS1xD(359)(6) <= CNStageIntLLROutputS1xD(372)(5);
  VNStageIntLLRInputS1xD(47)(3) <= CNStageIntLLROutputS1xD(373)(0);
  VNStageIntLLRInputS1xD(127)(6) <= CNStageIntLLROutputS1xD(373)(1);
  VNStageIntLLRInputS1xD(143)(6) <= CNStageIntLLROutputS1xD(373)(2);
  VNStageIntLLRInputS1xD(252)(5) <= CNStageIntLLROutputS1xD(373)(3);
  VNStageIntLLRInputS1xD(294)(6) <= CNStageIntLLROutputS1xD(373)(4);
  VNStageIntLLRInputS1xD(348)(6) <= CNStageIntLLROutputS1xD(373)(5);
  VNStageIntLLRInputS1xD(46)(6) <= CNStageIntLLROutputS1xD(374)(0);
  VNStageIntLLRInputS1xD(78)(6) <= CNStageIntLLROutputS1xD(374)(1);
  VNStageIntLLRInputS1xD(187)(5) <= CNStageIntLLROutputS1xD(374)(2);
  VNStageIntLLRInputS1xD(229)(4) <= CNStageIntLLROutputS1xD(374)(3);
  VNStageIntLLRInputS1xD(283)(6) <= CNStageIntLLROutputS1xD(374)(4);
  VNStageIntLLRInputS1xD(352)(6) <= CNStageIntLLROutputS1xD(374)(5);
  VNStageIntLLRInputS1xD(45)(6) <= CNStageIntLLROutputS1xD(375)(0);
  VNStageIntLLRInputS1xD(122)(5) <= CNStageIntLLROutputS1xD(375)(1);
  VNStageIntLLRInputS1xD(164)(5) <= CNStageIntLLROutputS1xD(375)(2);
  VNStageIntLLRInputS1xD(218)(6) <= CNStageIntLLROutputS1xD(375)(3);
  VNStageIntLLRInputS1xD(287)(6) <= CNStageIntLLROutputS1xD(375)(4);
  VNStageIntLLRInputS1xD(345)(5) <= CNStageIntLLROutputS1xD(375)(5);
  VNStageIntLLRInputS1xD(44)(6) <= CNStageIntLLROutputS1xD(376)(0);
  VNStageIntLLRInputS1xD(99)(6) <= CNStageIntLLROutputS1xD(376)(1);
  VNStageIntLLRInputS1xD(153)(6) <= CNStageIntLLROutputS1xD(376)(2);
  VNStageIntLLRInputS1xD(222)(3) <= CNStageIntLLROutputS1xD(376)(3);
  VNStageIntLLRInputS1xD(280)(6) <= CNStageIntLLROutputS1xD(376)(4);
  VNStageIntLLRInputS1xD(356)(5) <= CNStageIntLLROutputS1xD(376)(5);
  VNStageIntLLRInputS1xD(43)(5) <= CNStageIntLLROutputS1xD(377)(0);
  VNStageIntLLRInputS1xD(88)(6) <= CNStageIntLLROutputS1xD(377)(1);
  VNStageIntLLRInputS1xD(157)(5) <= CNStageIntLLROutputS1xD(377)(2);
  VNStageIntLLRInputS1xD(215)(6) <= CNStageIntLLROutputS1xD(377)(3);
  VNStageIntLLRInputS1xD(291)(5) <= CNStageIntLLROutputS1xD(377)(4);
  VNStageIntLLRInputS1xD(328)(4) <= CNStageIntLLROutputS1xD(377)(5);
  VNStageIntLLRInputS1xD(42)(6) <= CNStageIntLLROutputS1xD(378)(0);
  VNStageIntLLRInputS1xD(92)(6) <= CNStageIntLLROutputS1xD(378)(1);
  VNStageIntLLRInputS1xD(150)(5) <= CNStageIntLLROutputS1xD(378)(2);
  VNStageIntLLRInputS1xD(226)(2) <= CNStageIntLLROutputS1xD(378)(3);
  VNStageIntLLRInputS1xD(263)(6) <= CNStageIntLLROutputS1xD(378)(4);
  VNStageIntLLRInputS1xD(383)(6) <= CNStageIntLLROutputS1xD(378)(5);
  VNStageIntLLRInputS1xD(41)(6) <= CNStageIntLLROutputS1xD(379)(0);
  VNStageIntLLRInputS1xD(85)(5) <= CNStageIntLLROutputS1xD(379)(1);
  VNStageIntLLRInputS1xD(161)(6) <= CNStageIntLLROutputS1xD(379)(2);
  VNStageIntLLRInputS1xD(198)(6) <= CNStageIntLLROutputS1xD(379)(3);
  VNStageIntLLRInputS1xD(318)(3) <= CNStageIntLLROutputS1xD(379)(4);
  VNStageIntLLRInputS1xD(337)(6) <= CNStageIntLLROutputS1xD(379)(5);
  VNStageIntLLRInputS1xD(40)(4) <= CNStageIntLLROutputS1xD(380)(0);
  VNStageIntLLRInputS1xD(96)(5) <= CNStageIntLLROutputS1xD(380)(1);
  VNStageIntLLRInputS1xD(133)(4) <= CNStageIntLLROutputS1xD(380)(2);
  VNStageIntLLRInputS1xD(253)(5) <= CNStageIntLLROutputS1xD(380)(3);
  VNStageIntLLRInputS1xD(272)(6) <= CNStageIntLLROutputS1xD(380)(4);
  VNStageIntLLRInputS1xD(334)(4) <= CNStageIntLLROutputS1xD(380)(5);
  VNStageIntLLRInputS1xD(39)(6) <= CNStageIntLLROutputS1xD(381)(0);
  VNStageIntLLRInputS1xD(68)(5) <= CNStageIntLLROutputS1xD(381)(1);
  VNStageIntLLRInputS1xD(188)(4) <= CNStageIntLLROutputS1xD(381)(2);
  VNStageIntLLRInputS1xD(207)(5) <= CNStageIntLLROutputS1xD(381)(3);
  VNStageIntLLRInputS1xD(269)(5) <= CNStageIntLLROutputS1xD(381)(4);
  VNStageIntLLRInputS1xD(368)(2) <= CNStageIntLLROutputS1xD(381)(5);
  VNStageIntLLRInputS1xD(38)(6) <= CNStageIntLLROutputS1xD(382)(0);
  VNStageIntLLRInputS1xD(123)(4) <= CNStageIntLLROutputS1xD(382)(1);
  VNStageIntLLRInputS1xD(142)(4) <= CNStageIntLLROutputS1xD(382)(2);
  VNStageIntLLRInputS1xD(204)(6) <= CNStageIntLLROutputS1xD(382)(3);
  VNStageIntLLRInputS1xD(303)(6) <= CNStageIntLLROutputS1xD(382)(4);
  VNStageIntLLRInputS1xD(325)(6) <= CNStageIntLLROutputS1xD(382)(5);
  VNStageIntLLRInputS1xD(37)(6) <= CNStageIntLLROutputS1xD(383)(0);
  VNStageIntLLRInputS1xD(77)(4) <= CNStageIntLLROutputS1xD(383)(1);
  VNStageIntLLRInputS1xD(139)(6) <= CNStageIntLLROutputS1xD(383)(2);
  VNStageIntLLRInputS1xD(238)(6) <= CNStageIntLLROutputS1xD(383)(3);
  VNStageIntLLRInputS1xD(260)(5) <= CNStageIntLLROutputS1xD(383)(4);
  VNStageIntLLRInputS1xD(374)(6) <= CNStageIntLLROutputS1xD(383)(5);

  -- Check Nodes (Iteration 2)
  CNStageIntLLRInputS2xD(53)(0) <= VNStageIntLLROutputS1xD(0)(0);
  CNStageIntLLRInputS2xD(110)(0) <= VNStageIntLLROutputS1xD(0)(1);
  CNStageIntLLRInputS2xD(170)(0) <= VNStageIntLLROutputS1xD(0)(2);
  CNStageIntLLRInputS2xD(224)(0) <= VNStageIntLLROutputS1xD(0)(3);
  CNStageIntLLRInputS2xD(279)(0) <= VNStageIntLLROutputS1xD(0)(4);
  CNStageIntLLRInputS2xD(332)(0) <= VNStageIntLLROutputS1xD(0)(5);
  CNStageIntLLRInputS2xD(51)(0) <= VNStageIntLLROutputS1xD(1)(0);
  CNStageIntLLRInputS2xD(139)(0) <= VNStageIntLLROutputS1xD(1)(1);
  CNStageIntLLRInputS2xD(223)(0) <= VNStageIntLLROutputS1xD(1)(2);
  CNStageIntLLRInputS2xD(241)(0) <= VNStageIntLLROutputS1xD(1)(3);
  CNStageIntLLRInputS2xD(307)(0) <= VNStageIntLLROutputS1xD(1)(4);
  CNStageIntLLRInputS2xD(356)(0) <= VNStageIntLLROutputS1xD(1)(5);
  CNStageIntLLRInputS2xD(50)(0) <= VNStageIntLLROutputS1xD(2)(0);
  CNStageIntLLRInputS2xD(92)(0) <= VNStageIntLLROutputS1xD(2)(1);
  CNStageIntLLRInputS2xD(138)(0) <= VNStageIntLLROutputS1xD(2)(2);
  CNStageIntLLRInputS2xD(222)(0) <= VNStageIntLLROutputS1xD(2)(3);
  CNStageIntLLRInputS2xD(240)(0) <= VNStageIntLLROutputS1xD(2)(4);
  CNStageIntLLRInputS2xD(306)(0) <= VNStageIntLLROutputS1xD(2)(5);
  CNStageIntLLRInputS2xD(355)(0) <= VNStageIntLLROutputS1xD(2)(6);
  CNStageIntLLRInputS2xD(91)(0) <= VNStageIntLLROutputS1xD(3)(0);
  CNStageIntLLRInputS2xD(137)(0) <= VNStageIntLLROutputS1xD(3)(1);
  CNStageIntLLRInputS2xD(221)(0) <= VNStageIntLLROutputS1xD(3)(2);
  CNStageIntLLRInputS2xD(239)(0) <= VNStageIntLLROutputS1xD(3)(3);
  CNStageIntLLRInputS2xD(305)(0) <= VNStageIntLLROutputS1xD(3)(4);
  CNStageIntLLRInputS2xD(49)(0) <= VNStageIntLLROutputS1xD(4)(0);
  CNStageIntLLRInputS2xD(90)(0) <= VNStageIntLLROutputS1xD(4)(1);
  CNStageIntLLRInputS2xD(220)(0) <= VNStageIntLLROutputS1xD(4)(2);
  CNStageIntLLRInputS2xD(238)(0) <= VNStageIntLLROutputS1xD(4)(3);
  CNStageIntLLRInputS2xD(304)(0) <= VNStageIntLLROutputS1xD(4)(4);
  CNStageIntLLRInputS2xD(354)(0) <= VNStageIntLLROutputS1xD(4)(5);
  CNStageIntLLRInputS2xD(48)(0) <= VNStageIntLLROutputS1xD(5)(0);
  CNStageIntLLRInputS2xD(89)(0) <= VNStageIntLLROutputS1xD(5)(1);
  CNStageIntLLRInputS2xD(136)(0) <= VNStageIntLLROutputS1xD(5)(2);
  CNStageIntLLRInputS2xD(219)(0) <= VNStageIntLLROutputS1xD(5)(3);
  CNStageIntLLRInputS2xD(237)(0) <= VNStageIntLLROutputS1xD(5)(4);
  CNStageIntLLRInputS2xD(303)(0) <= VNStageIntLLROutputS1xD(5)(5);
  CNStageIntLLRInputS2xD(353)(0) <= VNStageIntLLROutputS1xD(5)(6);
  CNStageIntLLRInputS2xD(47)(0) <= VNStageIntLLROutputS1xD(6)(0);
  CNStageIntLLRInputS2xD(88)(0) <= VNStageIntLLROutputS1xD(6)(1);
  CNStageIntLLRInputS2xD(135)(0) <= VNStageIntLLROutputS1xD(6)(2);
  CNStageIntLLRInputS2xD(218)(0) <= VNStageIntLLROutputS1xD(6)(3);
  CNStageIntLLRInputS2xD(236)(0) <= VNStageIntLLROutputS1xD(6)(4);
  CNStageIntLLRInputS2xD(302)(0) <= VNStageIntLLROutputS1xD(6)(5);
  CNStageIntLLRInputS2xD(352)(0) <= VNStageIntLLROutputS1xD(6)(6);
  CNStageIntLLRInputS2xD(46)(0) <= VNStageIntLLROutputS1xD(7)(0);
  CNStageIntLLRInputS2xD(87)(0) <= VNStageIntLLROutputS1xD(7)(1);
  CNStageIntLLRInputS2xD(134)(0) <= VNStageIntLLROutputS1xD(7)(2);
  CNStageIntLLRInputS2xD(217)(0) <= VNStageIntLLROutputS1xD(7)(3);
  CNStageIntLLRInputS2xD(235)(0) <= VNStageIntLLROutputS1xD(7)(4);
  CNStageIntLLRInputS2xD(301)(0) <= VNStageIntLLROutputS1xD(7)(5);
  CNStageIntLLRInputS2xD(351)(0) <= VNStageIntLLROutputS1xD(7)(6);
  CNStageIntLLRInputS2xD(45)(0) <= VNStageIntLLROutputS1xD(8)(0);
  CNStageIntLLRInputS2xD(133)(0) <= VNStageIntLLROutputS1xD(8)(1);
  CNStageIntLLRInputS2xD(216)(0) <= VNStageIntLLROutputS1xD(8)(2);
  CNStageIntLLRInputS2xD(44)(0) <= VNStageIntLLROutputS1xD(9)(0);
  CNStageIntLLRInputS2xD(86)(0) <= VNStageIntLLROutputS1xD(9)(1);
  CNStageIntLLRInputS2xD(132)(0) <= VNStageIntLLROutputS1xD(9)(2);
  CNStageIntLLRInputS2xD(215)(0) <= VNStageIntLLROutputS1xD(9)(3);
  CNStageIntLLRInputS2xD(234)(0) <= VNStageIntLLROutputS1xD(9)(4);
  CNStageIntLLRInputS2xD(300)(0) <= VNStageIntLLROutputS1xD(9)(5);
  CNStageIntLLRInputS2xD(350)(0) <= VNStageIntLLROutputS1xD(9)(6);
  CNStageIntLLRInputS2xD(43)(0) <= VNStageIntLLROutputS1xD(10)(0);
  CNStageIntLLRInputS2xD(85)(0) <= VNStageIntLLROutputS1xD(10)(1);
  CNStageIntLLRInputS2xD(131)(0) <= VNStageIntLLROutputS1xD(10)(2);
  CNStageIntLLRInputS2xD(233)(0) <= VNStageIntLLROutputS1xD(10)(3);
  CNStageIntLLRInputS2xD(349)(0) <= VNStageIntLLROutputS1xD(10)(4);
  CNStageIntLLRInputS2xD(42)(0) <= VNStageIntLLROutputS1xD(11)(0);
  CNStageIntLLRInputS2xD(84)(0) <= VNStageIntLLROutputS1xD(11)(1);
  CNStageIntLLRInputS2xD(130)(0) <= VNStageIntLLROutputS1xD(11)(2);
  CNStageIntLLRInputS2xD(214)(0) <= VNStageIntLLROutputS1xD(11)(3);
  CNStageIntLLRInputS2xD(232)(0) <= VNStageIntLLROutputS1xD(11)(4);
  CNStageIntLLRInputS2xD(348)(0) <= VNStageIntLLROutputS1xD(11)(5);
  CNStageIntLLRInputS2xD(41)(0) <= VNStageIntLLROutputS1xD(12)(0);
  CNStageIntLLRInputS2xD(83)(0) <= VNStageIntLLROutputS1xD(12)(1);
  CNStageIntLLRInputS2xD(129)(0) <= VNStageIntLLROutputS1xD(12)(2);
  CNStageIntLLRInputS2xD(213)(0) <= VNStageIntLLROutputS1xD(12)(3);
  CNStageIntLLRInputS2xD(231)(0) <= VNStageIntLLROutputS1xD(12)(4);
  CNStageIntLLRInputS2xD(299)(0) <= VNStageIntLLROutputS1xD(12)(5);
  CNStageIntLLRInputS2xD(347)(0) <= VNStageIntLLROutputS1xD(12)(6);
  CNStageIntLLRInputS2xD(82)(0) <= VNStageIntLLROutputS1xD(13)(0);
  CNStageIntLLRInputS2xD(128)(0) <= VNStageIntLLROutputS1xD(13)(1);
  CNStageIntLLRInputS2xD(212)(0) <= VNStageIntLLROutputS1xD(13)(2);
  CNStageIntLLRInputS2xD(230)(0) <= VNStageIntLLROutputS1xD(13)(3);
  CNStageIntLLRInputS2xD(298)(0) <= VNStageIntLLROutputS1xD(13)(4);
  CNStageIntLLRInputS2xD(346)(0) <= VNStageIntLLROutputS1xD(13)(5);
  CNStageIntLLRInputS2xD(40)(0) <= VNStageIntLLROutputS1xD(14)(0);
  CNStageIntLLRInputS2xD(81)(0) <= VNStageIntLLROutputS1xD(14)(1);
  CNStageIntLLRInputS2xD(127)(0) <= VNStageIntLLROutputS1xD(14)(2);
  CNStageIntLLRInputS2xD(211)(0) <= VNStageIntLLROutputS1xD(14)(3);
  CNStageIntLLRInputS2xD(229)(0) <= VNStageIntLLROutputS1xD(14)(4);
  CNStageIntLLRInputS2xD(297)(0) <= VNStageIntLLROutputS1xD(14)(5);
  CNStageIntLLRInputS2xD(345)(0) <= VNStageIntLLROutputS1xD(14)(6);
  CNStageIntLLRInputS2xD(39)(0) <= VNStageIntLLROutputS1xD(15)(0);
  CNStageIntLLRInputS2xD(80)(0) <= VNStageIntLLROutputS1xD(15)(1);
  CNStageIntLLRInputS2xD(126)(0) <= VNStageIntLLROutputS1xD(15)(2);
  CNStageIntLLRInputS2xD(210)(0) <= VNStageIntLLROutputS1xD(15)(3);
  CNStageIntLLRInputS2xD(228)(0) <= VNStageIntLLROutputS1xD(15)(4);
  CNStageIntLLRInputS2xD(296)(0) <= VNStageIntLLROutputS1xD(15)(5);
  CNStageIntLLRInputS2xD(344)(0) <= VNStageIntLLROutputS1xD(15)(6);
  CNStageIntLLRInputS2xD(38)(0) <= VNStageIntLLROutputS1xD(16)(0);
  CNStageIntLLRInputS2xD(125)(0) <= VNStageIntLLROutputS1xD(16)(1);
  CNStageIntLLRInputS2xD(209)(0) <= VNStageIntLLROutputS1xD(16)(2);
  CNStageIntLLRInputS2xD(227)(0) <= VNStageIntLLROutputS1xD(16)(3);
  CNStageIntLLRInputS2xD(295)(0) <= VNStageIntLLROutputS1xD(16)(4);
  CNStageIntLLRInputS2xD(343)(0) <= VNStageIntLLROutputS1xD(16)(5);
  CNStageIntLLRInputS2xD(37)(0) <= VNStageIntLLROutputS1xD(17)(0);
  CNStageIntLLRInputS2xD(79)(0) <= VNStageIntLLROutputS1xD(17)(1);
  CNStageIntLLRInputS2xD(124)(0) <= VNStageIntLLROutputS1xD(17)(2);
  CNStageIntLLRInputS2xD(208)(0) <= VNStageIntLLROutputS1xD(17)(3);
  CNStageIntLLRInputS2xD(226)(0) <= VNStageIntLLROutputS1xD(17)(4);
  CNStageIntLLRInputS2xD(294)(0) <= VNStageIntLLROutputS1xD(17)(5);
  CNStageIntLLRInputS2xD(342)(0) <= VNStageIntLLROutputS1xD(17)(6);
  CNStageIntLLRInputS2xD(36)(0) <= VNStageIntLLROutputS1xD(18)(0);
  CNStageIntLLRInputS2xD(78)(0) <= VNStageIntLLROutputS1xD(18)(1);
  CNStageIntLLRInputS2xD(123)(0) <= VNStageIntLLROutputS1xD(18)(2);
  CNStageIntLLRInputS2xD(207)(0) <= VNStageIntLLROutputS1xD(18)(3);
  CNStageIntLLRInputS2xD(225)(0) <= VNStageIntLLROutputS1xD(18)(4);
  CNStageIntLLRInputS2xD(293)(0) <= VNStageIntLLROutputS1xD(18)(5);
  CNStageIntLLRInputS2xD(341)(0) <= VNStageIntLLROutputS1xD(18)(6);
  CNStageIntLLRInputS2xD(35)(0) <= VNStageIntLLROutputS1xD(19)(0);
  CNStageIntLLRInputS2xD(77)(0) <= VNStageIntLLROutputS1xD(19)(1);
  CNStageIntLLRInputS2xD(122)(0) <= VNStageIntLLROutputS1xD(19)(2);
  CNStageIntLLRInputS2xD(278)(0) <= VNStageIntLLROutputS1xD(19)(3);
  CNStageIntLLRInputS2xD(340)(0) <= VNStageIntLLROutputS1xD(19)(4);
  CNStageIntLLRInputS2xD(34)(0) <= VNStageIntLLROutputS1xD(20)(0);
  CNStageIntLLRInputS2xD(76)(0) <= VNStageIntLLROutputS1xD(20)(1);
  CNStageIntLLRInputS2xD(277)(0) <= VNStageIntLLROutputS1xD(20)(2);
  CNStageIntLLRInputS2xD(292)(0) <= VNStageIntLLROutputS1xD(20)(3);
  CNStageIntLLRInputS2xD(339)(0) <= VNStageIntLLROutputS1xD(20)(4);
  CNStageIntLLRInputS2xD(33)(0) <= VNStageIntLLROutputS1xD(21)(0);
  CNStageIntLLRInputS2xD(75)(0) <= VNStageIntLLROutputS1xD(21)(1);
  CNStageIntLLRInputS2xD(121)(0) <= VNStageIntLLROutputS1xD(21)(2);
  CNStageIntLLRInputS2xD(206)(0) <= VNStageIntLLROutputS1xD(21)(3);
  CNStageIntLLRInputS2xD(276)(0) <= VNStageIntLLROutputS1xD(21)(4);
  CNStageIntLLRInputS2xD(291)(0) <= VNStageIntLLROutputS1xD(21)(5);
  CNStageIntLLRInputS2xD(338)(0) <= VNStageIntLLROutputS1xD(21)(6);
  CNStageIntLLRInputS2xD(32)(0) <= VNStageIntLLROutputS1xD(22)(0);
  CNStageIntLLRInputS2xD(74)(0) <= VNStageIntLLROutputS1xD(22)(1);
  CNStageIntLLRInputS2xD(120)(0) <= VNStageIntLLROutputS1xD(22)(2);
  CNStageIntLLRInputS2xD(205)(0) <= VNStageIntLLROutputS1xD(22)(3);
  CNStageIntLLRInputS2xD(275)(0) <= VNStageIntLLROutputS1xD(22)(4);
  CNStageIntLLRInputS2xD(290)(0) <= VNStageIntLLROutputS1xD(22)(5);
  CNStageIntLLRInputS2xD(337)(0) <= VNStageIntLLROutputS1xD(22)(6);
  CNStageIntLLRInputS2xD(31)(0) <= VNStageIntLLROutputS1xD(23)(0);
  CNStageIntLLRInputS2xD(73)(0) <= VNStageIntLLROutputS1xD(23)(1);
  CNStageIntLLRInputS2xD(119)(0) <= VNStageIntLLROutputS1xD(23)(2);
  CNStageIntLLRInputS2xD(204)(0) <= VNStageIntLLROutputS1xD(23)(3);
  CNStageIntLLRInputS2xD(274)(0) <= VNStageIntLLROutputS1xD(23)(4);
  CNStageIntLLRInputS2xD(289)(0) <= VNStageIntLLROutputS1xD(23)(5);
  CNStageIntLLRInputS2xD(336)(0) <= VNStageIntLLROutputS1xD(23)(6);
  CNStageIntLLRInputS2xD(30)(0) <= VNStageIntLLROutputS1xD(24)(0);
  CNStageIntLLRInputS2xD(72)(0) <= VNStageIntLLROutputS1xD(24)(1);
  CNStageIntLLRInputS2xD(118)(0) <= VNStageIntLLROutputS1xD(24)(2);
  CNStageIntLLRInputS2xD(203)(0) <= VNStageIntLLROutputS1xD(24)(3);
  CNStageIntLLRInputS2xD(273)(0) <= VNStageIntLLROutputS1xD(24)(4);
  CNStageIntLLRInputS2xD(288)(0) <= VNStageIntLLROutputS1xD(24)(5);
  CNStageIntLLRInputS2xD(335)(0) <= VNStageIntLLROutputS1xD(24)(6);
  CNStageIntLLRInputS2xD(29)(0) <= VNStageIntLLROutputS1xD(25)(0);
  CNStageIntLLRInputS2xD(71)(0) <= VNStageIntLLROutputS1xD(25)(1);
  CNStageIntLLRInputS2xD(117)(0) <= VNStageIntLLROutputS1xD(25)(2);
  CNStageIntLLRInputS2xD(202)(0) <= VNStageIntLLROutputS1xD(25)(3);
  CNStageIntLLRInputS2xD(287)(0) <= VNStageIntLLROutputS1xD(25)(4);
  CNStageIntLLRInputS2xD(28)(0) <= VNStageIntLLROutputS1xD(26)(0);
  CNStageIntLLRInputS2xD(70)(0) <= VNStageIntLLROutputS1xD(26)(1);
  CNStageIntLLRInputS2xD(116)(0) <= VNStageIntLLROutputS1xD(26)(2);
  CNStageIntLLRInputS2xD(201)(0) <= VNStageIntLLROutputS1xD(26)(3);
  CNStageIntLLRInputS2xD(272)(0) <= VNStageIntLLROutputS1xD(26)(4);
  CNStageIntLLRInputS2xD(286)(0) <= VNStageIntLLROutputS1xD(26)(5);
  CNStageIntLLRInputS2xD(334)(0) <= VNStageIntLLROutputS1xD(26)(6);
  CNStageIntLLRInputS2xD(27)(0) <= VNStageIntLLROutputS1xD(27)(0);
  CNStageIntLLRInputS2xD(69)(0) <= VNStageIntLLROutputS1xD(27)(1);
  CNStageIntLLRInputS2xD(115)(0) <= VNStageIntLLROutputS1xD(27)(2);
  CNStageIntLLRInputS2xD(200)(0) <= VNStageIntLLROutputS1xD(27)(3);
  CNStageIntLLRInputS2xD(285)(0) <= VNStageIntLLROutputS1xD(27)(4);
  CNStageIntLLRInputS2xD(26)(0) <= VNStageIntLLROutputS1xD(28)(0);
  CNStageIntLLRInputS2xD(68)(0) <= VNStageIntLLROutputS1xD(28)(1);
  CNStageIntLLRInputS2xD(114)(0) <= VNStageIntLLROutputS1xD(28)(2);
  CNStageIntLLRInputS2xD(199)(0) <= VNStageIntLLROutputS1xD(28)(3);
  CNStageIntLLRInputS2xD(271)(0) <= VNStageIntLLROutputS1xD(28)(4);
  CNStageIntLLRInputS2xD(333)(0) <= VNStageIntLLROutputS1xD(28)(5);
  CNStageIntLLRInputS2xD(25)(0) <= VNStageIntLLROutputS1xD(29)(0);
  CNStageIntLLRInputS2xD(67)(0) <= VNStageIntLLROutputS1xD(29)(1);
  CNStageIntLLRInputS2xD(113)(0) <= VNStageIntLLROutputS1xD(29)(2);
  CNStageIntLLRInputS2xD(270)(0) <= VNStageIntLLROutputS1xD(29)(3);
  CNStageIntLLRInputS2xD(24)(0) <= VNStageIntLLROutputS1xD(30)(0);
  CNStageIntLLRInputS2xD(66)(0) <= VNStageIntLLROutputS1xD(30)(1);
  CNStageIntLLRInputS2xD(112)(0) <= VNStageIntLLROutputS1xD(30)(2);
  CNStageIntLLRInputS2xD(198)(0) <= VNStageIntLLROutputS1xD(30)(3);
  CNStageIntLLRInputS2xD(269)(0) <= VNStageIntLLROutputS1xD(30)(4);
  CNStageIntLLRInputS2xD(284)(0) <= VNStageIntLLROutputS1xD(30)(5);
  CNStageIntLLRInputS2xD(23)(0) <= VNStageIntLLROutputS1xD(31)(0);
  CNStageIntLLRInputS2xD(65)(0) <= VNStageIntLLROutputS1xD(31)(1);
  CNStageIntLLRInputS2xD(197)(0) <= VNStageIntLLROutputS1xD(31)(2);
  CNStageIntLLRInputS2xD(283)(0) <= VNStageIntLLROutputS1xD(31)(3);
  CNStageIntLLRInputS2xD(22)(0) <= VNStageIntLLROutputS1xD(32)(0);
  CNStageIntLLRInputS2xD(64)(0) <= VNStageIntLLROutputS1xD(32)(1);
  CNStageIntLLRInputS2xD(111)(0) <= VNStageIntLLROutputS1xD(32)(2);
  CNStageIntLLRInputS2xD(268)(0) <= VNStageIntLLROutputS1xD(32)(3);
  CNStageIntLLRInputS2xD(21)(0) <= VNStageIntLLROutputS1xD(33)(0);
  CNStageIntLLRInputS2xD(63)(0) <= VNStageIntLLROutputS1xD(33)(1);
  CNStageIntLLRInputS2xD(169)(0) <= VNStageIntLLROutputS1xD(33)(2);
  CNStageIntLLRInputS2xD(196)(0) <= VNStageIntLLROutputS1xD(33)(3);
  CNStageIntLLRInputS2xD(267)(0) <= VNStageIntLLROutputS1xD(33)(4);
  CNStageIntLLRInputS2xD(282)(0) <= VNStageIntLLROutputS1xD(33)(5);
  CNStageIntLLRInputS2xD(20)(0) <= VNStageIntLLROutputS1xD(34)(0);
  CNStageIntLLRInputS2xD(62)(0) <= VNStageIntLLROutputS1xD(34)(1);
  CNStageIntLLRInputS2xD(168)(0) <= VNStageIntLLROutputS1xD(34)(2);
  CNStageIntLLRInputS2xD(195)(0) <= VNStageIntLLROutputS1xD(34)(3);
  CNStageIntLLRInputS2xD(266)(0) <= VNStageIntLLROutputS1xD(34)(4);
  CNStageIntLLRInputS2xD(281)(0) <= VNStageIntLLROutputS1xD(34)(5);
  CNStageIntLLRInputS2xD(19)(0) <= VNStageIntLLROutputS1xD(35)(0);
  CNStageIntLLRInputS2xD(61)(0) <= VNStageIntLLROutputS1xD(35)(1);
  CNStageIntLLRInputS2xD(167)(0) <= VNStageIntLLROutputS1xD(35)(2);
  CNStageIntLLRInputS2xD(194)(0) <= VNStageIntLLROutputS1xD(35)(3);
  CNStageIntLLRInputS2xD(265)(0) <= VNStageIntLLROutputS1xD(35)(4);
  CNStageIntLLRInputS2xD(280)(0) <= VNStageIntLLROutputS1xD(35)(5);
  CNStageIntLLRInputS2xD(18)(0) <= VNStageIntLLROutputS1xD(36)(0);
  CNStageIntLLRInputS2xD(60)(0) <= VNStageIntLLROutputS1xD(36)(1);
  CNStageIntLLRInputS2xD(166)(0) <= VNStageIntLLROutputS1xD(36)(2);
  CNStageIntLLRInputS2xD(264)(0) <= VNStageIntLLROutputS1xD(36)(3);
  CNStageIntLLRInputS2xD(17)(0) <= VNStageIntLLROutputS1xD(37)(0);
  CNStageIntLLRInputS2xD(59)(0) <= VNStageIntLLROutputS1xD(37)(1);
  CNStageIntLLRInputS2xD(165)(0) <= VNStageIntLLROutputS1xD(37)(2);
  CNStageIntLLRInputS2xD(193)(0) <= VNStageIntLLROutputS1xD(37)(3);
  CNStageIntLLRInputS2xD(263)(0) <= VNStageIntLLROutputS1xD(37)(4);
  CNStageIntLLRInputS2xD(331)(0) <= VNStageIntLLROutputS1xD(37)(5);
  CNStageIntLLRInputS2xD(383)(0) <= VNStageIntLLROutputS1xD(37)(6);
  CNStageIntLLRInputS2xD(16)(0) <= VNStageIntLLROutputS1xD(38)(0);
  CNStageIntLLRInputS2xD(58)(0) <= VNStageIntLLROutputS1xD(38)(1);
  CNStageIntLLRInputS2xD(164)(0) <= VNStageIntLLROutputS1xD(38)(2);
  CNStageIntLLRInputS2xD(192)(0) <= VNStageIntLLROutputS1xD(38)(3);
  CNStageIntLLRInputS2xD(262)(0) <= VNStageIntLLROutputS1xD(38)(4);
  CNStageIntLLRInputS2xD(330)(0) <= VNStageIntLLROutputS1xD(38)(5);
  CNStageIntLLRInputS2xD(382)(0) <= VNStageIntLLROutputS1xD(38)(6);
  CNStageIntLLRInputS2xD(15)(0) <= VNStageIntLLROutputS1xD(39)(0);
  CNStageIntLLRInputS2xD(57)(0) <= VNStageIntLLROutputS1xD(39)(1);
  CNStageIntLLRInputS2xD(163)(0) <= VNStageIntLLROutputS1xD(39)(2);
  CNStageIntLLRInputS2xD(191)(0) <= VNStageIntLLROutputS1xD(39)(3);
  CNStageIntLLRInputS2xD(261)(0) <= VNStageIntLLROutputS1xD(39)(4);
  CNStageIntLLRInputS2xD(329)(0) <= VNStageIntLLROutputS1xD(39)(5);
  CNStageIntLLRInputS2xD(381)(0) <= VNStageIntLLROutputS1xD(39)(6);
  CNStageIntLLRInputS2xD(14)(0) <= VNStageIntLLROutputS1xD(40)(0);
  CNStageIntLLRInputS2xD(56)(0) <= VNStageIntLLROutputS1xD(40)(1);
  CNStageIntLLRInputS2xD(162)(0) <= VNStageIntLLROutputS1xD(40)(2);
  CNStageIntLLRInputS2xD(260)(0) <= VNStageIntLLROutputS1xD(40)(3);
  CNStageIntLLRInputS2xD(380)(0) <= VNStageIntLLROutputS1xD(40)(4);
  CNStageIntLLRInputS2xD(13)(0) <= VNStageIntLLROutputS1xD(41)(0);
  CNStageIntLLRInputS2xD(55)(0) <= VNStageIntLLROutputS1xD(41)(1);
  CNStageIntLLRInputS2xD(161)(0) <= VNStageIntLLROutputS1xD(41)(2);
  CNStageIntLLRInputS2xD(190)(0) <= VNStageIntLLROutputS1xD(41)(3);
  CNStageIntLLRInputS2xD(259)(0) <= VNStageIntLLROutputS1xD(41)(4);
  CNStageIntLLRInputS2xD(328)(0) <= VNStageIntLLROutputS1xD(41)(5);
  CNStageIntLLRInputS2xD(379)(0) <= VNStageIntLLROutputS1xD(41)(6);
  CNStageIntLLRInputS2xD(12)(0) <= VNStageIntLLROutputS1xD(42)(0);
  CNStageIntLLRInputS2xD(54)(0) <= VNStageIntLLROutputS1xD(42)(1);
  CNStageIntLLRInputS2xD(160)(0) <= VNStageIntLLROutputS1xD(42)(2);
  CNStageIntLLRInputS2xD(189)(0) <= VNStageIntLLROutputS1xD(42)(3);
  CNStageIntLLRInputS2xD(258)(0) <= VNStageIntLLROutputS1xD(42)(4);
  CNStageIntLLRInputS2xD(327)(0) <= VNStageIntLLROutputS1xD(42)(5);
  CNStageIntLLRInputS2xD(378)(0) <= VNStageIntLLROutputS1xD(42)(6);
  CNStageIntLLRInputS2xD(109)(0) <= VNStageIntLLROutputS1xD(43)(0);
  CNStageIntLLRInputS2xD(159)(0) <= VNStageIntLLROutputS1xD(43)(1);
  CNStageIntLLRInputS2xD(188)(0) <= VNStageIntLLROutputS1xD(43)(2);
  CNStageIntLLRInputS2xD(257)(0) <= VNStageIntLLROutputS1xD(43)(3);
  CNStageIntLLRInputS2xD(326)(0) <= VNStageIntLLROutputS1xD(43)(4);
  CNStageIntLLRInputS2xD(377)(0) <= VNStageIntLLROutputS1xD(43)(5);
  CNStageIntLLRInputS2xD(11)(0) <= VNStageIntLLROutputS1xD(44)(0);
  CNStageIntLLRInputS2xD(108)(0) <= VNStageIntLLROutputS1xD(44)(1);
  CNStageIntLLRInputS2xD(158)(0) <= VNStageIntLLROutputS1xD(44)(2);
  CNStageIntLLRInputS2xD(187)(0) <= VNStageIntLLROutputS1xD(44)(3);
  CNStageIntLLRInputS2xD(256)(0) <= VNStageIntLLROutputS1xD(44)(4);
  CNStageIntLLRInputS2xD(325)(0) <= VNStageIntLLROutputS1xD(44)(5);
  CNStageIntLLRInputS2xD(376)(0) <= VNStageIntLLROutputS1xD(44)(6);
  CNStageIntLLRInputS2xD(10)(0) <= VNStageIntLLROutputS1xD(45)(0);
  CNStageIntLLRInputS2xD(107)(0) <= VNStageIntLLROutputS1xD(45)(1);
  CNStageIntLLRInputS2xD(157)(0) <= VNStageIntLLROutputS1xD(45)(2);
  CNStageIntLLRInputS2xD(186)(0) <= VNStageIntLLROutputS1xD(45)(3);
  CNStageIntLLRInputS2xD(255)(0) <= VNStageIntLLROutputS1xD(45)(4);
  CNStageIntLLRInputS2xD(324)(0) <= VNStageIntLLROutputS1xD(45)(5);
  CNStageIntLLRInputS2xD(375)(0) <= VNStageIntLLROutputS1xD(45)(6);
  CNStageIntLLRInputS2xD(9)(0) <= VNStageIntLLROutputS1xD(46)(0);
  CNStageIntLLRInputS2xD(106)(0) <= VNStageIntLLROutputS1xD(46)(1);
  CNStageIntLLRInputS2xD(156)(0) <= VNStageIntLLROutputS1xD(46)(2);
  CNStageIntLLRInputS2xD(185)(0) <= VNStageIntLLROutputS1xD(46)(3);
  CNStageIntLLRInputS2xD(254)(0) <= VNStageIntLLROutputS1xD(46)(4);
  CNStageIntLLRInputS2xD(323)(0) <= VNStageIntLLROutputS1xD(46)(5);
  CNStageIntLLRInputS2xD(374)(0) <= VNStageIntLLROutputS1xD(46)(6);
  CNStageIntLLRInputS2xD(8)(0) <= VNStageIntLLROutputS1xD(47)(0);
  CNStageIntLLRInputS2xD(155)(0) <= VNStageIntLLROutputS1xD(47)(1);
  CNStageIntLLRInputS2xD(253)(0) <= VNStageIntLLROutputS1xD(47)(2);
  CNStageIntLLRInputS2xD(373)(0) <= VNStageIntLLROutputS1xD(47)(3);
  CNStageIntLLRInputS2xD(7)(0) <= VNStageIntLLROutputS1xD(48)(0);
  CNStageIntLLRInputS2xD(154)(0) <= VNStageIntLLROutputS1xD(48)(1);
  CNStageIntLLRInputS2xD(322)(0) <= VNStageIntLLROutputS1xD(48)(2);
  CNStageIntLLRInputS2xD(372)(0) <= VNStageIntLLROutputS1xD(48)(3);
  CNStageIntLLRInputS2xD(6)(0) <= VNStageIntLLROutputS1xD(49)(0);
  CNStageIntLLRInputS2xD(105)(0) <= VNStageIntLLROutputS1xD(49)(1);
  CNStageIntLLRInputS2xD(153)(0) <= VNStageIntLLROutputS1xD(49)(2);
  CNStageIntLLRInputS2xD(184)(0) <= VNStageIntLLROutputS1xD(49)(3);
  CNStageIntLLRInputS2xD(252)(0) <= VNStageIntLLROutputS1xD(49)(4);
  CNStageIntLLRInputS2xD(321)(0) <= VNStageIntLLROutputS1xD(49)(5);
  CNStageIntLLRInputS2xD(371)(0) <= VNStageIntLLROutputS1xD(49)(6);
  CNStageIntLLRInputS2xD(5)(0) <= VNStageIntLLROutputS1xD(50)(0);
  CNStageIntLLRInputS2xD(104)(0) <= VNStageIntLLROutputS1xD(50)(1);
  CNStageIntLLRInputS2xD(152)(0) <= VNStageIntLLROutputS1xD(50)(2);
  CNStageIntLLRInputS2xD(183)(0) <= VNStageIntLLROutputS1xD(50)(3);
  CNStageIntLLRInputS2xD(251)(0) <= VNStageIntLLROutputS1xD(50)(4);
  CNStageIntLLRInputS2xD(320)(0) <= VNStageIntLLROutputS1xD(50)(5);
  CNStageIntLLRInputS2xD(370)(0) <= VNStageIntLLROutputS1xD(50)(6);
  CNStageIntLLRInputS2xD(4)(0) <= VNStageIntLLROutputS1xD(51)(0);
  CNStageIntLLRInputS2xD(103)(0) <= VNStageIntLLROutputS1xD(51)(1);
  CNStageIntLLRInputS2xD(182)(0) <= VNStageIntLLROutputS1xD(51)(2);
  CNStageIntLLRInputS2xD(250)(0) <= VNStageIntLLROutputS1xD(51)(3);
  CNStageIntLLRInputS2xD(319)(0) <= VNStageIntLLROutputS1xD(51)(4);
  CNStageIntLLRInputS2xD(369)(0) <= VNStageIntLLROutputS1xD(51)(5);
  CNStageIntLLRInputS2xD(102)(0) <= VNStageIntLLROutputS1xD(52)(0);
  CNStageIntLLRInputS2xD(151)(0) <= VNStageIntLLROutputS1xD(52)(1);
  CNStageIntLLRInputS2xD(181)(0) <= VNStageIntLLROutputS1xD(52)(2);
  CNStageIntLLRInputS2xD(318)(0) <= VNStageIntLLROutputS1xD(52)(3);
  CNStageIntLLRInputS2xD(368)(0) <= VNStageIntLLROutputS1xD(52)(4);
  CNStageIntLLRInputS2xD(3)(0) <= VNStageIntLLROutputS1xD(53)(0);
  CNStageIntLLRInputS2xD(150)(0) <= VNStageIntLLROutputS1xD(53)(1);
  CNStageIntLLRInputS2xD(180)(0) <= VNStageIntLLROutputS1xD(53)(2);
  CNStageIntLLRInputS2xD(249)(0) <= VNStageIntLLROutputS1xD(53)(3);
  CNStageIntLLRInputS2xD(317)(0) <= VNStageIntLLROutputS1xD(53)(4);
  CNStageIntLLRInputS2xD(367)(0) <= VNStageIntLLROutputS1xD(53)(5);
  CNStageIntLLRInputS2xD(2)(0) <= VNStageIntLLROutputS1xD(54)(0);
  CNStageIntLLRInputS2xD(101)(0) <= VNStageIntLLROutputS1xD(54)(1);
  CNStageIntLLRInputS2xD(149)(0) <= VNStageIntLLROutputS1xD(54)(2);
  CNStageIntLLRInputS2xD(179)(0) <= VNStageIntLLROutputS1xD(54)(3);
  CNStageIntLLRInputS2xD(316)(0) <= VNStageIntLLROutputS1xD(54)(4);
  CNStageIntLLRInputS2xD(366)(0) <= VNStageIntLLROutputS1xD(54)(5);
  CNStageIntLLRInputS2xD(1)(0) <= VNStageIntLLROutputS1xD(55)(0);
  CNStageIntLLRInputS2xD(100)(0) <= VNStageIntLLROutputS1xD(55)(1);
  CNStageIntLLRInputS2xD(148)(0) <= VNStageIntLLROutputS1xD(55)(2);
  CNStageIntLLRInputS2xD(178)(0) <= VNStageIntLLROutputS1xD(55)(3);
  CNStageIntLLRInputS2xD(248)(0) <= VNStageIntLLROutputS1xD(55)(4);
  CNStageIntLLRInputS2xD(315)(0) <= VNStageIntLLROutputS1xD(55)(5);
  CNStageIntLLRInputS2xD(365)(0) <= VNStageIntLLROutputS1xD(55)(6);
  CNStageIntLLRInputS2xD(0)(0) <= VNStageIntLLROutputS1xD(56)(0);
  CNStageIntLLRInputS2xD(99)(0) <= VNStageIntLLROutputS1xD(56)(1);
  CNStageIntLLRInputS2xD(147)(0) <= VNStageIntLLROutputS1xD(56)(2);
  CNStageIntLLRInputS2xD(177)(0) <= VNStageIntLLROutputS1xD(56)(3);
  CNStageIntLLRInputS2xD(247)(0) <= VNStageIntLLROutputS1xD(56)(4);
  CNStageIntLLRInputS2xD(314)(0) <= VNStageIntLLROutputS1xD(56)(5);
  CNStageIntLLRInputS2xD(364)(0) <= VNStageIntLLROutputS1xD(56)(6);
  CNStageIntLLRInputS2xD(98)(0) <= VNStageIntLLROutputS1xD(57)(0);
  CNStageIntLLRInputS2xD(146)(0) <= VNStageIntLLROutputS1xD(57)(1);
  CNStageIntLLRInputS2xD(176)(0) <= VNStageIntLLROutputS1xD(57)(2);
  CNStageIntLLRInputS2xD(246)(0) <= VNStageIntLLROutputS1xD(57)(3);
  CNStageIntLLRInputS2xD(313)(0) <= VNStageIntLLROutputS1xD(57)(4);
  CNStageIntLLRInputS2xD(363)(0) <= VNStageIntLLROutputS1xD(57)(5);
  CNStageIntLLRInputS2xD(97)(0) <= VNStageIntLLROutputS1xD(58)(0);
  CNStageIntLLRInputS2xD(145)(0) <= VNStageIntLLROutputS1xD(58)(1);
  CNStageIntLLRInputS2xD(175)(0) <= VNStageIntLLROutputS1xD(58)(2);
  CNStageIntLLRInputS2xD(312)(0) <= VNStageIntLLROutputS1xD(58)(3);
  CNStageIntLLRInputS2xD(362)(0) <= VNStageIntLLROutputS1xD(58)(4);
  CNStageIntLLRInputS2xD(144)(0) <= VNStageIntLLROutputS1xD(59)(0);
  CNStageIntLLRInputS2xD(174)(0) <= VNStageIntLLROutputS1xD(59)(1);
  CNStageIntLLRInputS2xD(245)(0) <= VNStageIntLLROutputS1xD(59)(2);
  CNStageIntLLRInputS2xD(311)(0) <= VNStageIntLLROutputS1xD(59)(3);
  CNStageIntLLRInputS2xD(361)(0) <= VNStageIntLLROutputS1xD(59)(4);
  CNStageIntLLRInputS2xD(96)(0) <= VNStageIntLLROutputS1xD(60)(0);
  CNStageIntLLRInputS2xD(143)(0) <= VNStageIntLLROutputS1xD(60)(1);
  CNStageIntLLRInputS2xD(173)(0) <= VNStageIntLLROutputS1xD(60)(2);
  CNStageIntLLRInputS2xD(244)(0) <= VNStageIntLLROutputS1xD(60)(3);
  CNStageIntLLRInputS2xD(310)(0) <= VNStageIntLLROutputS1xD(60)(4);
  CNStageIntLLRInputS2xD(360)(0) <= VNStageIntLLROutputS1xD(60)(5);
  CNStageIntLLRInputS2xD(95)(0) <= VNStageIntLLROutputS1xD(61)(0);
  CNStageIntLLRInputS2xD(142)(0) <= VNStageIntLLROutputS1xD(61)(1);
  CNStageIntLLRInputS2xD(172)(0) <= VNStageIntLLROutputS1xD(61)(2);
  CNStageIntLLRInputS2xD(243)(0) <= VNStageIntLLROutputS1xD(61)(3);
  CNStageIntLLRInputS2xD(309)(0) <= VNStageIntLLROutputS1xD(61)(4);
  CNStageIntLLRInputS2xD(359)(0) <= VNStageIntLLROutputS1xD(61)(5);
  CNStageIntLLRInputS2xD(94)(0) <= VNStageIntLLROutputS1xD(62)(0);
  CNStageIntLLRInputS2xD(141)(0) <= VNStageIntLLROutputS1xD(62)(1);
  CNStageIntLLRInputS2xD(171)(0) <= VNStageIntLLROutputS1xD(62)(2);
  CNStageIntLLRInputS2xD(242)(0) <= VNStageIntLLROutputS1xD(62)(3);
  CNStageIntLLRInputS2xD(308)(0) <= VNStageIntLLROutputS1xD(62)(4);
  CNStageIntLLRInputS2xD(358)(0) <= VNStageIntLLROutputS1xD(62)(5);
  CNStageIntLLRInputS2xD(52)(0) <= VNStageIntLLROutputS1xD(63)(0);
  CNStageIntLLRInputS2xD(93)(0) <= VNStageIntLLROutputS1xD(63)(1);
  CNStageIntLLRInputS2xD(140)(0) <= VNStageIntLLROutputS1xD(63)(2);
  CNStageIntLLRInputS2xD(357)(0) <= VNStageIntLLROutputS1xD(63)(3);
  CNStageIntLLRInputS2xD(53)(1) <= VNStageIntLLROutputS1xD(64)(0);
  CNStageIntLLRInputS2xD(109)(1) <= VNStageIntLLROutputS1xD(64)(1);
  CNStageIntLLRInputS2xD(130)(1) <= VNStageIntLLROutputS1xD(64)(2);
  CNStageIntLLRInputS2xD(245)(1) <= VNStageIntLLROutputS1xD(64)(3);
  CNStageIntLLRInputS2xD(299)(1) <= VNStageIntLLROutputS1xD(64)(4);
  CNStageIntLLRInputS2xD(342)(1) <= VNStageIntLLROutputS1xD(64)(5);
  CNStageIntLLRInputS2xD(51)(1) <= VNStageIntLLROutputS1xD(65)(0);
  CNStageIntLLRInputS2xD(74)(1) <= VNStageIntLLROutputS1xD(65)(1);
  CNStageIntLLRInputS2xD(141)(1) <= VNStageIntLLROutputS1xD(65)(2);
  CNStageIntLLRInputS2xD(189)(1) <= VNStageIntLLROutputS1xD(65)(3);
  CNStageIntLLRInputS2xD(286)(1) <= VNStageIntLLROutputS1xD(65)(4);
  CNStageIntLLRInputS2xD(50)(1) <= VNStageIntLLROutputS1xD(66)(0);
  CNStageIntLLRInputS2xD(66)(1) <= VNStageIntLLROutputS1xD(66)(1);
  CNStageIntLLRInputS2xD(155)(1) <= VNStageIntLLROutputS1xD(66)(2);
  CNStageIntLLRInputS2xD(244)(1) <= VNStageIntLLROutputS1xD(66)(3);
  CNStageIntLLRInputS2xD(97)(1) <= VNStageIntLLROutputS1xD(67)(0);
  CNStageIntLLRInputS2xD(275)(1) <= VNStageIntLLROutputS1xD(67)(1);
  CNStageIntLLRInputS2xD(322)(1) <= VNStageIntLLROutputS1xD(67)(2);
  CNStageIntLLRInputS2xD(365)(1) <= VNStageIntLLROutputS1xD(67)(3);
  CNStageIntLLRInputS2xD(49)(1) <= VNStageIntLLROutputS1xD(68)(0);
  CNStageIntLLRInputS2xD(112)(1) <= VNStageIntLLROutputS1xD(68)(1);
  CNStageIntLLRInputS2xD(210)(1) <= VNStageIntLLROutputS1xD(68)(2);
  CNStageIntLLRInputS2xD(256)(1) <= VNStageIntLLROutputS1xD(68)(3);
  CNStageIntLLRInputS2xD(318)(1) <= VNStageIntLLROutputS1xD(68)(4);
  CNStageIntLLRInputS2xD(381)(1) <= VNStageIntLLROutputS1xD(68)(5);
  CNStageIntLLRInputS2xD(48)(1) <= VNStageIntLLROutputS1xD(69)(0);
  CNStageIntLLRInputS2xD(101)(1) <= VNStageIntLLROutputS1xD(69)(1);
  CNStageIntLLRInputS2xD(135)(1) <= VNStageIntLLROutputS1xD(69)(2);
  CNStageIntLLRInputS2xD(215)(1) <= VNStageIntLLROutputS1xD(69)(3);
  CNStageIntLLRInputS2xD(259)(1) <= VNStageIntLLROutputS1xD(69)(4);
  CNStageIntLLRInputS2xD(283)(1) <= VNStageIntLLROutputS1xD(69)(5);
  CNStageIntLLRInputS2xD(351)(1) <= VNStageIntLLROutputS1xD(69)(6);
  CNStageIntLLRInputS2xD(47)(1) <= VNStageIntLLROutputS1xD(70)(0);
  CNStageIntLLRInputS2xD(104)(1) <= VNStageIntLLROutputS1xD(70)(1);
  CNStageIntLLRInputS2xD(136)(1) <= VNStageIntLLROutputS1xD(70)(2);
  CNStageIntLLRInputS2xD(206)(1) <= VNStageIntLLROutputS1xD(70)(3);
  CNStageIntLLRInputS2xD(246)(1) <= VNStageIntLLROutputS1xD(70)(4);
  CNStageIntLLRInputS2xD(301)(1) <= VNStageIntLLROutputS1xD(70)(5);
  CNStageIntLLRInputS2xD(46)(1) <= VNStageIntLLROutputS1xD(71)(0);
  CNStageIntLLRInputS2xD(95)(1) <= VNStageIntLLROutputS1xD(71)(1);
  CNStageIntLLRInputS2xD(176)(1) <= VNStageIntLLROutputS1xD(71)(2);
  CNStageIntLLRInputS2xD(276)(1) <= VNStageIntLLROutputS1xD(71)(3);
  CNStageIntLLRInputS2xD(302)(1) <= VNStageIntLLROutputS1xD(71)(4);
  CNStageIntLLRInputS2xD(353)(1) <= VNStageIntLLROutputS1xD(71)(5);
  CNStageIntLLRInputS2xD(45)(1) <= VNStageIntLLROutputS1xD(72)(0);
  CNStageIntLLRInputS2xD(75)(1) <= VNStageIntLLROutputS1xD(72)(1);
  CNStageIntLLRInputS2xD(162)(1) <= VNStageIntLLROutputS1xD(72)(2);
  CNStageIntLLRInputS2xD(183)(1) <= VNStageIntLLROutputS1xD(72)(3);
  CNStageIntLLRInputS2xD(243)(1) <= VNStageIntLLROutputS1xD(72)(4);
  CNStageIntLLRInputS2xD(367)(1) <= VNStageIntLLROutputS1xD(72)(5);
  CNStageIntLLRInputS2xD(44)(1) <= VNStageIntLLROutputS1xD(73)(0);
  CNStageIntLLRInputS2xD(56)(1) <= VNStageIntLLROutputS1xD(73)(1);
  CNStageIntLLRInputS2xD(121)(1) <= VNStageIntLLROutputS1xD(73)(2);
  CNStageIntLLRInputS2xD(219)(1) <= VNStageIntLLROutputS1xD(73)(3);
  CNStageIntLLRInputS2xD(328)(1) <= VNStageIntLLROutputS1xD(73)(4);
  CNStageIntLLRInputS2xD(363)(1) <= VNStageIntLLROutputS1xD(73)(5);
  CNStageIntLLRInputS2xD(43)(1) <= VNStageIntLLROutputS1xD(74)(0);
  CNStageIntLLRInputS2xD(70)(1) <= VNStageIntLLROutputS1xD(74)(1);
  CNStageIntLLRInputS2xD(125)(1) <= VNStageIntLLROutputS1xD(74)(2);
  CNStageIntLLRInputS2xD(221)(1) <= VNStageIntLLROutputS1xD(74)(3);
  CNStageIntLLRInputS2xD(290)(1) <= VNStageIntLLROutputS1xD(74)(4);
  CNStageIntLLRInputS2xD(42)(1) <= VNStageIntLLROutputS1xD(75)(0);
  CNStageIntLLRInputS2xD(81)(1) <= VNStageIntLLROutputS1xD(75)(1);
  CNStageIntLLRInputS2xD(170)(1) <= VNStageIntLLROutputS1xD(75)(2);
  CNStageIntLLRInputS2xD(192)(1) <= VNStageIntLLROutputS1xD(75)(3);
  CNStageIntLLRInputS2xD(278)(1) <= VNStageIntLLROutputS1xD(75)(4);
  CNStageIntLLRInputS2xD(294)(1) <= VNStageIntLLROutputS1xD(75)(5);
  CNStageIntLLRInputS2xD(347)(1) <= VNStageIntLLROutputS1xD(75)(6);
  CNStageIntLLRInputS2xD(41)(1) <= VNStageIntLLROutputS1xD(76)(0);
  CNStageIntLLRInputS2xD(106)(1) <= VNStageIntLLROutputS1xD(76)(1);
  CNStageIntLLRInputS2xD(124)(1) <= VNStageIntLLROutputS1xD(76)(2);
  CNStageIntLLRInputS2xD(174)(1) <= VNStageIntLLROutputS1xD(76)(3);
  CNStageIntLLRInputS2xD(270)(1) <= VNStageIntLLROutputS1xD(76)(4);
  CNStageIntLLRInputS2xD(332)(1) <= VNStageIntLLROutputS1xD(76)(5);
  CNStageIntLLRInputS2xD(348)(1) <= VNStageIntLLROutputS1xD(76)(6);
  CNStageIntLLRInputS2xD(119)(1) <= VNStageIntLLROutputS1xD(77)(0);
  CNStageIntLLRInputS2xD(185)(1) <= VNStageIntLLROutputS1xD(77)(1);
  CNStageIntLLRInputS2xD(257)(1) <= VNStageIntLLROutputS1xD(77)(2);
  CNStageIntLLRInputS2xD(293)(1) <= VNStageIntLLROutputS1xD(77)(3);
  CNStageIntLLRInputS2xD(383)(1) <= VNStageIntLLROutputS1xD(77)(4);
  CNStageIntLLRInputS2xD(40)(1) <= VNStageIntLLROutputS1xD(78)(0);
  CNStageIntLLRInputS2xD(84)(1) <= VNStageIntLLROutputS1xD(78)(1);
  CNStageIntLLRInputS2xD(159)(1) <= VNStageIntLLROutputS1xD(78)(2);
  CNStageIntLLRInputS2xD(193)(1) <= VNStageIntLLROutputS1xD(78)(3);
  CNStageIntLLRInputS2xD(274)(1) <= VNStageIntLLROutputS1xD(78)(4);
  CNStageIntLLRInputS2xD(288)(1) <= VNStageIntLLROutputS1xD(78)(5);
  CNStageIntLLRInputS2xD(374)(1) <= VNStageIntLLROutputS1xD(78)(6);
  CNStageIntLLRInputS2xD(39)(1) <= VNStageIntLLROutputS1xD(79)(0);
  CNStageIntLLRInputS2xD(99)(1) <= VNStageIntLLROutputS1xD(79)(1);
  CNStageIntLLRInputS2xD(167)(1) <= VNStageIntLLROutputS1xD(79)(2);
  CNStageIntLLRInputS2xD(220)(1) <= VNStageIntLLROutputS1xD(79)(3);
  CNStageIntLLRInputS2xD(325)(1) <= VNStageIntLLROutputS1xD(79)(4);
  CNStageIntLLRInputS2xD(38)(1) <= VNStageIntLLROutputS1xD(80)(0);
  CNStageIntLLRInputS2xD(62)(1) <= VNStageIntLLROutputS1xD(80)(1);
  CNStageIntLLRInputS2xD(131)(1) <= VNStageIntLLROutputS1xD(80)(2);
  CNStageIntLLRInputS2xD(182)(1) <= VNStageIntLLROutputS1xD(80)(3);
  CNStageIntLLRInputS2xD(248)(1) <= VNStageIntLLROutputS1xD(80)(4);
  CNStageIntLLRInputS2xD(337)(1) <= VNStageIntLLROutputS1xD(80)(5);
  CNStageIntLLRInputS2xD(37)(1) <= VNStageIntLLROutputS1xD(81)(0);
  CNStageIntLLRInputS2xD(72)(1) <= VNStageIntLLROutputS1xD(81)(1);
  CNStageIntLLRInputS2xD(129)(1) <= VNStageIntLLROutputS1xD(81)(2);
  CNStageIntLLRInputS2xD(262)(1) <= VNStageIntLLROutputS1xD(81)(3);
  CNStageIntLLRInputS2xD(36)(1) <= VNStageIntLLROutputS1xD(82)(0);
  CNStageIntLLRInputS2xD(67)(1) <= VNStageIntLLROutputS1xD(82)(1);
  CNStageIntLLRInputS2xD(165)(1) <= VNStageIntLLROutputS1xD(82)(2);
  CNStageIntLLRInputS2xD(188)(1) <= VNStageIntLLROutputS1xD(82)(3);
  CNStageIntLLRInputS2xD(254)(1) <= VNStageIntLLROutputS1xD(82)(4);
  CNStageIntLLRInputS2xD(298)(1) <= VNStageIntLLROutputS1xD(82)(5);
  CNStageIntLLRInputS2xD(336)(1) <= VNStageIntLLROutputS1xD(82)(6);
  CNStageIntLLRInputS2xD(35)(1) <= VNStageIntLLROutputS1xD(83)(0);
  CNStageIntLLRInputS2xD(73)(1) <= VNStageIntLLROutputS1xD(83)(1);
  CNStageIntLLRInputS2xD(144)(1) <= VNStageIntLLROutputS1xD(83)(2);
  CNStageIntLLRInputS2xD(208)(1) <= VNStageIntLLROutputS1xD(83)(3);
  CNStageIntLLRInputS2xD(232)(1) <= VNStageIntLLROutputS1xD(83)(4);
  CNStageIntLLRInputS2xD(330)(1) <= VNStageIntLLROutputS1xD(83)(5);
  CNStageIntLLRInputS2xD(34)(1) <= VNStageIntLLROutputS1xD(84)(0);
  CNStageIntLLRInputS2xD(61)(1) <= VNStageIntLLROutputS1xD(84)(1);
  CNStageIntLLRInputS2xD(147)(1) <= VNStageIntLLROutputS1xD(84)(2);
  CNStageIntLLRInputS2xD(222)(1) <= VNStageIntLLROutputS1xD(84)(3);
  CNStageIntLLRInputS2xD(310)(1) <= VNStageIntLLROutputS1xD(84)(4);
  CNStageIntLLRInputS2xD(371)(1) <= VNStageIntLLROutputS1xD(84)(5);
  CNStageIntLLRInputS2xD(33)(1) <= VNStageIntLLROutputS1xD(85)(0);
  CNStageIntLLRInputS2xD(132)(1) <= VNStageIntLLROutputS1xD(85)(1);
  CNStageIntLLRInputS2xD(218)(1) <= VNStageIntLLROutputS1xD(85)(2);
  CNStageIntLLRInputS2xD(235)(1) <= VNStageIntLLROutputS1xD(85)(3);
  CNStageIntLLRInputS2xD(313)(1) <= VNStageIntLLROutputS1xD(85)(4);
  CNStageIntLLRInputS2xD(379)(1) <= VNStageIntLLROutputS1xD(85)(5);
  CNStageIntLLRInputS2xD(32)(1) <= VNStageIntLLROutputS1xD(86)(0);
  CNStageIntLLRInputS2xD(166)(1) <= VNStageIntLLROutputS1xD(86)(1);
  CNStageIntLLRInputS2xD(239)(1) <= VNStageIntLLROutputS1xD(86)(2);
  CNStageIntLLRInputS2xD(343)(1) <= VNStageIntLLROutputS1xD(86)(3);
  CNStageIntLLRInputS2xD(31)(1) <= VNStageIntLLROutputS1xD(87)(0);
  CNStageIntLLRInputS2xD(77)(1) <= VNStageIntLLROutputS1xD(87)(1);
  CNStageIntLLRInputS2xD(128)(1) <= VNStageIntLLROutputS1xD(87)(2);
  CNStageIntLLRInputS2xD(203)(1) <= VNStageIntLLROutputS1xD(87)(3);
  CNStageIntLLRInputS2xD(229)(1) <= VNStageIntLLROutputS1xD(87)(4);
  CNStageIntLLRInputS2xD(331)(1) <= VNStageIntLLROutputS1xD(87)(5);
  CNStageIntLLRInputS2xD(341)(1) <= VNStageIntLLROutputS1xD(87)(6);
  CNStageIntLLRInputS2xD(30)(1) <= VNStageIntLLROutputS1xD(88)(0);
  CNStageIntLLRInputS2xD(79)(1) <= VNStageIntLLROutputS1xD(88)(1);
  CNStageIntLLRInputS2xD(156)(1) <= VNStageIntLLROutputS1xD(88)(2);
  CNStageIntLLRInputS2xD(204)(1) <= VNStageIntLLROutputS1xD(88)(3);
  CNStageIntLLRInputS2xD(263)(1) <= VNStageIntLLROutputS1xD(88)(4);
  CNStageIntLLRInputS2xD(297)(1) <= VNStageIntLLROutputS1xD(88)(5);
  CNStageIntLLRInputS2xD(377)(1) <= VNStageIntLLROutputS1xD(88)(6);
  CNStageIntLLRInputS2xD(29)(1) <= VNStageIntLLROutputS1xD(89)(0);
  CNStageIntLLRInputS2xD(102)(1) <= VNStageIntLLROutputS1xD(89)(1);
  CNStageIntLLRInputS2xD(140)(1) <= VNStageIntLLROutputS1xD(89)(2);
  CNStageIntLLRInputS2xD(184)(1) <= VNStageIntLLROutputS1xD(89)(3);
  CNStageIntLLRInputS2xD(247)(1) <= VNStageIntLLROutputS1xD(89)(4);
  CNStageIntLLRInputS2xD(355)(1) <= VNStageIntLLROutputS1xD(89)(5);
  CNStageIntLLRInputS2xD(28)(1) <= VNStageIntLLROutputS1xD(90)(0);
  CNStageIntLLRInputS2xD(85)(1) <= VNStageIntLLROutputS1xD(90)(1);
  CNStageIntLLRInputS2xD(168)(1) <= VNStageIntLLROutputS1xD(90)(2);
  CNStageIntLLRInputS2xD(175)(1) <= VNStageIntLLROutputS1xD(90)(3);
  CNStageIntLLRInputS2xD(258)(1) <= VNStageIntLLROutputS1xD(90)(4);
  CNStageIntLLRInputS2xD(307)(1) <= VNStageIntLLROutputS1xD(90)(5);
  CNStageIntLLRInputS2xD(358)(1) <= VNStageIntLLROutputS1xD(90)(6);
  CNStageIntLLRInputS2xD(27)(1) <= VNStageIntLLROutputS1xD(91)(0);
  CNStageIntLLRInputS2xD(96)(1) <= VNStageIntLLROutputS1xD(91)(1);
  CNStageIntLLRInputS2xD(158)(1) <= VNStageIntLLROutputS1xD(91)(2);
  CNStageIntLLRInputS2xD(191)(1) <= VNStageIntLLROutputS1xD(91)(3);
  CNStageIntLLRInputS2xD(269)(1) <= VNStageIntLLROutputS1xD(91)(4);
  CNStageIntLLRInputS2xD(280)(1) <= VNStageIntLLROutputS1xD(91)(5);
  CNStageIntLLRInputS2xD(344)(1) <= VNStageIntLLROutputS1xD(91)(6);
  CNStageIntLLRInputS2xD(26)(1) <= VNStageIntLLROutputS1xD(92)(0);
  CNStageIntLLRInputS2xD(103)(1) <= VNStageIntLLROutputS1xD(92)(1);
  CNStageIntLLRInputS2xD(145)(1) <= VNStageIntLLROutputS1xD(92)(2);
  CNStageIntLLRInputS2xD(195)(1) <= VNStageIntLLROutputS1xD(92)(3);
  CNStageIntLLRInputS2xD(242)(1) <= VNStageIntLLROutputS1xD(92)(4);
  CNStageIntLLRInputS2xD(324)(1) <= VNStageIntLLROutputS1xD(92)(5);
  CNStageIntLLRInputS2xD(378)(1) <= VNStageIntLLROutputS1xD(92)(6);
  CNStageIntLLRInputS2xD(25)(1) <= VNStageIntLLROutputS1xD(93)(0);
  CNStageIntLLRInputS2xD(78)(1) <= VNStageIntLLROutputS1xD(93)(1);
  CNStageIntLLRInputS2xD(164)(1) <= VNStageIntLLROutputS1xD(93)(2);
  CNStageIntLLRInputS2xD(224)(1) <= VNStageIntLLROutputS1xD(93)(3);
  CNStageIntLLRInputS2xD(231)(1) <= VNStageIntLLROutputS1xD(93)(4);
  CNStageIntLLRInputS2xD(311)(1) <= VNStageIntLLROutputS1xD(93)(5);
  CNStageIntLLRInputS2xD(340)(1) <= VNStageIntLLROutputS1xD(93)(6);
  CNStageIntLLRInputS2xD(24)(1) <= VNStageIntLLROutputS1xD(94)(0);
  CNStageIntLLRInputS2xD(92)(1) <= VNStageIntLLROutputS1xD(94)(1);
  CNStageIntLLRInputS2xD(194)(1) <= VNStageIntLLROutputS1xD(94)(2);
  CNStageIntLLRInputS2xD(329)(1) <= VNStageIntLLROutputS1xD(94)(3);
  CNStageIntLLRInputS2xD(368)(1) <= VNStageIntLLROutputS1xD(94)(4);
  CNStageIntLLRInputS2xD(23)(1) <= VNStageIntLLROutputS1xD(95)(0);
  CNStageIntLLRInputS2xD(63)(1) <= VNStageIntLLROutputS1xD(95)(1);
  CNStageIntLLRInputS2xD(134)(1) <= VNStageIntLLROutputS1xD(95)(2);
  CNStageIntLLRInputS2xD(190)(1) <= VNStageIntLLROutputS1xD(95)(3);
  CNStageIntLLRInputS2xD(234)(1) <= VNStageIntLLROutputS1xD(95)(4);
  CNStageIntLLRInputS2xD(303)(1) <= VNStageIntLLROutputS1xD(95)(5);
  CNStageIntLLRInputS2xD(352)(1) <= VNStageIntLLROutputS1xD(95)(6);
  CNStageIntLLRInputS2xD(22)(1) <= VNStageIntLLROutputS1xD(96)(0);
  CNStageIntLLRInputS2xD(98)(1) <= VNStageIntLLROutputS1xD(96)(1);
  CNStageIntLLRInputS2xD(150)(1) <= VNStageIntLLROutputS1xD(96)(2);
  CNStageIntLLRInputS2xD(172)(1) <= VNStageIntLLROutputS1xD(96)(3);
  CNStageIntLLRInputS2xD(251)(1) <= VNStageIntLLROutputS1xD(96)(4);
  CNStageIntLLRInputS2xD(380)(1) <= VNStageIntLLROutputS1xD(96)(5);
  CNStageIntLLRInputS2xD(21)(1) <= VNStageIntLLROutputS1xD(97)(0);
  CNStageIntLLRInputS2xD(65)(1) <= VNStageIntLLROutputS1xD(97)(1);
  CNStageIntLLRInputS2xD(142)(1) <= VNStageIntLLROutputS1xD(97)(2);
  CNStageIntLLRInputS2xD(180)(1) <= VNStageIntLLROutputS1xD(97)(3);
  CNStageIntLLRInputS2xD(260)(1) <= VNStageIntLLROutputS1xD(97)(4);
  CNStageIntLLRInputS2xD(316)(1) <= VNStageIntLLROutputS1xD(97)(5);
  CNStageIntLLRInputS2xD(370)(1) <= VNStageIntLLROutputS1xD(97)(6);
  CNStageIntLLRInputS2xD(20)(1) <= VNStageIntLLROutputS1xD(98)(0);
  CNStageIntLLRInputS2xD(116)(1) <= VNStageIntLLROutputS1xD(98)(1);
  CNStageIntLLRInputS2xD(199)(1) <= VNStageIntLLROutputS1xD(98)(2);
  CNStageIntLLRInputS2xD(255)(1) <= VNStageIntLLROutputS1xD(98)(3);
  CNStageIntLLRInputS2xD(308)(1) <= VNStageIntLLROutputS1xD(98)(4);
  CNStageIntLLRInputS2xD(356)(1) <= VNStageIntLLROutputS1xD(98)(5);
  CNStageIntLLRInputS2xD(19)(1) <= VNStageIntLLROutputS1xD(99)(0);
  CNStageIntLLRInputS2xD(76)(1) <= VNStageIntLLROutputS1xD(99)(1);
  CNStageIntLLRInputS2xD(126)(1) <= VNStageIntLLROutputS1xD(99)(2);
  CNStageIntLLRInputS2xD(198)(1) <= VNStageIntLLROutputS1xD(99)(3);
  CNStageIntLLRInputS2xD(261)(1) <= VNStageIntLLROutputS1xD(99)(4);
  CNStageIntLLRInputS2xD(285)(1) <= VNStageIntLLROutputS1xD(99)(5);
  CNStageIntLLRInputS2xD(376)(1) <= VNStageIntLLROutputS1xD(99)(6);
  CNStageIntLLRInputS2xD(18)(1) <= VNStageIntLLROutputS1xD(100)(0);
  CNStageIntLLRInputS2xD(94)(1) <= VNStageIntLLROutputS1xD(100)(1);
  CNStageIntLLRInputS2xD(120)(1) <= VNStageIntLLROutputS1xD(100)(2);
  CNStageIntLLRInputS2xD(178)(1) <= VNStageIntLLROutputS1xD(100)(3);
  CNStageIntLLRInputS2xD(250)(1) <= VNStageIntLLROutputS1xD(100)(4);
  CNStageIntLLRInputS2xD(295)(1) <= VNStageIntLLROutputS1xD(100)(5);
  CNStageIntLLRInputS2xD(349)(1) <= VNStageIntLLROutputS1xD(100)(6);
  CNStageIntLLRInputS2xD(17)(1) <= VNStageIntLLROutputS1xD(101)(0);
  CNStageIntLLRInputS2xD(58)(1) <= VNStageIntLLROutputS1xD(101)(1);
  CNStageIntLLRInputS2xD(123)(1) <= VNStageIntLLROutputS1xD(101)(2);
  CNStageIntLLRInputS2xD(211)(1) <= VNStageIntLLROutputS1xD(101)(3);
  CNStageIntLLRInputS2xD(273)(1) <= VNStageIntLLROutputS1xD(101)(4);
  CNStageIntLLRInputS2xD(289)(1) <= VNStageIntLLROutputS1xD(101)(5);
  CNStageIntLLRInputS2xD(346)(1) <= VNStageIntLLROutputS1xD(101)(6);
  CNStageIntLLRInputS2xD(16)(1) <= VNStageIntLLROutputS1xD(102)(0);
  CNStageIntLLRInputS2xD(59)(1) <= VNStageIntLLROutputS1xD(102)(1);
  CNStageIntLLRInputS2xD(113)(1) <= VNStageIntLLROutputS1xD(102)(2);
  CNStageIntLLRInputS2xD(214)(1) <= VNStageIntLLROutputS1xD(102)(3);
  CNStageIntLLRInputS2xD(226)(1) <= VNStageIntLLROutputS1xD(102)(4);
  CNStageIntLLRInputS2xD(361)(1) <= VNStageIntLLROutputS1xD(102)(5);
  CNStageIntLLRInputS2xD(15)(1) <= VNStageIntLLROutputS1xD(103)(0);
  CNStageIntLLRInputS2xD(93)(1) <= VNStageIntLLROutputS1xD(103)(1);
  CNStageIntLLRInputS2xD(151)(1) <= VNStageIntLLROutputS1xD(103)(2);
  CNStageIntLLRInputS2xD(200)(1) <= VNStageIntLLROutputS1xD(103)(3);
  CNStageIntLLRInputS2xD(265)(1) <= VNStageIntLLROutputS1xD(103)(4);
  CNStageIntLLRInputS2xD(284)(1) <= VNStageIntLLROutputS1xD(103)(5);
  CNStageIntLLRInputS2xD(354)(1) <= VNStageIntLLROutputS1xD(103)(6);
  CNStageIntLLRInputS2xD(14)(1) <= VNStageIntLLROutputS1xD(104)(0);
  CNStageIntLLRInputS2xD(86)(1) <= VNStageIntLLROutputS1xD(104)(1);
  CNStageIntLLRInputS2xD(133)(1) <= VNStageIntLLROutputS1xD(104)(2);
  CNStageIntLLRInputS2xD(179)(1) <= VNStageIntLLROutputS1xD(104)(3);
  CNStageIntLLRInputS2xD(267)(1) <= VNStageIntLLROutputS1xD(104)(4);
  CNStageIntLLRInputS2xD(317)(1) <= VNStageIntLLROutputS1xD(104)(5);
  CNStageIntLLRInputS2xD(13)(1) <= VNStageIntLLROutputS1xD(105)(0);
  CNStageIntLLRInputS2xD(146)(1) <= VNStageIntLLROutputS1xD(105)(1);
  CNStageIntLLRInputS2xD(197)(1) <= VNStageIntLLROutputS1xD(105)(2);
  CNStageIntLLRInputS2xD(237)(1) <= VNStageIntLLROutputS1xD(105)(3);
  CNStageIntLLRInputS2xD(300)(1) <= VNStageIntLLROutputS1xD(105)(4);
  CNStageIntLLRInputS2xD(338)(1) <= VNStageIntLLROutputS1xD(105)(5);
  CNStageIntLLRInputS2xD(12)(1) <= VNStageIntLLROutputS1xD(106)(0);
  CNStageIntLLRInputS2xD(157)(1) <= VNStageIntLLROutputS1xD(106)(1);
  CNStageIntLLRInputS2xD(223)(1) <= VNStageIntLLROutputS1xD(106)(2);
  CNStageIntLLRInputS2xD(272)(1) <= VNStageIntLLROutputS1xD(106)(3);
  CNStageIntLLRInputS2xD(312)(1) <= VNStageIntLLROutputS1xD(106)(4);
  CNStageIntLLRInputS2xD(333)(1) <= VNStageIntLLROutputS1xD(106)(5);
  CNStageIntLLRInputS2xD(110)(1) <= VNStageIntLLROutputS1xD(107)(0);
  CNStageIntLLRInputS2xD(127)(1) <= VNStageIntLLROutputS1xD(107)(1);
  CNStageIntLLRInputS2xD(207)(1) <= VNStageIntLLROutputS1xD(107)(2);
  CNStageIntLLRInputS2xD(230)(1) <= VNStageIntLLROutputS1xD(107)(3);
  CNStageIntLLRInputS2xD(323)(1) <= VNStageIntLLROutputS1xD(107)(4);
  CNStageIntLLRInputS2xD(335)(1) <= VNStageIntLLROutputS1xD(107)(5);
  CNStageIntLLRInputS2xD(11)(1) <= VNStageIntLLROutputS1xD(108)(0);
  CNStageIntLLRInputS2xD(105)(1) <= VNStageIntLLROutputS1xD(108)(1);
  CNStageIntLLRInputS2xD(115)(1) <= VNStageIntLLROutputS1xD(108)(2);
  CNStageIntLLRInputS2xD(181)(1) <= VNStageIntLLROutputS1xD(108)(3);
  CNStageIntLLRInputS2xD(238)(1) <= VNStageIntLLROutputS1xD(108)(4);
  CNStageIntLLRInputS2xD(296)(1) <= VNStageIntLLROutputS1xD(108)(5);
  CNStageIntLLRInputS2xD(10)(1) <= VNStageIntLLROutputS1xD(109)(0);
  CNStageIntLLRInputS2xD(100)(1) <= VNStageIntLLROutputS1xD(109)(1);
  CNStageIntLLRInputS2xD(160)(1) <= VNStageIntLLROutputS1xD(109)(2);
  CNStageIntLLRInputS2xD(171)(1) <= VNStageIntLLROutputS1xD(109)(3);
  CNStageIntLLRInputS2xD(266)(1) <= VNStageIntLLROutputS1xD(109)(4);
  CNStageIntLLRInputS2xD(362)(1) <= VNStageIntLLROutputS1xD(109)(5);
  CNStageIntLLRInputS2xD(9)(1) <= VNStageIntLLROutputS1xD(110)(0);
  CNStageIntLLRInputS2xD(83)(1) <= VNStageIntLLROutputS1xD(110)(1);
  CNStageIntLLRInputS2xD(118)(1) <= VNStageIntLLROutputS1xD(110)(2);
  CNStageIntLLRInputS2xD(212)(1) <= VNStageIntLLROutputS1xD(110)(3);
  CNStageIntLLRInputS2xD(225)(1) <= VNStageIntLLROutputS1xD(110)(4);
  CNStageIntLLRInputS2xD(326)(1) <= VNStageIntLLROutputS1xD(110)(5);
  CNStageIntLLRInputS2xD(345)(1) <= VNStageIntLLROutputS1xD(110)(6);
  CNStageIntLLRInputS2xD(8)(1) <= VNStageIntLLROutputS1xD(111)(0);
  CNStageIntLLRInputS2xD(90)(1) <= VNStageIntLLROutputS1xD(111)(1);
  CNStageIntLLRInputS2xD(138)(1) <= VNStageIntLLROutputS1xD(111)(2);
  CNStageIntLLRInputS2xD(177)(1) <= VNStageIntLLROutputS1xD(111)(3);
  CNStageIntLLRInputS2xD(252)(1) <= VNStageIntLLROutputS1xD(111)(4);
  CNStageIntLLRInputS2xD(287)(1) <= VNStageIntLLROutputS1xD(111)(5);
  CNStageIntLLRInputS2xD(357)(1) <= VNStageIntLLROutputS1xD(111)(6);
  CNStageIntLLRInputS2xD(7)(1) <= VNStageIntLLROutputS1xD(112)(0);
  CNStageIntLLRInputS2xD(54)(1) <= VNStageIntLLROutputS1xD(112)(1);
  CNStageIntLLRInputS2xD(148)(1) <= VNStageIntLLROutputS1xD(112)(2);
  CNStageIntLLRInputS2xD(205)(1) <= VNStageIntLLROutputS1xD(112)(3);
  CNStageIntLLRInputS2xD(233)(1) <= VNStageIntLLROutputS1xD(112)(4);
  CNStageIntLLRInputS2xD(305)(1) <= VNStageIntLLROutputS1xD(112)(5);
  CNStageIntLLRInputS2xD(369)(1) <= VNStageIntLLROutputS1xD(112)(6);
  CNStageIntLLRInputS2xD(6)(1) <= VNStageIntLLROutputS1xD(113)(0);
  CNStageIntLLRInputS2xD(108)(1) <= VNStageIntLLROutputS1xD(113)(1);
  CNStageIntLLRInputS2xD(143)(1) <= VNStageIntLLROutputS1xD(113)(2);
  CNStageIntLLRInputS2xD(202)(1) <= VNStageIntLLROutputS1xD(113)(3);
  CNStageIntLLRInputS2xD(253)(1) <= VNStageIntLLROutputS1xD(113)(4);
  CNStageIntLLRInputS2xD(314)(1) <= VNStageIntLLROutputS1xD(113)(5);
  CNStageIntLLRInputS2xD(339)(1) <= VNStageIntLLROutputS1xD(113)(6);
  CNStageIntLLRInputS2xD(5)(1) <= VNStageIntLLROutputS1xD(114)(0);
  CNStageIntLLRInputS2xD(88)(1) <= VNStageIntLLROutputS1xD(114)(1);
  CNStageIntLLRInputS2xD(149)(1) <= VNStageIntLLROutputS1xD(114)(2);
  CNStageIntLLRInputS2xD(216)(1) <= VNStageIntLLROutputS1xD(114)(3);
  CNStageIntLLRInputS2xD(268)(1) <= VNStageIntLLROutputS1xD(114)(4);
  CNStageIntLLRInputS2xD(309)(1) <= VNStageIntLLROutputS1xD(114)(5);
  CNStageIntLLRInputS2xD(4)(1) <= VNStageIntLLROutputS1xD(115)(0);
  CNStageIntLLRInputS2xD(68)(1) <= VNStageIntLLROutputS1xD(115)(1);
  CNStageIntLLRInputS2xD(137)(1) <= VNStageIntLLROutputS1xD(115)(2);
  CNStageIntLLRInputS2xD(209)(1) <= VNStageIntLLROutputS1xD(115)(3);
  CNStageIntLLRInputS2xD(264)(1) <= VNStageIntLLROutputS1xD(115)(4);
  CNStageIntLLRInputS2xD(315)(1) <= VNStageIntLLROutputS1xD(115)(5);
  CNStageIntLLRInputS2xD(372)(1) <= VNStageIntLLROutputS1xD(115)(6);
  CNStageIntLLRInputS2xD(71)(1) <= VNStageIntLLROutputS1xD(116)(0);
  CNStageIntLLRInputS2xD(163)(1) <= VNStageIntLLROutputS1xD(116)(1);
  CNStageIntLLRInputS2xD(187)(1) <= VNStageIntLLROutputS1xD(116)(2);
  CNStageIntLLRInputS2xD(228)(1) <= VNStageIntLLROutputS1xD(116)(3);
  CNStageIntLLRInputS2xD(304)(1) <= VNStageIntLLROutputS1xD(116)(4);
  CNStageIntLLRInputS2xD(3)(1) <= VNStageIntLLROutputS1xD(117)(0);
  CNStageIntLLRInputS2xD(55)(1) <= VNStageIntLLROutputS1xD(117)(1);
  CNStageIntLLRInputS2xD(111)(1) <= VNStageIntLLROutputS1xD(117)(2);
  CNStageIntLLRInputS2xD(196)(1) <= VNStageIntLLROutputS1xD(117)(3);
  CNStageIntLLRInputS2xD(2)(1) <= VNStageIntLLROutputS1xD(118)(0);
  CNStageIntLLRInputS2xD(89)(1) <= VNStageIntLLROutputS1xD(118)(1);
  CNStageIntLLRInputS2xD(152)(1) <= VNStageIntLLROutputS1xD(118)(2);
  CNStageIntLLRInputS2xD(249)(1) <= VNStageIntLLROutputS1xD(118)(3);
  CNStageIntLLRInputS2xD(282)(1) <= VNStageIntLLROutputS1xD(118)(4);
  CNStageIntLLRInputS2xD(359)(1) <= VNStageIntLLROutputS1xD(118)(5);
  CNStageIntLLRInputS2xD(1)(1) <= VNStageIntLLROutputS1xD(119)(0);
  CNStageIntLLRInputS2xD(107)(1) <= VNStageIntLLROutputS1xD(119)(1);
  CNStageIntLLRInputS2xD(154)(1) <= VNStageIntLLROutputS1xD(119)(2);
  CNStageIntLLRInputS2xD(227)(1) <= VNStageIntLLROutputS1xD(119)(3);
  CNStageIntLLRInputS2xD(319)(1) <= VNStageIntLLROutputS1xD(119)(4);
  CNStageIntLLRInputS2xD(0)(1) <= VNStageIntLLROutputS1xD(120)(0);
  CNStageIntLLRInputS2xD(80)(1) <= VNStageIntLLROutputS1xD(120)(1);
  CNStageIntLLRInputS2xD(321)(1) <= VNStageIntLLROutputS1xD(120)(2);
  CNStageIntLLRInputS2xD(360)(1) <= VNStageIntLLROutputS1xD(120)(3);
  CNStageIntLLRInputS2xD(64)(1) <= VNStageIntLLROutputS1xD(121)(0);
  CNStageIntLLRInputS2xD(161)(1) <= VNStageIntLLROutputS1xD(121)(1);
  CNStageIntLLRInputS2xD(217)(1) <= VNStageIntLLROutputS1xD(121)(2);
  CNStageIntLLRInputS2xD(236)(1) <= VNStageIntLLROutputS1xD(121)(3);
  CNStageIntLLRInputS2xD(291)(1) <= VNStageIntLLROutputS1xD(121)(4);
  CNStageIntLLRInputS2xD(350)(1) <= VNStageIntLLROutputS1xD(121)(5);
  CNStageIntLLRInputS2xD(91)(1) <= VNStageIntLLROutputS1xD(122)(0);
  CNStageIntLLRInputS2xD(114)(1) <= VNStageIntLLROutputS1xD(122)(1);
  CNStageIntLLRInputS2xD(201)(1) <= VNStageIntLLROutputS1xD(122)(2);
  CNStageIntLLRInputS2xD(241)(1) <= VNStageIntLLROutputS1xD(122)(3);
  CNStageIntLLRInputS2xD(327)(1) <= VNStageIntLLROutputS1xD(122)(4);
  CNStageIntLLRInputS2xD(375)(1) <= VNStageIntLLROutputS1xD(122)(5);
  CNStageIntLLRInputS2xD(82)(1) <= VNStageIntLLROutputS1xD(123)(0);
  CNStageIntLLRInputS2xD(122)(1) <= VNStageIntLLROutputS1xD(123)(1);
  CNStageIntLLRInputS2xD(213)(1) <= VNStageIntLLROutputS1xD(123)(2);
  CNStageIntLLRInputS2xD(279)(1) <= VNStageIntLLROutputS1xD(123)(3);
  CNStageIntLLRInputS2xD(382)(1) <= VNStageIntLLROutputS1xD(123)(4);
  CNStageIntLLRInputS2xD(69)(1) <= VNStageIntLLROutputS1xD(124)(0);
  CNStageIntLLRInputS2xD(153)(1) <= VNStageIntLLROutputS1xD(124)(1);
  CNStageIntLLRInputS2xD(240)(1) <= VNStageIntLLROutputS1xD(124)(2);
  CNStageIntLLRInputS2xD(292)(1) <= VNStageIntLLROutputS1xD(124)(3);
  CNStageIntLLRInputS2xD(364)(1) <= VNStageIntLLROutputS1xD(124)(4);
  CNStageIntLLRInputS2xD(87)(1) <= VNStageIntLLROutputS1xD(125)(0);
  CNStageIntLLRInputS2xD(169)(1) <= VNStageIntLLROutputS1xD(125)(1);
  CNStageIntLLRInputS2xD(320)(1) <= VNStageIntLLROutputS1xD(125)(2);
  CNStageIntLLRInputS2xD(366)(1) <= VNStageIntLLROutputS1xD(125)(3);
  CNStageIntLLRInputS2xD(60)(1) <= VNStageIntLLROutputS1xD(126)(0);
  CNStageIntLLRInputS2xD(139)(1) <= VNStageIntLLROutputS1xD(126)(1);
  CNStageIntLLRInputS2xD(186)(1) <= VNStageIntLLROutputS1xD(126)(2);
  CNStageIntLLRInputS2xD(271)(1) <= VNStageIntLLROutputS1xD(126)(3);
  CNStageIntLLRInputS2xD(281)(1) <= VNStageIntLLROutputS1xD(126)(4);
  CNStageIntLLRInputS2xD(334)(1) <= VNStageIntLLROutputS1xD(126)(5);
  CNStageIntLLRInputS2xD(52)(1) <= VNStageIntLLROutputS1xD(127)(0);
  CNStageIntLLRInputS2xD(57)(1) <= VNStageIntLLROutputS1xD(127)(1);
  CNStageIntLLRInputS2xD(117)(1) <= VNStageIntLLROutputS1xD(127)(2);
  CNStageIntLLRInputS2xD(173)(1) <= VNStageIntLLROutputS1xD(127)(3);
  CNStageIntLLRInputS2xD(277)(1) <= VNStageIntLLROutputS1xD(127)(4);
  CNStageIntLLRInputS2xD(306)(1) <= VNStageIntLLROutputS1xD(127)(5);
  CNStageIntLLRInputS2xD(373)(1) <= VNStageIntLLROutputS1xD(127)(6);
  CNStageIntLLRInputS2xD(53)(2) <= VNStageIntLLROutputS1xD(128)(0);
  CNStageIntLLRInputS2xD(108)(2) <= VNStageIntLLROutputS1xD(128)(1);
  CNStageIntLLRInputS2xD(129)(2) <= VNStageIntLLROutputS1xD(128)(2);
  CNStageIntLLRInputS2xD(198)(2) <= VNStageIntLLROutputS1xD(128)(3);
  CNStageIntLLRInputS2xD(244)(2) <= VNStageIntLLROutputS1xD(128)(4);
  CNStageIntLLRInputS2xD(298)(2) <= VNStageIntLLROutputS1xD(128)(5);
  CNStageIntLLRInputS2xD(341)(2) <= VNStageIntLLROutputS1xD(128)(6);
  CNStageIntLLRInputS2xD(51)(2) <= VNStageIntLLROutputS1xD(129)(0);
  CNStageIntLLRInputS2xD(56)(2) <= VNStageIntLLROutputS1xD(129)(1);
  CNStageIntLLRInputS2xD(116)(2) <= VNStageIntLLROutputS1xD(129)(2);
  CNStageIntLLRInputS2xD(172)(2) <= VNStageIntLLROutputS1xD(129)(3);
  CNStageIntLLRInputS2xD(276)(2) <= VNStageIntLLROutputS1xD(129)(4);
  CNStageIntLLRInputS2xD(305)(2) <= VNStageIntLLROutputS1xD(129)(5);
  CNStageIntLLRInputS2xD(372)(2) <= VNStageIntLLROutputS1xD(129)(6);
  CNStageIntLLRInputS2xD(50)(2) <= VNStageIntLLROutputS1xD(130)(0);
  CNStageIntLLRInputS2xD(73)(2) <= VNStageIntLLROutputS1xD(130)(1);
  CNStageIntLLRInputS2xD(140)(2) <= VNStageIntLLROutputS1xD(130)(2);
  CNStageIntLLRInputS2xD(188)(2) <= VNStageIntLLROutputS1xD(130)(3);
  CNStageIntLLRInputS2xD(245)(2) <= VNStageIntLLROutputS1xD(130)(4);
  CNStageIntLLRInputS2xD(285)(2) <= VNStageIntLLROutputS1xD(130)(5);
  CNStageIntLLRInputS2xD(65)(2) <= VNStageIntLLROutputS1xD(131)(0);
  CNStageIntLLRInputS2xD(154)(2) <= VNStageIntLLROutputS1xD(131)(1);
  CNStageIntLLRInputS2xD(206)(2) <= VNStageIntLLROutputS1xD(131)(2);
  CNStageIntLLRInputS2xD(243)(2) <= VNStageIntLLROutputS1xD(131)(3);
  CNStageIntLLRInputS2xD(307)(2) <= VNStageIntLLROutputS1xD(131)(4);
  CNStageIntLLRInputS2xD(334)(2) <= VNStageIntLLROutputS1xD(131)(5);
  CNStageIntLLRInputS2xD(49)(2) <= VNStageIntLLROutputS1xD(132)(0);
  CNStageIntLLRInputS2xD(151)(2) <= VNStageIntLLROutputS1xD(132)(1);
  CNStageIntLLRInputS2xD(214)(2) <= VNStageIntLLROutputS1xD(132)(2);
  CNStageIntLLRInputS2xD(274)(2) <= VNStageIntLLROutputS1xD(132)(3);
  CNStageIntLLRInputS2xD(321)(2) <= VNStageIntLLROutputS1xD(132)(4);
  CNStageIntLLRInputS2xD(364)(2) <= VNStageIntLLROutputS1xD(132)(5);
  CNStageIntLLRInputS2xD(48)(2) <= VNStageIntLLROutputS1xD(133)(0);
  CNStageIntLLRInputS2xD(209)(2) <= VNStageIntLLROutputS1xD(133)(1);
  CNStageIntLLRInputS2xD(255)(2) <= VNStageIntLLROutputS1xD(133)(2);
  CNStageIntLLRInputS2xD(317)(2) <= VNStageIntLLROutputS1xD(133)(3);
  CNStageIntLLRInputS2xD(380)(2) <= VNStageIntLLROutputS1xD(133)(4);
  CNStageIntLLRInputS2xD(47)(2) <= VNStageIntLLROutputS1xD(134)(0);
  CNStageIntLLRInputS2xD(100)(2) <= VNStageIntLLROutputS1xD(134)(1);
  CNStageIntLLRInputS2xD(134)(2) <= VNStageIntLLROutputS1xD(134)(2);
  CNStageIntLLRInputS2xD(258)(2) <= VNStageIntLLROutputS1xD(134)(3);
  CNStageIntLLRInputS2xD(46)(2) <= VNStageIntLLROutputS1xD(135)(0);
  CNStageIntLLRInputS2xD(103)(2) <= VNStageIntLLROutputS1xD(135)(1);
  CNStageIntLLRInputS2xD(135)(2) <= VNStageIntLLROutputS1xD(135)(2);
  CNStageIntLLRInputS2xD(205)(2) <= VNStageIntLLROutputS1xD(135)(3);
  CNStageIntLLRInputS2xD(45)(2) <= VNStageIntLLROutputS1xD(136)(0);
  CNStageIntLLRInputS2xD(94)(2) <= VNStageIntLLROutputS1xD(136)(1);
  CNStageIntLLRInputS2xD(111)(2) <= VNStageIntLLROutputS1xD(136)(2);
  CNStageIntLLRInputS2xD(175)(2) <= VNStageIntLLROutputS1xD(136)(3);
  CNStageIntLLRInputS2xD(275)(2) <= VNStageIntLLROutputS1xD(136)(4);
  CNStageIntLLRInputS2xD(301)(2) <= VNStageIntLLROutputS1xD(136)(5);
  CNStageIntLLRInputS2xD(352)(2) <= VNStageIntLLROutputS1xD(136)(6);
  CNStageIntLLRInputS2xD(44)(2) <= VNStageIntLLROutputS1xD(137)(0);
  CNStageIntLLRInputS2xD(74)(2) <= VNStageIntLLROutputS1xD(137)(1);
  CNStageIntLLRInputS2xD(161)(2) <= VNStageIntLLROutputS1xD(137)(2);
  CNStageIntLLRInputS2xD(182)(2) <= VNStageIntLLROutputS1xD(137)(3);
  CNStageIntLLRInputS2xD(242)(2) <= VNStageIntLLROutputS1xD(137)(4);
  CNStageIntLLRInputS2xD(282)(2) <= VNStageIntLLROutputS1xD(137)(5);
  CNStageIntLLRInputS2xD(366)(2) <= VNStageIntLLROutputS1xD(137)(6);
  CNStageIntLLRInputS2xD(43)(2) <= VNStageIntLLROutputS1xD(138)(0);
  CNStageIntLLRInputS2xD(55)(2) <= VNStageIntLLROutputS1xD(138)(1);
  CNStageIntLLRInputS2xD(120)(2) <= VNStageIntLLROutputS1xD(138)(2);
  CNStageIntLLRInputS2xD(218)(2) <= VNStageIntLLROutputS1xD(138)(3);
  CNStageIntLLRInputS2xD(268)(2) <= VNStageIntLLROutputS1xD(138)(4);
  CNStageIntLLRInputS2xD(327)(2) <= VNStageIntLLROutputS1xD(138)(5);
  CNStageIntLLRInputS2xD(362)(2) <= VNStageIntLLROutputS1xD(138)(6);
  CNStageIntLLRInputS2xD(42)(2) <= VNStageIntLLROutputS1xD(139)(0);
  CNStageIntLLRInputS2xD(69)(2) <= VNStageIntLLROutputS1xD(139)(1);
  CNStageIntLLRInputS2xD(124)(2) <= VNStageIntLLROutputS1xD(139)(2);
  CNStageIntLLRInputS2xD(220)(2) <= VNStageIntLLROutputS1xD(139)(3);
  CNStageIntLLRInputS2xD(252)(2) <= VNStageIntLLROutputS1xD(139)(4);
  CNStageIntLLRInputS2xD(289)(2) <= VNStageIntLLROutputS1xD(139)(5);
  CNStageIntLLRInputS2xD(383)(2) <= VNStageIntLLROutputS1xD(139)(6);
  CNStageIntLLRInputS2xD(41)(2) <= VNStageIntLLROutputS1xD(140)(0);
  CNStageIntLLRInputS2xD(80)(2) <= VNStageIntLLROutputS1xD(140)(1);
  CNStageIntLLRInputS2xD(170)(2) <= VNStageIntLLROutputS1xD(140)(2);
  CNStageIntLLRInputS2xD(191)(2) <= VNStageIntLLROutputS1xD(140)(3);
  CNStageIntLLRInputS2xD(277)(2) <= VNStageIntLLROutputS1xD(140)(4);
  CNStageIntLLRInputS2xD(293)(2) <= VNStageIntLLROutputS1xD(140)(5);
  CNStageIntLLRInputS2xD(346)(2) <= VNStageIntLLROutputS1xD(140)(6);
  CNStageIntLLRInputS2xD(123)(2) <= VNStageIntLLROutputS1xD(141)(0);
  CNStageIntLLRInputS2xD(173)(2) <= VNStageIntLLROutputS1xD(141)(1);
  CNStageIntLLRInputS2xD(269)(2) <= VNStageIntLLROutputS1xD(141)(2);
  CNStageIntLLRInputS2xD(332)(2) <= VNStageIntLLROutputS1xD(141)(3);
  CNStageIntLLRInputS2xD(347)(2) <= VNStageIntLLROutputS1xD(141)(4);
  CNStageIntLLRInputS2xD(40)(2) <= VNStageIntLLROutputS1xD(142)(0);
  CNStageIntLLRInputS2xD(96)(2) <= VNStageIntLLROutputS1xD(142)(1);
  CNStageIntLLRInputS2xD(118)(2) <= VNStageIntLLROutputS1xD(142)(2);
  CNStageIntLLRInputS2xD(256)(2) <= VNStageIntLLROutputS1xD(142)(3);
  CNStageIntLLRInputS2xD(382)(2) <= VNStageIntLLROutputS1xD(142)(4);
  CNStageIntLLRInputS2xD(39)(2) <= VNStageIntLLROutputS1xD(143)(0);
  CNStageIntLLRInputS2xD(83)(2) <= VNStageIntLLROutputS1xD(143)(1);
  CNStageIntLLRInputS2xD(158)(2) <= VNStageIntLLROutputS1xD(143)(2);
  CNStageIntLLRInputS2xD(192)(2) <= VNStageIntLLROutputS1xD(143)(3);
  CNStageIntLLRInputS2xD(273)(2) <= VNStageIntLLROutputS1xD(143)(4);
  CNStageIntLLRInputS2xD(287)(2) <= VNStageIntLLROutputS1xD(143)(5);
  CNStageIntLLRInputS2xD(373)(2) <= VNStageIntLLROutputS1xD(143)(6);
  CNStageIntLLRInputS2xD(38)(2) <= VNStageIntLLROutputS1xD(144)(0);
  CNStageIntLLRInputS2xD(98)(2) <= VNStageIntLLROutputS1xD(144)(1);
  CNStageIntLLRInputS2xD(166)(2) <= VNStageIntLLROutputS1xD(144)(2);
  CNStageIntLLRInputS2xD(219)(2) <= VNStageIntLLROutputS1xD(144)(3);
  CNStageIntLLRInputS2xD(249)(2) <= VNStageIntLLROutputS1xD(144)(4);
  CNStageIntLLRInputS2xD(324)(2) <= VNStageIntLLROutputS1xD(144)(5);
  CNStageIntLLRInputS2xD(333)(2) <= VNStageIntLLROutputS1xD(144)(6);
  CNStageIntLLRInputS2xD(37)(2) <= VNStageIntLLROutputS1xD(145)(0);
  CNStageIntLLRInputS2xD(61)(2) <= VNStageIntLLROutputS1xD(145)(1);
  CNStageIntLLRInputS2xD(130)(2) <= VNStageIntLLROutputS1xD(145)(2);
  CNStageIntLLRInputS2xD(181)(2) <= VNStageIntLLROutputS1xD(145)(3);
  CNStageIntLLRInputS2xD(247)(2) <= VNStageIntLLROutputS1xD(145)(4);
  CNStageIntLLRInputS2xD(331)(2) <= VNStageIntLLROutputS1xD(145)(5);
  CNStageIntLLRInputS2xD(336)(2) <= VNStageIntLLROutputS1xD(145)(6);
  CNStageIntLLRInputS2xD(36)(2) <= VNStageIntLLROutputS1xD(146)(0);
  CNStageIntLLRInputS2xD(71)(2) <= VNStageIntLLROutputS1xD(146)(1);
  CNStageIntLLRInputS2xD(128)(2) <= VNStageIntLLROutputS1xD(146)(2);
  CNStageIntLLRInputS2xD(261)(2) <= VNStageIntLLROutputS1xD(146)(3);
  CNStageIntLLRInputS2xD(299)(2) <= VNStageIntLLROutputS1xD(146)(4);
  CNStageIntLLRInputS2xD(35)(2) <= VNStageIntLLROutputS1xD(147)(0);
  CNStageIntLLRInputS2xD(66)(2) <= VNStageIntLLROutputS1xD(147)(1);
  CNStageIntLLRInputS2xD(164)(2) <= VNStageIntLLROutputS1xD(147)(2);
  CNStageIntLLRInputS2xD(187)(2) <= VNStageIntLLROutputS1xD(147)(3);
  CNStageIntLLRInputS2xD(253)(2) <= VNStageIntLLROutputS1xD(147)(4);
  CNStageIntLLRInputS2xD(297)(2) <= VNStageIntLLROutputS1xD(147)(5);
  CNStageIntLLRInputS2xD(335)(2) <= VNStageIntLLROutputS1xD(147)(6);
  CNStageIntLLRInputS2xD(34)(2) <= VNStageIntLLROutputS1xD(148)(0);
  CNStageIntLLRInputS2xD(72)(2) <= VNStageIntLLROutputS1xD(148)(1);
  CNStageIntLLRInputS2xD(143)(2) <= VNStageIntLLROutputS1xD(148)(2);
  CNStageIntLLRInputS2xD(207)(2) <= VNStageIntLLROutputS1xD(148)(3);
  CNStageIntLLRInputS2xD(231)(2) <= VNStageIntLLROutputS1xD(148)(4);
  CNStageIntLLRInputS2xD(329)(2) <= VNStageIntLLROutputS1xD(148)(5);
  CNStageIntLLRInputS2xD(33)(2) <= VNStageIntLLROutputS1xD(149)(0);
  CNStageIntLLRInputS2xD(60)(2) <= VNStageIntLLROutputS1xD(149)(1);
  CNStageIntLLRInputS2xD(146)(2) <= VNStageIntLLROutputS1xD(149)(2);
  CNStageIntLLRInputS2xD(221)(2) <= VNStageIntLLROutputS1xD(149)(3);
  CNStageIntLLRInputS2xD(241)(2) <= VNStageIntLLROutputS1xD(149)(4);
  CNStageIntLLRInputS2xD(309)(2) <= VNStageIntLLROutputS1xD(149)(5);
  CNStageIntLLRInputS2xD(370)(2) <= VNStageIntLLROutputS1xD(149)(6);
  CNStageIntLLRInputS2xD(32)(2) <= VNStageIntLLROutputS1xD(150)(0);
  CNStageIntLLRInputS2xD(86)(2) <= VNStageIntLLROutputS1xD(150)(1);
  CNStageIntLLRInputS2xD(131)(2) <= VNStageIntLLROutputS1xD(150)(2);
  CNStageIntLLRInputS2xD(217)(2) <= VNStageIntLLROutputS1xD(150)(3);
  CNStageIntLLRInputS2xD(312)(2) <= VNStageIntLLROutputS1xD(150)(4);
  CNStageIntLLRInputS2xD(378)(2) <= VNStageIntLLROutputS1xD(150)(5);
  CNStageIntLLRInputS2xD(31)(2) <= VNStageIntLLROutputS1xD(151)(0);
  CNStageIntLLRInputS2xD(92)(2) <= VNStageIntLLROutputS1xD(151)(1);
  CNStageIntLLRInputS2xD(165)(2) <= VNStageIntLLROutputS1xD(151)(2);
  CNStageIntLLRInputS2xD(184)(2) <= VNStageIntLLROutputS1xD(151)(3);
  CNStageIntLLRInputS2xD(238)(2) <= VNStageIntLLROutputS1xD(151)(4);
  CNStageIntLLRInputS2xD(342)(2) <= VNStageIntLLROutputS1xD(151)(5);
  CNStageIntLLRInputS2xD(30)(2) <= VNStageIntLLROutputS1xD(152)(0);
  CNStageIntLLRInputS2xD(76)(2) <= VNStageIntLLROutputS1xD(152)(1);
  CNStageIntLLRInputS2xD(127)(2) <= VNStageIntLLROutputS1xD(152)(2);
  CNStageIntLLRInputS2xD(202)(2) <= VNStageIntLLROutputS1xD(152)(3);
  CNStageIntLLRInputS2xD(228)(2) <= VNStageIntLLROutputS1xD(152)(4);
  CNStageIntLLRInputS2xD(330)(2) <= VNStageIntLLROutputS1xD(152)(5);
  CNStageIntLLRInputS2xD(340)(2) <= VNStageIntLLROutputS1xD(152)(6);
  CNStageIntLLRInputS2xD(29)(2) <= VNStageIntLLROutputS1xD(153)(0);
  CNStageIntLLRInputS2xD(78)(2) <= VNStageIntLLROutputS1xD(153)(1);
  CNStageIntLLRInputS2xD(155)(2) <= VNStageIntLLROutputS1xD(153)(2);
  CNStageIntLLRInputS2xD(203)(2) <= VNStageIntLLROutputS1xD(153)(3);
  CNStageIntLLRInputS2xD(262)(2) <= VNStageIntLLROutputS1xD(153)(4);
  CNStageIntLLRInputS2xD(296)(2) <= VNStageIntLLROutputS1xD(153)(5);
  CNStageIntLLRInputS2xD(376)(2) <= VNStageIntLLROutputS1xD(153)(6);
  CNStageIntLLRInputS2xD(28)(2) <= VNStageIntLLROutputS1xD(154)(0);
  CNStageIntLLRInputS2xD(139)(2) <= VNStageIntLLROutputS1xD(154)(1);
  CNStageIntLLRInputS2xD(183)(2) <= VNStageIntLLROutputS1xD(154)(2);
  CNStageIntLLRInputS2xD(246)(2) <= VNStageIntLLROutputS1xD(154)(3);
  CNStageIntLLRInputS2xD(322)(2) <= VNStageIntLLROutputS1xD(154)(4);
  CNStageIntLLRInputS2xD(27)(2) <= VNStageIntLLROutputS1xD(155)(0);
  CNStageIntLLRInputS2xD(84)(2) <= VNStageIntLLROutputS1xD(155)(1);
  CNStageIntLLRInputS2xD(167)(2) <= VNStageIntLLROutputS1xD(155)(2);
  CNStageIntLLRInputS2xD(174)(2) <= VNStageIntLLROutputS1xD(155)(3);
  CNStageIntLLRInputS2xD(257)(2) <= VNStageIntLLROutputS1xD(155)(4);
  CNStageIntLLRInputS2xD(306)(2) <= VNStageIntLLROutputS1xD(155)(5);
  CNStageIntLLRInputS2xD(357)(2) <= VNStageIntLLROutputS1xD(155)(6);
  CNStageIntLLRInputS2xD(26)(2) <= VNStageIntLLROutputS1xD(156)(0);
  CNStageIntLLRInputS2xD(95)(2) <= VNStageIntLLROutputS1xD(156)(1);
  CNStageIntLLRInputS2xD(157)(2) <= VNStageIntLLROutputS1xD(156)(2);
  CNStageIntLLRInputS2xD(343)(2) <= VNStageIntLLROutputS1xD(156)(3);
  CNStageIntLLRInputS2xD(25)(2) <= VNStageIntLLROutputS1xD(157)(0);
  CNStageIntLLRInputS2xD(102)(2) <= VNStageIntLLROutputS1xD(157)(1);
  CNStageIntLLRInputS2xD(144)(2) <= VNStageIntLLROutputS1xD(157)(2);
  CNStageIntLLRInputS2xD(194)(2) <= VNStageIntLLROutputS1xD(157)(3);
  CNStageIntLLRInputS2xD(323)(2) <= VNStageIntLLROutputS1xD(157)(4);
  CNStageIntLLRInputS2xD(377)(2) <= VNStageIntLLROutputS1xD(157)(5);
  CNStageIntLLRInputS2xD(24)(2) <= VNStageIntLLROutputS1xD(158)(0);
  CNStageIntLLRInputS2xD(77)(2) <= VNStageIntLLROutputS1xD(158)(1);
  CNStageIntLLRInputS2xD(163)(2) <= VNStageIntLLROutputS1xD(158)(2);
  CNStageIntLLRInputS2xD(224)(2) <= VNStageIntLLROutputS1xD(158)(3);
  CNStageIntLLRInputS2xD(230)(2) <= VNStageIntLLROutputS1xD(158)(4);
  CNStageIntLLRInputS2xD(310)(2) <= VNStageIntLLROutputS1xD(158)(5);
  CNStageIntLLRInputS2xD(339)(2) <= VNStageIntLLROutputS1xD(158)(6);
  CNStageIntLLRInputS2xD(23)(2) <= VNStageIntLLROutputS1xD(159)(0);
  CNStageIntLLRInputS2xD(91)(2) <= VNStageIntLLROutputS1xD(159)(1);
  CNStageIntLLRInputS2xD(136)(2) <= VNStageIntLLROutputS1xD(159)(2);
  CNStageIntLLRInputS2xD(271)(2) <= VNStageIntLLROutputS1xD(159)(3);
  CNStageIntLLRInputS2xD(367)(2) <= VNStageIntLLROutputS1xD(159)(4);
  CNStageIntLLRInputS2xD(22)(2) <= VNStageIntLLROutputS1xD(160)(0);
  CNStageIntLLRInputS2xD(62)(2) <= VNStageIntLLROutputS1xD(160)(1);
  CNStageIntLLRInputS2xD(133)(2) <= VNStageIntLLROutputS1xD(160)(2);
  CNStageIntLLRInputS2xD(189)(2) <= VNStageIntLLROutputS1xD(160)(3);
  CNStageIntLLRInputS2xD(233)(2) <= VNStageIntLLROutputS1xD(160)(4);
  CNStageIntLLRInputS2xD(302)(2) <= VNStageIntLLROutputS1xD(160)(5);
  CNStageIntLLRInputS2xD(351)(2) <= VNStageIntLLROutputS1xD(160)(6);
  CNStageIntLLRInputS2xD(21)(2) <= VNStageIntLLROutputS1xD(161)(0);
  CNStageIntLLRInputS2xD(97)(2) <= VNStageIntLLROutputS1xD(161)(1);
  CNStageIntLLRInputS2xD(149)(2) <= VNStageIntLLROutputS1xD(161)(2);
  CNStageIntLLRInputS2xD(171)(2) <= VNStageIntLLROutputS1xD(161)(3);
  CNStageIntLLRInputS2xD(250)(2) <= VNStageIntLLROutputS1xD(161)(4);
  CNStageIntLLRInputS2xD(300)(2) <= VNStageIntLLROutputS1xD(161)(5);
  CNStageIntLLRInputS2xD(379)(2) <= VNStageIntLLROutputS1xD(161)(6);
  CNStageIntLLRInputS2xD(20)(2) <= VNStageIntLLROutputS1xD(162)(0);
  CNStageIntLLRInputS2xD(64)(2) <= VNStageIntLLROutputS1xD(162)(1);
  CNStageIntLLRInputS2xD(141)(2) <= VNStageIntLLROutputS1xD(162)(2);
  CNStageIntLLRInputS2xD(179)(2) <= VNStageIntLLROutputS1xD(162)(3);
  CNStageIntLLRInputS2xD(259)(2) <= VNStageIntLLROutputS1xD(162)(4);
  CNStageIntLLRInputS2xD(315)(2) <= VNStageIntLLROutputS1xD(162)(5);
  CNStageIntLLRInputS2xD(369)(2) <= VNStageIntLLROutputS1xD(162)(6);
  CNStageIntLLRInputS2xD(19)(2) <= VNStageIntLLROutputS1xD(163)(0);
  CNStageIntLLRInputS2xD(79)(2) <= VNStageIntLLROutputS1xD(163)(1);
  CNStageIntLLRInputS2xD(115)(2) <= VNStageIntLLROutputS1xD(163)(2);
  CNStageIntLLRInputS2xD(254)(2) <= VNStageIntLLROutputS1xD(163)(3);
  CNStageIntLLRInputS2xD(355)(2) <= VNStageIntLLROutputS1xD(163)(4);
  CNStageIntLLRInputS2xD(18)(2) <= VNStageIntLLROutputS1xD(164)(0);
  CNStageIntLLRInputS2xD(75)(2) <= VNStageIntLLROutputS1xD(164)(1);
  CNStageIntLLRInputS2xD(125)(2) <= VNStageIntLLROutputS1xD(164)(2);
  CNStageIntLLRInputS2xD(197)(2) <= VNStageIntLLROutputS1xD(164)(3);
  CNStageIntLLRInputS2xD(260)(2) <= VNStageIntLLROutputS1xD(164)(4);
  CNStageIntLLRInputS2xD(375)(2) <= VNStageIntLLROutputS1xD(164)(5);
  CNStageIntLLRInputS2xD(17)(2) <= VNStageIntLLROutputS1xD(165)(0);
  CNStageIntLLRInputS2xD(93)(2) <= VNStageIntLLROutputS1xD(165)(1);
  CNStageIntLLRInputS2xD(119)(2) <= VNStageIntLLROutputS1xD(165)(2);
  CNStageIntLLRInputS2xD(177)(2) <= VNStageIntLLROutputS1xD(165)(3);
  CNStageIntLLRInputS2xD(294)(2) <= VNStageIntLLROutputS1xD(165)(4);
  CNStageIntLLRInputS2xD(348)(2) <= VNStageIntLLROutputS1xD(165)(5);
  CNStageIntLLRInputS2xD(16)(2) <= VNStageIntLLROutputS1xD(166)(0);
  CNStageIntLLRInputS2xD(57)(2) <= VNStageIntLLROutputS1xD(166)(1);
  CNStageIntLLRInputS2xD(122)(2) <= VNStageIntLLROutputS1xD(166)(2);
  CNStageIntLLRInputS2xD(210)(2) <= VNStageIntLLROutputS1xD(166)(3);
  CNStageIntLLRInputS2xD(288)(2) <= VNStageIntLLROutputS1xD(166)(4);
  CNStageIntLLRInputS2xD(345)(2) <= VNStageIntLLROutputS1xD(166)(5);
  CNStageIntLLRInputS2xD(15)(2) <= VNStageIntLLROutputS1xD(167)(0);
  CNStageIntLLRInputS2xD(58)(2) <= VNStageIntLLROutputS1xD(167)(1);
  CNStageIntLLRInputS2xD(112)(2) <= VNStageIntLLROutputS1xD(167)(2);
  CNStageIntLLRInputS2xD(213)(2) <= VNStageIntLLROutputS1xD(167)(3);
  CNStageIntLLRInputS2xD(225)(2) <= VNStageIntLLROutputS1xD(167)(4);
  CNStageIntLLRInputS2xD(292)(2) <= VNStageIntLLROutputS1xD(167)(5);
  CNStageIntLLRInputS2xD(360)(2) <= VNStageIntLLROutputS1xD(167)(6);
  CNStageIntLLRInputS2xD(14)(2) <= VNStageIntLLROutputS1xD(168)(0);
  CNStageIntLLRInputS2xD(150)(2) <= VNStageIntLLROutputS1xD(168)(1);
  CNStageIntLLRInputS2xD(199)(2) <= VNStageIntLLROutputS1xD(168)(2);
  CNStageIntLLRInputS2xD(264)(2) <= VNStageIntLLROutputS1xD(168)(3);
  CNStageIntLLRInputS2xD(283)(2) <= VNStageIntLLROutputS1xD(168)(4);
  CNStageIntLLRInputS2xD(353)(2) <= VNStageIntLLROutputS1xD(168)(5);
  CNStageIntLLRInputS2xD(13)(2) <= VNStageIntLLROutputS1xD(169)(0);
  CNStageIntLLRInputS2xD(85)(2) <= VNStageIntLLROutputS1xD(169)(1);
  CNStageIntLLRInputS2xD(132)(2) <= VNStageIntLLROutputS1xD(169)(2);
  CNStageIntLLRInputS2xD(178)(2) <= VNStageIntLLROutputS1xD(169)(3);
  CNStageIntLLRInputS2xD(266)(2) <= VNStageIntLLROutputS1xD(169)(4);
  CNStageIntLLRInputS2xD(316)(2) <= VNStageIntLLROutputS1xD(169)(5);
  CNStageIntLLRInputS2xD(12)(2) <= VNStageIntLLROutputS1xD(170)(0);
  CNStageIntLLRInputS2xD(101)(2) <= VNStageIntLLROutputS1xD(170)(1);
  CNStageIntLLRInputS2xD(145)(2) <= VNStageIntLLROutputS1xD(170)(2);
  CNStageIntLLRInputS2xD(236)(2) <= VNStageIntLLROutputS1xD(170)(3);
  CNStageIntLLRInputS2xD(337)(2) <= VNStageIntLLROutputS1xD(170)(4);
  CNStageIntLLRInputS2xD(105)(2) <= VNStageIntLLROutputS1xD(171)(0);
  CNStageIntLLRInputS2xD(156)(2) <= VNStageIntLLROutputS1xD(171)(1);
  CNStageIntLLRInputS2xD(222)(2) <= VNStageIntLLROutputS1xD(171)(2);
  CNStageIntLLRInputS2xD(311)(2) <= VNStageIntLLROutputS1xD(171)(3);
  CNStageIntLLRInputS2xD(11)(2) <= VNStageIntLLROutputS1xD(172)(0);
  CNStageIntLLRInputS2xD(110)(2) <= VNStageIntLLROutputS1xD(172)(1);
  CNStageIntLLRInputS2xD(126)(2) <= VNStageIntLLROutputS1xD(172)(2);
  CNStageIntLLRInputS2xD(229)(2) <= VNStageIntLLROutputS1xD(172)(3);
  CNStageIntLLRInputS2xD(10)(2) <= VNStageIntLLROutputS1xD(173)(0);
  CNStageIntLLRInputS2xD(104)(2) <= VNStageIntLLROutputS1xD(173)(1);
  CNStageIntLLRInputS2xD(114)(2) <= VNStageIntLLROutputS1xD(173)(2);
  CNStageIntLLRInputS2xD(180)(2) <= VNStageIntLLROutputS1xD(173)(3);
  CNStageIntLLRInputS2xD(237)(2) <= VNStageIntLLROutputS1xD(173)(4);
  CNStageIntLLRInputS2xD(295)(2) <= VNStageIntLLROutputS1xD(173)(5);
  CNStageIntLLRInputS2xD(9)(2) <= VNStageIntLLROutputS1xD(174)(0);
  CNStageIntLLRInputS2xD(99)(2) <= VNStageIntLLROutputS1xD(174)(1);
  CNStageIntLLRInputS2xD(159)(2) <= VNStageIntLLROutputS1xD(174)(2);
  CNStageIntLLRInputS2xD(265)(2) <= VNStageIntLLROutputS1xD(174)(3);
  CNStageIntLLRInputS2xD(361)(2) <= VNStageIntLLROutputS1xD(174)(4);
  CNStageIntLLRInputS2xD(8)(2) <= VNStageIntLLROutputS1xD(175)(0);
  CNStageIntLLRInputS2xD(82)(2) <= VNStageIntLLROutputS1xD(175)(1);
  CNStageIntLLRInputS2xD(117)(2) <= VNStageIntLLROutputS1xD(175)(2);
  CNStageIntLLRInputS2xD(211)(2) <= VNStageIntLLROutputS1xD(175)(3);
  CNStageIntLLRInputS2xD(278)(2) <= VNStageIntLLROutputS1xD(175)(4);
  CNStageIntLLRInputS2xD(325)(2) <= VNStageIntLLROutputS1xD(175)(5);
  CNStageIntLLRInputS2xD(344)(2) <= VNStageIntLLROutputS1xD(175)(6);
  CNStageIntLLRInputS2xD(7)(2) <= VNStageIntLLROutputS1xD(176)(0);
  CNStageIntLLRInputS2xD(89)(2) <= VNStageIntLLROutputS1xD(176)(1);
  CNStageIntLLRInputS2xD(137)(2) <= VNStageIntLLROutputS1xD(176)(2);
  CNStageIntLLRInputS2xD(176)(2) <= VNStageIntLLROutputS1xD(176)(3);
  CNStageIntLLRInputS2xD(251)(2) <= VNStageIntLLROutputS1xD(176)(4);
  CNStageIntLLRInputS2xD(286)(2) <= VNStageIntLLROutputS1xD(176)(5);
  CNStageIntLLRInputS2xD(356)(2) <= VNStageIntLLROutputS1xD(176)(6);
  CNStageIntLLRInputS2xD(6)(2) <= VNStageIntLLROutputS1xD(177)(0);
  CNStageIntLLRInputS2xD(109)(2) <= VNStageIntLLROutputS1xD(177)(1);
  CNStageIntLLRInputS2xD(147)(2) <= VNStageIntLLROutputS1xD(177)(2);
  CNStageIntLLRInputS2xD(204)(2) <= VNStageIntLLROutputS1xD(177)(3);
  CNStageIntLLRInputS2xD(232)(2) <= VNStageIntLLROutputS1xD(177)(4);
  CNStageIntLLRInputS2xD(304)(2) <= VNStageIntLLROutputS1xD(177)(5);
  CNStageIntLLRInputS2xD(368)(2) <= VNStageIntLLROutputS1xD(177)(6);
  CNStageIntLLRInputS2xD(5)(2) <= VNStageIntLLROutputS1xD(178)(0);
  CNStageIntLLRInputS2xD(107)(2) <= VNStageIntLLROutputS1xD(178)(1);
  CNStageIntLLRInputS2xD(142)(2) <= VNStageIntLLROutputS1xD(178)(2);
  CNStageIntLLRInputS2xD(201)(2) <= VNStageIntLLROutputS1xD(178)(3);
  CNStageIntLLRInputS2xD(313)(2) <= VNStageIntLLROutputS1xD(178)(4);
  CNStageIntLLRInputS2xD(338)(2) <= VNStageIntLLROutputS1xD(178)(5);
  CNStageIntLLRInputS2xD(4)(2) <= VNStageIntLLROutputS1xD(179)(0);
  CNStageIntLLRInputS2xD(87)(2) <= VNStageIntLLROutputS1xD(179)(1);
  CNStageIntLLRInputS2xD(148)(2) <= VNStageIntLLROutputS1xD(179)(2);
  CNStageIntLLRInputS2xD(215)(2) <= VNStageIntLLROutputS1xD(179)(3);
  CNStageIntLLRInputS2xD(267)(2) <= VNStageIntLLROutputS1xD(179)(4);
  CNStageIntLLRInputS2xD(308)(2) <= VNStageIntLLROutputS1xD(179)(5);
  CNStageIntLLRInputS2xD(67)(2) <= VNStageIntLLROutputS1xD(180)(0);
  CNStageIntLLRInputS2xD(208)(2) <= VNStageIntLLROutputS1xD(180)(1);
  CNStageIntLLRInputS2xD(263)(2) <= VNStageIntLLROutputS1xD(180)(2);
  CNStageIntLLRInputS2xD(314)(2) <= VNStageIntLLROutputS1xD(180)(3);
  CNStageIntLLRInputS2xD(371)(2) <= VNStageIntLLROutputS1xD(180)(4);
  CNStageIntLLRInputS2xD(3)(2) <= VNStageIntLLROutputS1xD(181)(0);
  CNStageIntLLRInputS2xD(70)(2) <= VNStageIntLLROutputS1xD(181)(1);
  CNStageIntLLRInputS2xD(162)(2) <= VNStageIntLLROutputS1xD(181)(2);
  CNStageIntLLRInputS2xD(186)(2) <= VNStageIntLLROutputS1xD(181)(3);
  CNStageIntLLRInputS2xD(227)(2) <= VNStageIntLLROutputS1xD(181)(4);
  CNStageIntLLRInputS2xD(303)(2) <= VNStageIntLLROutputS1xD(181)(5);
  CNStageIntLLRInputS2xD(2)(2) <= VNStageIntLLROutputS1xD(182)(0);
  CNStageIntLLRInputS2xD(54)(2) <= VNStageIntLLROutputS1xD(182)(1);
  CNStageIntLLRInputS2xD(169)(2) <= VNStageIntLLROutputS1xD(182)(2);
  CNStageIntLLRInputS2xD(195)(2) <= VNStageIntLLROutputS1xD(182)(3);
  CNStageIntLLRInputS2xD(248)(2) <= VNStageIntLLROutputS1xD(182)(4);
  CNStageIntLLRInputS2xD(328)(2) <= VNStageIntLLROutputS1xD(182)(5);
  CNStageIntLLRInputS2xD(350)(2) <= VNStageIntLLROutputS1xD(182)(6);
  CNStageIntLLRInputS2xD(1)(2) <= VNStageIntLLROutputS1xD(183)(0);
  CNStageIntLLRInputS2xD(88)(2) <= VNStageIntLLROutputS1xD(183)(1);
  CNStageIntLLRInputS2xD(190)(2) <= VNStageIntLLROutputS1xD(183)(2);
  CNStageIntLLRInputS2xD(281)(2) <= VNStageIntLLROutputS1xD(183)(3);
  CNStageIntLLRInputS2xD(358)(2) <= VNStageIntLLROutputS1xD(183)(4);
  CNStageIntLLRInputS2xD(0)(2) <= VNStageIntLLROutputS1xD(184)(0);
  CNStageIntLLRInputS2xD(106)(2) <= VNStageIntLLROutputS1xD(184)(1);
  CNStageIntLLRInputS2xD(153)(2) <= VNStageIntLLROutputS1xD(184)(2);
  CNStageIntLLRInputS2xD(193)(2) <= VNStageIntLLROutputS1xD(184)(3);
  CNStageIntLLRInputS2xD(226)(2) <= VNStageIntLLROutputS1xD(184)(4);
  CNStageIntLLRInputS2xD(318)(2) <= VNStageIntLLROutputS1xD(184)(5);
  CNStageIntLLRInputS2xD(354)(2) <= VNStageIntLLROutputS1xD(184)(6);
  CNStageIntLLRInputS2xD(121)(2) <= VNStageIntLLROutputS1xD(185)(0);
  CNStageIntLLRInputS2xD(272)(2) <= VNStageIntLLROutputS1xD(185)(1);
  CNStageIntLLRInputS2xD(320)(2) <= VNStageIntLLROutputS1xD(185)(2);
  CNStageIntLLRInputS2xD(359)(2) <= VNStageIntLLROutputS1xD(185)(3);
  CNStageIntLLRInputS2xD(63)(2) <= VNStageIntLLROutputS1xD(186)(0);
  CNStageIntLLRInputS2xD(160)(2) <= VNStageIntLLROutputS1xD(186)(1);
  CNStageIntLLRInputS2xD(216)(2) <= VNStageIntLLROutputS1xD(186)(2);
  CNStageIntLLRInputS2xD(235)(2) <= VNStageIntLLROutputS1xD(186)(3);
  CNStageIntLLRInputS2xD(290)(2) <= VNStageIntLLROutputS1xD(186)(4);
  CNStageIntLLRInputS2xD(349)(2) <= VNStageIntLLROutputS1xD(186)(5);
  CNStageIntLLRInputS2xD(90)(2) <= VNStageIntLLROutputS1xD(187)(0);
  CNStageIntLLRInputS2xD(113)(2) <= VNStageIntLLROutputS1xD(187)(1);
  CNStageIntLLRInputS2xD(200)(2) <= VNStageIntLLROutputS1xD(187)(2);
  CNStageIntLLRInputS2xD(240)(2) <= VNStageIntLLROutputS1xD(187)(3);
  CNStageIntLLRInputS2xD(326)(2) <= VNStageIntLLROutputS1xD(187)(4);
  CNStageIntLLRInputS2xD(374)(2) <= VNStageIntLLROutputS1xD(187)(5);
  CNStageIntLLRInputS2xD(81)(2) <= VNStageIntLLROutputS1xD(188)(0);
  CNStageIntLLRInputS2xD(212)(2) <= VNStageIntLLROutputS1xD(188)(1);
  CNStageIntLLRInputS2xD(279)(2) <= VNStageIntLLROutputS1xD(188)(2);
  CNStageIntLLRInputS2xD(284)(2) <= VNStageIntLLROutputS1xD(188)(3);
  CNStageIntLLRInputS2xD(381)(2) <= VNStageIntLLROutputS1xD(188)(4);
  CNStageIntLLRInputS2xD(68)(2) <= VNStageIntLLROutputS1xD(189)(0);
  CNStageIntLLRInputS2xD(152)(2) <= VNStageIntLLROutputS1xD(189)(1);
  CNStageIntLLRInputS2xD(223)(2) <= VNStageIntLLROutputS1xD(189)(2);
  CNStageIntLLRInputS2xD(239)(2) <= VNStageIntLLROutputS1xD(189)(3);
  CNStageIntLLRInputS2xD(291)(2) <= VNStageIntLLROutputS1xD(189)(4);
  CNStageIntLLRInputS2xD(363)(2) <= VNStageIntLLROutputS1xD(189)(5);
  CNStageIntLLRInputS2xD(168)(2) <= VNStageIntLLROutputS1xD(190)(0);
  CNStageIntLLRInputS2xD(196)(2) <= VNStageIntLLROutputS1xD(190)(1);
  CNStageIntLLRInputS2xD(234)(2) <= VNStageIntLLROutputS1xD(190)(2);
  CNStageIntLLRInputS2xD(319)(2) <= VNStageIntLLROutputS1xD(190)(3);
  CNStageIntLLRInputS2xD(365)(2) <= VNStageIntLLROutputS1xD(190)(4);
  CNStageIntLLRInputS2xD(52)(2) <= VNStageIntLLROutputS1xD(191)(0);
  CNStageIntLLRInputS2xD(59)(2) <= VNStageIntLLROutputS1xD(191)(1);
  CNStageIntLLRInputS2xD(138)(2) <= VNStageIntLLROutputS1xD(191)(2);
  CNStageIntLLRInputS2xD(185)(2) <= VNStageIntLLROutputS1xD(191)(3);
  CNStageIntLLRInputS2xD(270)(2) <= VNStageIntLLROutputS1xD(191)(4);
  CNStageIntLLRInputS2xD(280)(2) <= VNStageIntLLROutputS1xD(191)(5);
  CNStageIntLLRInputS2xD(53)(3) <= VNStageIntLLROutputS1xD(192)(0);
  CNStageIntLLRInputS2xD(107)(3) <= VNStageIntLLROutputS1xD(192)(1);
  CNStageIntLLRInputS2xD(128)(3) <= VNStageIntLLROutputS1xD(192)(2);
  CNStageIntLLRInputS2xD(197)(3) <= VNStageIntLLROutputS1xD(192)(3);
  CNStageIntLLRInputS2xD(243)(3) <= VNStageIntLLROutputS1xD(192)(4);
  CNStageIntLLRInputS2xD(297)(3) <= VNStageIntLLROutputS1xD(192)(5);
  CNStageIntLLRInputS2xD(340)(3) <= VNStageIntLLROutputS1xD(192)(6);
  CNStageIntLLRInputS2xD(51)(3) <= VNStageIntLLROutputS1xD(193)(0);
  CNStageIntLLRInputS2xD(58)(3) <= VNStageIntLLROutputS1xD(193)(1);
  CNStageIntLLRInputS2xD(137)(3) <= VNStageIntLLROutputS1xD(193)(2);
  CNStageIntLLRInputS2xD(269)(3) <= VNStageIntLLROutputS1xD(193)(3);
  CNStageIntLLRInputS2xD(333)(3) <= VNStageIntLLROutputS1xD(193)(4);
  CNStageIntLLRInputS2xD(50)(3) <= VNStageIntLLROutputS1xD(194)(0);
  CNStageIntLLRInputS2xD(55)(3) <= VNStageIntLLROutputS1xD(194)(1);
  CNStageIntLLRInputS2xD(115)(3) <= VNStageIntLLROutputS1xD(194)(2);
  CNStageIntLLRInputS2xD(171)(3) <= VNStageIntLLROutputS1xD(194)(3);
  CNStageIntLLRInputS2xD(275)(3) <= VNStageIntLLROutputS1xD(194)(4);
  CNStageIntLLRInputS2xD(304)(3) <= VNStageIntLLROutputS1xD(194)(5);
  CNStageIntLLRInputS2xD(371)(3) <= VNStageIntLLROutputS1xD(194)(6);
  CNStageIntLLRInputS2xD(72)(3) <= VNStageIntLLROutputS1xD(195)(0);
  CNStageIntLLRInputS2xD(139)(3) <= VNStageIntLLROutputS1xD(195)(1);
  CNStageIntLLRInputS2xD(187)(3) <= VNStageIntLLROutputS1xD(195)(2);
  CNStageIntLLRInputS2xD(244)(3) <= VNStageIntLLROutputS1xD(195)(3);
  CNStageIntLLRInputS2xD(49)(3) <= VNStageIntLLROutputS1xD(196)(0);
  CNStageIntLLRInputS2xD(64)(3) <= VNStageIntLLROutputS1xD(196)(1);
  CNStageIntLLRInputS2xD(153)(3) <= VNStageIntLLROutputS1xD(196)(2);
  CNStageIntLLRInputS2xD(205)(3) <= VNStageIntLLROutputS1xD(196)(3);
  CNStageIntLLRInputS2xD(242)(3) <= VNStageIntLLROutputS1xD(196)(4);
  CNStageIntLLRInputS2xD(306)(3) <= VNStageIntLLROutputS1xD(196)(5);
  CNStageIntLLRInputS2xD(48)(3) <= VNStageIntLLROutputS1xD(197)(0);
  CNStageIntLLRInputS2xD(96)(3) <= VNStageIntLLROutputS1xD(197)(1);
  CNStageIntLLRInputS2xD(150)(3) <= VNStageIntLLROutputS1xD(197)(2);
  CNStageIntLLRInputS2xD(213)(3) <= VNStageIntLLROutputS1xD(197)(3);
  CNStageIntLLRInputS2xD(273)(3) <= VNStageIntLLROutputS1xD(197)(4);
  CNStageIntLLRInputS2xD(320)(3) <= VNStageIntLLROutputS1xD(197)(5);
  CNStageIntLLRInputS2xD(363)(3) <= VNStageIntLLROutputS1xD(197)(6);
  CNStageIntLLRInputS2xD(47)(3) <= VNStageIntLLROutputS1xD(198)(0);
  CNStageIntLLRInputS2xD(105)(3) <= VNStageIntLLROutputS1xD(198)(1);
  CNStageIntLLRInputS2xD(111)(3) <= VNStageIntLLROutputS1xD(198)(2);
  CNStageIntLLRInputS2xD(208)(3) <= VNStageIntLLROutputS1xD(198)(3);
  CNStageIntLLRInputS2xD(254)(3) <= VNStageIntLLROutputS1xD(198)(4);
  CNStageIntLLRInputS2xD(316)(3) <= VNStageIntLLROutputS1xD(198)(5);
  CNStageIntLLRInputS2xD(379)(3) <= VNStageIntLLROutputS1xD(198)(6);
  CNStageIntLLRInputS2xD(46)(3) <= VNStageIntLLROutputS1xD(199)(0);
  CNStageIntLLRInputS2xD(99)(3) <= VNStageIntLLROutputS1xD(199)(1);
  CNStageIntLLRInputS2xD(133)(3) <= VNStageIntLLROutputS1xD(199)(2);
  CNStageIntLLRInputS2xD(214)(3) <= VNStageIntLLROutputS1xD(199)(3);
  CNStageIntLLRInputS2xD(257)(3) <= VNStageIntLLROutputS1xD(199)(4);
  CNStageIntLLRInputS2xD(282)(3) <= VNStageIntLLROutputS1xD(199)(5);
  CNStageIntLLRInputS2xD(350)(3) <= VNStageIntLLROutputS1xD(199)(6);
  CNStageIntLLRInputS2xD(45)(3) <= VNStageIntLLROutputS1xD(200)(0);
  CNStageIntLLRInputS2xD(102)(3) <= VNStageIntLLROutputS1xD(200)(1);
  CNStageIntLLRInputS2xD(134)(3) <= VNStageIntLLROutputS1xD(200)(2);
  CNStageIntLLRInputS2xD(204)(3) <= VNStageIntLLROutputS1xD(200)(3);
  CNStageIntLLRInputS2xD(245)(3) <= VNStageIntLLROutputS1xD(200)(4);
  CNStageIntLLRInputS2xD(300)(3) <= VNStageIntLLROutputS1xD(200)(5);
  CNStageIntLLRInputS2xD(44)(3) <= VNStageIntLLROutputS1xD(201)(0);
  CNStageIntLLRInputS2xD(93)(3) <= VNStageIntLLROutputS1xD(201)(1);
  CNStageIntLLRInputS2xD(169)(3) <= VNStageIntLLROutputS1xD(201)(2);
  CNStageIntLLRInputS2xD(174)(3) <= VNStageIntLLROutputS1xD(201)(3);
  CNStageIntLLRInputS2xD(274)(3) <= VNStageIntLLROutputS1xD(201)(4);
  CNStageIntLLRInputS2xD(351)(3) <= VNStageIntLLROutputS1xD(201)(5);
  CNStageIntLLRInputS2xD(43)(3) <= VNStageIntLLROutputS1xD(202)(0);
  CNStageIntLLRInputS2xD(73)(3) <= VNStageIntLLROutputS1xD(202)(1);
  CNStageIntLLRInputS2xD(160)(3) <= VNStageIntLLROutputS1xD(202)(2);
  CNStageIntLLRInputS2xD(181)(3) <= VNStageIntLLROutputS1xD(202)(3);
  CNStageIntLLRInputS2xD(281)(3) <= VNStageIntLLROutputS1xD(202)(4);
  CNStageIntLLRInputS2xD(365)(3) <= VNStageIntLLROutputS1xD(202)(5);
  CNStageIntLLRInputS2xD(42)(3) <= VNStageIntLLROutputS1xD(203)(0);
  CNStageIntLLRInputS2xD(54)(3) <= VNStageIntLLROutputS1xD(203)(1);
  CNStageIntLLRInputS2xD(119)(3) <= VNStageIntLLROutputS1xD(203)(2);
  CNStageIntLLRInputS2xD(217)(3) <= VNStageIntLLROutputS1xD(203)(3);
  CNStageIntLLRInputS2xD(267)(3) <= VNStageIntLLROutputS1xD(203)(4);
  CNStageIntLLRInputS2xD(326)(3) <= VNStageIntLLROutputS1xD(203)(5);
  CNStageIntLLRInputS2xD(361)(3) <= VNStageIntLLROutputS1xD(203)(6);
  CNStageIntLLRInputS2xD(41)(3) <= VNStageIntLLROutputS1xD(204)(0);
  CNStageIntLLRInputS2xD(68)(3) <= VNStageIntLLROutputS1xD(204)(1);
  CNStageIntLLRInputS2xD(123)(3) <= VNStageIntLLROutputS1xD(204)(2);
  CNStageIntLLRInputS2xD(219)(3) <= VNStageIntLLROutputS1xD(204)(3);
  CNStageIntLLRInputS2xD(251)(3) <= VNStageIntLLROutputS1xD(204)(4);
  CNStageIntLLRInputS2xD(288)(3) <= VNStageIntLLROutputS1xD(204)(5);
  CNStageIntLLRInputS2xD(382)(3) <= VNStageIntLLROutputS1xD(204)(6);
  CNStageIntLLRInputS2xD(170)(3) <= VNStageIntLLROutputS1xD(205)(0);
  CNStageIntLLRInputS2xD(276)(3) <= VNStageIntLLROutputS1xD(205)(1);
  CNStageIntLLRInputS2xD(345)(3) <= VNStageIntLLROutputS1xD(205)(2);
  CNStageIntLLRInputS2xD(40)(3) <= VNStageIntLLROutputS1xD(206)(0);
  CNStageIntLLRInputS2xD(122)(3) <= VNStageIntLLROutputS1xD(206)(1);
  CNStageIntLLRInputS2xD(172)(3) <= VNStageIntLLROutputS1xD(206)(2);
  CNStageIntLLRInputS2xD(332)(3) <= VNStageIntLLROutputS1xD(206)(3);
  CNStageIntLLRInputS2xD(346)(3) <= VNStageIntLLROutputS1xD(206)(4);
  CNStageIntLLRInputS2xD(39)(3) <= VNStageIntLLROutputS1xD(207)(0);
  CNStageIntLLRInputS2xD(95)(3) <= VNStageIntLLROutputS1xD(207)(1);
  CNStageIntLLRInputS2xD(117)(3) <= VNStageIntLLROutputS1xD(207)(2);
  CNStageIntLLRInputS2xD(255)(3) <= VNStageIntLLROutputS1xD(207)(3);
  CNStageIntLLRInputS2xD(292)(3) <= VNStageIntLLROutputS1xD(207)(4);
  CNStageIntLLRInputS2xD(381)(3) <= VNStageIntLLROutputS1xD(207)(5);
  CNStageIntLLRInputS2xD(38)(3) <= VNStageIntLLROutputS1xD(208)(0);
  CNStageIntLLRInputS2xD(82)(3) <= VNStageIntLLROutputS1xD(208)(1);
  CNStageIntLLRInputS2xD(157)(3) <= VNStageIntLLROutputS1xD(208)(2);
  CNStageIntLLRInputS2xD(191)(3) <= VNStageIntLLROutputS1xD(208)(3);
  CNStageIntLLRInputS2xD(286)(3) <= VNStageIntLLROutputS1xD(208)(4);
  CNStageIntLLRInputS2xD(372)(3) <= VNStageIntLLROutputS1xD(208)(5);
  CNStageIntLLRInputS2xD(37)(3) <= VNStageIntLLROutputS1xD(209)(0);
  CNStageIntLLRInputS2xD(97)(3) <= VNStageIntLLROutputS1xD(209)(1);
  CNStageIntLLRInputS2xD(165)(3) <= VNStageIntLLROutputS1xD(209)(2);
  CNStageIntLLRInputS2xD(218)(3) <= VNStageIntLLROutputS1xD(209)(3);
  CNStageIntLLRInputS2xD(323)(3) <= VNStageIntLLROutputS1xD(209)(4);
  CNStageIntLLRInputS2xD(36)(3) <= VNStageIntLLROutputS1xD(210)(0);
  CNStageIntLLRInputS2xD(60)(3) <= VNStageIntLLROutputS1xD(210)(1);
  CNStageIntLLRInputS2xD(129)(3) <= VNStageIntLLROutputS1xD(210)(2);
  CNStageIntLLRInputS2xD(180)(3) <= VNStageIntLLROutputS1xD(210)(3);
  CNStageIntLLRInputS2xD(246)(3) <= VNStageIntLLROutputS1xD(210)(4);
  CNStageIntLLRInputS2xD(330)(3) <= VNStageIntLLROutputS1xD(210)(5);
  CNStageIntLLRInputS2xD(335)(3) <= VNStageIntLLROutputS1xD(210)(6);
  CNStageIntLLRInputS2xD(35)(3) <= VNStageIntLLROutputS1xD(211)(0);
  CNStageIntLLRInputS2xD(70)(3) <= VNStageIntLLROutputS1xD(211)(1);
  CNStageIntLLRInputS2xD(127)(3) <= VNStageIntLLROutputS1xD(211)(2);
  CNStageIntLLRInputS2xD(206)(3) <= VNStageIntLLROutputS1xD(211)(3);
  CNStageIntLLRInputS2xD(260)(3) <= VNStageIntLLROutputS1xD(211)(4);
  CNStageIntLLRInputS2xD(298)(3) <= VNStageIntLLROutputS1xD(211)(5);
  CNStageIntLLRInputS2xD(34)(3) <= VNStageIntLLROutputS1xD(212)(0);
  CNStageIntLLRInputS2xD(65)(3) <= VNStageIntLLROutputS1xD(212)(1);
  CNStageIntLLRInputS2xD(163)(3) <= VNStageIntLLROutputS1xD(212)(2);
  CNStageIntLLRInputS2xD(186)(3) <= VNStageIntLLROutputS1xD(212)(3);
  CNStageIntLLRInputS2xD(296)(3) <= VNStageIntLLROutputS1xD(212)(4);
  CNStageIntLLRInputS2xD(33)(3) <= VNStageIntLLROutputS1xD(213)(0);
  CNStageIntLLRInputS2xD(71)(3) <= VNStageIntLLROutputS1xD(213)(1);
  CNStageIntLLRInputS2xD(142)(3) <= VNStageIntLLROutputS1xD(213)(2);
  CNStageIntLLRInputS2xD(230)(3) <= VNStageIntLLROutputS1xD(213)(3);
  CNStageIntLLRInputS2xD(32)(3) <= VNStageIntLLROutputS1xD(214)(0);
  CNStageIntLLRInputS2xD(59)(3) <= VNStageIntLLROutputS1xD(214)(1);
  CNStageIntLLRInputS2xD(145)(3) <= VNStageIntLLROutputS1xD(214)(2);
  CNStageIntLLRInputS2xD(220)(3) <= VNStageIntLLROutputS1xD(214)(3);
  CNStageIntLLRInputS2xD(240)(3) <= VNStageIntLLROutputS1xD(214)(4);
  CNStageIntLLRInputS2xD(308)(3) <= VNStageIntLLROutputS1xD(214)(5);
  CNStageIntLLRInputS2xD(369)(3) <= VNStageIntLLROutputS1xD(214)(6);
  CNStageIntLLRInputS2xD(31)(3) <= VNStageIntLLROutputS1xD(215)(0);
  CNStageIntLLRInputS2xD(85)(3) <= VNStageIntLLROutputS1xD(215)(1);
  CNStageIntLLRInputS2xD(130)(3) <= VNStageIntLLROutputS1xD(215)(2);
  CNStageIntLLRInputS2xD(216)(3) <= VNStageIntLLROutputS1xD(215)(3);
  CNStageIntLLRInputS2xD(234)(3) <= VNStageIntLLROutputS1xD(215)(4);
  CNStageIntLLRInputS2xD(311)(3) <= VNStageIntLLROutputS1xD(215)(5);
  CNStageIntLLRInputS2xD(377)(3) <= VNStageIntLLROutputS1xD(215)(6);
  CNStageIntLLRInputS2xD(30)(3) <= VNStageIntLLROutputS1xD(216)(0);
  CNStageIntLLRInputS2xD(91)(3) <= VNStageIntLLROutputS1xD(216)(1);
  CNStageIntLLRInputS2xD(164)(3) <= VNStageIntLLROutputS1xD(216)(2);
  CNStageIntLLRInputS2xD(183)(3) <= VNStageIntLLROutputS1xD(216)(3);
  CNStageIntLLRInputS2xD(237)(3) <= VNStageIntLLROutputS1xD(216)(4);
  CNStageIntLLRInputS2xD(299)(3) <= VNStageIntLLROutputS1xD(216)(5);
  CNStageIntLLRInputS2xD(341)(3) <= VNStageIntLLROutputS1xD(216)(6);
  CNStageIntLLRInputS2xD(29)(3) <= VNStageIntLLROutputS1xD(217)(0);
  CNStageIntLLRInputS2xD(75)(3) <= VNStageIntLLROutputS1xD(217)(1);
  CNStageIntLLRInputS2xD(126)(3) <= VNStageIntLLROutputS1xD(217)(2);
  CNStageIntLLRInputS2xD(201)(3) <= VNStageIntLLROutputS1xD(217)(3);
  CNStageIntLLRInputS2xD(227)(3) <= VNStageIntLLROutputS1xD(217)(4);
  CNStageIntLLRInputS2xD(329)(3) <= VNStageIntLLROutputS1xD(217)(5);
  CNStageIntLLRInputS2xD(339)(3) <= VNStageIntLLROutputS1xD(217)(6);
  CNStageIntLLRInputS2xD(28)(3) <= VNStageIntLLROutputS1xD(218)(0);
  CNStageIntLLRInputS2xD(77)(3) <= VNStageIntLLROutputS1xD(218)(1);
  CNStageIntLLRInputS2xD(154)(3) <= VNStageIntLLROutputS1xD(218)(2);
  CNStageIntLLRInputS2xD(202)(3) <= VNStageIntLLROutputS1xD(218)(3);
  CNStageIntLLRInputS2xD(261)(3) <= VNStageIntLLROutputS1xD(218)(4);
  CNStageIntLLRInputS2xD(295)(3) <= VNStageIntLLROutputS1xD(218)(5);
  CNStageIntLLRInputS2xD(375)(3) <= VNStageIntLLROutputS1xD(218)(6);
  CNStageIntLLRInputS2xD(27)(3) <= VNStageIntLLROutputS1xD(219)(0);
  CNStageIntLLRInputS2xD(101)(3) <= VNStageIntLLROutputS1xD(219)(1);
  CNStageIntLLRInputS2xD(138)(3) <= VNStageIntLLROutputS1xD(219)(2);
  CNStageIntLLRInputS2xD(182)(3) <= VNStageIntLLROutputS1xD(219)(3);
  CNStageIntLLRInputS2xD(321)(3) <= VNStageIntLLROutputS1xD(219)(4);
  CNStageIntLLRInputS2xD(354)(3) <= VNStageIntLLROutputS1xD(219)(5);
  CNStageIntLLRInputS2xD(26)(3) <= VNStageIntLLROutputS1xD(220)(0);
  CNStageIntLLRInputS2xD(83)(3) <= VNStageIntLLROutputS1xD(220)(1);
  CNStageIntLLRInputS2xD(166)(3) <= VNStageIntLLROutputS1xD(220)(2);
  CNStageIntLLRInputS2xD(173)(3) <= VNStageIntLLROutputS1xD(220)(3);
  CNStageIntLLRInputS2xD(256)(3) <= VNStageIntLLROutputS1xD(220)(4);
  CNStageIntLLRInputS2xD(305)(3) <= VNStageIntLLROutputS1xD(220)(5);
  CNStageIntLLRInputS2xD(356)(3) <= VNStageIntLLROutputS1xD(220)(6);
  CNStageIntLLRInputS2xD(25)(3) <= VNStageIntLLROutputS1xD(221)(0);
  CNStageIntLLRInputS2xD(94)(3) <= VNStageIntLLROutputS1xD(221)(1);
  CNStageIntLLRInputS2xD(156)(3) <= VNStageIntLLROutputS1xD(221)(2);
  CNStageIntLLRInputS2xD(190)(3) <= VNStageIntLLROutputS1xD(221)(3);
  CNStageIntLLRInputS2xD(268)(3) <= VNStageIntLLROutputS1xD(221)(4);
  CNStageIntLLRInputS2xD(331)(3) <= VNStageIntLLROutputS1xD(221)(5);
  CNStageIntLLRInputS2xD(342)(3) <= VNStageIntLLROutputS1xD(221)(6);
  CNStageIntLLRInputS2xD(24)(3) <= VNStageIntLLROutputS1xD(222)(0);
  CNStageIntLLRInputS2xD(143)(3) <= VNStageIntLLROutputS1xD(222)(1);
  CNStageIntLLRInputS2xD(241)(3) <= VNStageIntLLROutputS1xD(222)(2);
  CNStageIntLLRInputS2xD(376)(3) <= VNStageIntLLROutputS1xD(222)(3);
  CNStageIntLLRInputS2xD(23)(3) <= VNStageIntLLROutputS1xD(223)(0);
  CNStageIntLLRInputS2xD(76)(3) <= VNStageIntLLROutputS1xD(223)(1);
  CNStageIntLLRInputS2xD(162)(3) <= VNStageIntLLROutputS1xD(223)(2);
  CNStageIntLLRInputS2xD(224)(3) <= VNStageIntLLROutputS1xD(223)(3);
  CNStageIntLLRInputS2xD(229)(3) <= VNStageIntLLROutputS1xD(223)(4);
  CNStageIntLLRInputS2xD(309)(3) <= VNStageIntLLROutputS1xD(223)(5);
  CNStageIntLLRInputS2xD(338)(3) <= VNStageIntLLROutputS1xD(223)(6);
  CNStageIntLLRInputS2xD(22)(3) <= VNStageIntLLROutputS1xD(224)(0);
  CNStageIntLLRInputS2xD(90)(3) <= VNStageIntLLROutputS1xD(224)(1);
  CNStageIntLLRInputS2xD(135)(3) <= VNStageIntLLROutputS1xD(224)(2);
  CNStageIntLLRInputS2xD(193)(3) <= VNStageIntLLROutputS1xD(224)(3);
  CNStageIntLLRInputS2xD(270)(3) <= VNStageIntLLROutputS1xD(224)(4);
  CNStageIntLLRInputS2xD(328)(3) <= VNStageIntLLROutputS1xD(224)(5);
  CNStageIntLLRInputS2xD(366)(3) <= VNStageIntLLROutputS1xD(224)(6);
  CNStageIntLLRInputS2xD(21)(3) <= VNStageIntLLROutputS1xD(225)(0);
  CNStageIntLLRInputS2xD(61)(3) <= VNStageIntLLROutputS1xD(225)(1);
  CNStageIntLLRInputS2xD(132)(3) <= VNStageIntLLROutputS1xD(225)(2);
  CNStageIntLLRInputS2xD(188)(3) <= VNStageIntLLROutputS1xD(225)(3);
  CNStageIntLLRInputS2xD(232)(3) <= VNStageIntLLROutputS1xD(225)(4);
  CNStageIntLLRInputS2xD(301)(3) <= VNStageIntLLROutputS1xD(225)(5);
  CNStageIntLLRInputS2xD(20)(3) <= VNStageIntLLROutputS1xD(226)(0);
  CNStageIntLLRInputS2xD(148)(3) <= VNStageIntLLROutputS1xD(226)(1);
  CNStageIntLLRInputS2xD(378)(3) <= VNStageIntLLROutputS1xD(226)(2);
  CNStageIntLLRInputS2xD(19)(3) <= VNStageIntLLROutputS1xD(227)(0);
  CNStageIntLLRInputS2xD(63)(3) <= VNStageIntLLROutputS1xD(227)(1);
  CNStageIntLLRInputS2xD(140)(3) <= VNStageIntLLROutputS1xD(227)(2);
  CNStageIntLLRInputS2xD(178)(3) <= VNStageIntLLROutputS1xD(227)(3);
  CNStageIntLLRInputS2xD(258)(3) <= VNStageIntLLROutputS1xD(227)(4);
  CNStageIntLLRInputS2xD(314)(3) <= VNStageIntLLROutputS1xD(227)(5);
  CNStageIntLLRInputS2xD(368)(3) <= VNStageIntLLROutputS1xD(227)(6);
  CNStageIntLLRInputS2xD(18)(3) <= VNStageIntLLROutputS1xD(228)(0);
  CNStageIntLLRInputS2xD(78)(3) <= VNStageIntLLROutputS1xD(228)(1);
  CNStageIntLLRInputS2xD(114)(3) <= VNStageIntLLROutputS1xD(228)(2);
  CNStageIntLLRInputS2xD(198)(3) <= VNStageIntLLROutputS1xD(228)(3);
  CNStageIntLLRInputS2xD(253)(3) <= VNStageIntLLROutputS1xD(228)(4);
  CNStageIntLLRInputS2xD(307)(3) <= VNStageIntLLROutputS1xD(228)(5);
  CNStageIntLLRInputS2xD(17)(3) <= VNStageIntLLROutputS1xD(229)(0);
  CNStageIntLLRInputS2xD(74)(3) <= VNStageIntLLROutputS1xD(229)(1);
  CNStageIntLLRInputS2xD(124)(3) <= VNStageIntLLROutputS1xD(229)(2);
  CNStageIntLLRInputS2xD(259)(3) <= VNStageIntLLROutputS1xD(229)(3);
  CNStageIntLLRInputS2xD(374)(3) <= VNStageIntLLROutputS1xD(229)(4);
  CNStageIntLLRInputS2xD(16)(3) <= VNStageIntLLROutputS1xD(230)(0);
  CNStageIntLLRInputS2xD(118)(3) <= VNStageIntLLROutputS1xD(230)(1);
  CNStageIntLLRInputS2xD(176)(3) <= VNStageIntLLROutputS1xD(230)(2);
  CNStageIntLLRInputS2xD(249)(3) <= VNStageIntLLROutputS1xD(230)(3);
  CNStageIntLLRInputS2xD(293)(3) <= VNStageIntLLROutputS1xD(230)(4);
  CNStageIntLLRInputS2xD(347)(3) <= VNStageIntLLROutputS1xD(230)(5);
  CNStageIntLLRInputS2xD(15)(3) <= VNStageIntLLROutputS1xD(231)(0);
  CNStageIntLLRInputS2xD(56)(3) <= VNStageIntLLROutputS1xD(231)(1);
  CNStageIntLLRInputS2xD(209)(3) <= VNStageIntLLROutputS1xD(231)(2);
  CNStageIntLLRInputS2xD(272)(3) <= VNStageIntLLROutputS1xD(231)(3);
  CNStageIntLLRInputS2xD(287)(3) <= VNStageIntLLROutputS1xD(231)(4);
  CNStageIntLLRInputS2xD(344)(3) <= VNStageIntLLROutputS1xD(231)(5);
  CNStageIntLLRInputS2xD(14)(3) <= VNStageIntLLROutputS1xD(232)(0);
  CNStageIntLLRInputS2xD(57)(3) <= VNStageIntLLROutputS1xD(232)(1);
  CNStageIntLLRInputS2xD(212)(3) <= VNStageIntLLROutputS1xD(232)(2);
  CNStageIntLLRInputS2xD(278)(3) <= VNStageIntLLROutputS1xD(232)(3);
  CNStageIntLLRInputS2xD(291)(3) <= VNStageIntLLROutputS1xD(232)(4);
  CNStageIntLLRInputS2xD(359)(3) <= VNStageIntLLROutputS1xD(232)(5);
  CNStageIntLLRInputS2xD(13)(3) <= VNStageIntLLROutputS1xD(233)(0);
  CNStageIntLLRInputS2xD(92)(3) <= VNStageIntLLROutputS1xD(233)(1);
  CNStageIntLLRInputS2xD(149)(3) <= VNStageIntLLROutputS1xD(233)(2);
  CNStageIntLLRInputS2xD(263)(3) <= VNStageIntLLROutputS1xD(233)(3);
  CNStageIntLLRInputS2xD(352)(3) <= VNStageIntLLROutputS1xD(233)(4);
  CNStageIntLLRInputS2xD(12)(3) <= VNStageIntLLROutputS1xD(234)(0);
  CNStageIntLLRInputS2xD(84)(3) <= VNStageIntLLROutputS1xD(234)(1);
  CNStageIntLLRInputS2xD(131)(3) <= VNStageIntLLROutputS1xD(234)(2);
  CNStageIntLLRInputS2xD(177)(3) <= VNStageIntLLROutputS1xD(234)(3);
  CNStageIntLLRInputS2xD(265)(3) <= VNStageIntLLROutputS1xD(234)(4);
  CNStageIntLLRInputS2xD(315)(3) <= VNStageIntLLROutputS1xD(234)(5);
  CNStageIntLLRInputS2xD(100)(3) <= VNStageIntLLROutputS1xD(235)(0);
  CNStageIntLLRInputS2xD(144)(3) <= VNStageIntLLROutputS1xD(235)(1);
  CNStageIntLLRInputS2xD(196)(3) <= VNStageIntLLROutputS1xD(235)(2);
  CNStageIntLLRInputS2xD(235)(3) <= VNStageIntLLROutputS1xD(235)(3);
  CNStageIntLLRInputS2xD(336)(3) <= VNStageIntLLROutputS1xD(235)(4);
  CNStageIntLLRInputS2xD(11)(3) <= VNStageIntLLROutputS1xD(236)(0);
  CNStageIntLLRInputS2xD(104)(3) <= VNStageIntLLROutputS1xD(236)(1);
  CNStageIntLLRInputS2xD(155)(3) <= VNStageIntLLROutputS1xD(236)(2);
  CNStageIntLLRInputS2xD(221)(3) <= VNStageIntLLROutputS1xD(236)(3);
  CNStageIntLLRInputS2xD(271)(3) <= VNStageIntLLROutputS1xD(236)(4);
  CNStageIntLLRInputS2xD(310)(3) <= VNStageIntLLROutputS1xD(236)(5);
  CNStageIntLLRInputS2xD(10)(3) <= VNStageIntLLROutputS1xD(237)(0);
  CNStageIntLLRInputS2xD(110)(3) <= VNStageIntLLROutputS1xD(237)(1);
  CNStageIntLLRInputS2xD(125)(3) <= VNStageIntLLROutputS1xD(237)(2);
  CNStageIntLLRInputS2xD(228)(3) <= VNStageIntLLROutputS1xD(237)(3);
  CNStageIntLLRInputS2xD(322)(3) <= VNStageIntLLROutputS1xD(237)(4);
  CNStageIntLLRInputS2xD(334)(3) <= VNStageIntLLROutputS1xD(237)(5);
  CNStageIntLLRInputS2xD(9)(3) <= VNStageIntLLROutputS1xD(238)(0);
  CNStageIntLLRInputS2xD(103)(3) <= VNStageIntLLROutputS1xD(238)(1);
  CNStageIntLLRInputS2xD(113)(3) <= VNStageIntLLROutputS1xD(238)(2);
  CNStageIntLLRInputS2xD(179)(3) <= VNStageIntLLROutputS1xD(238)(3);
  CNStageIntLLRInputS2xD(236)(3) <= VNStageIntLLROutputS1xD(238)(4);
  CNStageIntLLRInputS2xD(294)(3) <= VNStageIntLLROutputS1xD(238)(5);
  CNStageIntLLRInputS2xD(383)(3) <= VNStageIntLLROutputS1xD(238)(6);
  CNStageIntLLRInputS2xD(8)(3) <= VNStageIntLLROutputS1xD(239)(0);
  CNStageIntLLRInputS2xD(98)(3) <= VNStageIntLLROutputS1xD(239)(1);
  CNStageIntLLRInputS2xD(158)(3) <= VNStageIntLLROutputS1xD(239)(2);
  CNStageIntLLRInputS2xD(223)(3) <= VNStageIntLLROutputS1xD(239)(3);
  CNStageIntLLRInputS2xD(264)(3) <= VNStageIntLLROutputS1xD(239)(4);
  CNStageIntLLRInputS2xD(284)(3) <= VNStageIntLLROutputS1xD(239)(5);
  CNStageIntLLRInputS2xD(360)(3) <= VNStageIntLLROutputS1xD(239)(6);
  CNStageIntLLRInputS2xD(7)(3) <= VNStageIntLLROutputS1xD(240)(0);
  CNStageIntLLRInputS2xD(81)(3) <= VNStageIntLLROutputS1xD(240)(1);
  CNStageIntLLRInputS2xD(116)(3) <= VNStageIntLLROutputS1xD(240)(2);
  CNStageIntLLRInputS2xD(210)(3) <= VNStageIntLLROutputS1xD(240)(3);
  CNStageIntLLRInputS2xD(277)(3) <= VNStageIntLLROutputS1xD(240)(4);
  CNStageIntLLRInputS2xD(324)(3) <= VNStageIntLLROutputS1xD(240)(5);
  CNStageIntLLRInputS2xD(343)(3) <= VNStageIntLLROutputS1xD(240)(6);
  CNStageIntLLRInputS2xD(6)(3) <= VNStageIntLLROutputS1xD(241)(0);
  CNStageIntLLRInputS2xD(88)(3) <= VNStageIntLLROutputS1xD(241)(1);
  CNStageIntLLRInputS2xD(175)(3) <= VNStageIntLLROutputS1xD(241)(2);
  CNStageIntLLRInputS2xD(250)(3) <= VNStageIntLLROutputS1xD(241)(3);
  CNStageIntLLRInputS2xD(285)(3) <= VNStageIntLLROutputS1xD(241)(4);
  CNStageIntLLRInputS2xD(355)(3) <= VNStageIntLLROutputS1xD(241)(5);
  CNStageIntLLRInputS2xD(5)(3) <= VNStageIntLLROutputS1xD(242)(0);
  CNStageIntLLRInputS2xD(108)(3) <= VNStageIntLLROutputS1xD(242)(1);
  CNStageIntLLRInputS2xD(146)(3) <= VNStageIntLLROutputS1xD(242)(2);
  CNStageIntLLRInputS2xD(203)(3) <= VNStageIntLLROutputS1xD(242)(3);
  CNStageIntLLRInputS2xD(231)(3) <= VNStageIntLLROutputS1xD(242)(4);
  CNStageIntLLRInputS2xD(303)(3) <= VNStageIntLLROutputS1xD(242)(5);
  CNStageIntLLRInputS2xD(367)(3) <= VNStageIntLLROutputS1xD(242)(6);
  CNStageIntLLRInputS2xD(4)(3) <= VNStageIntLLROutputS1xD(243)(0);
  CNStageIntLLRInputS2xD(106)(3) <= VNStageIntLLROutputS1xD(243)(1);
  CNStageIntLLRInputS2xD(141)(3) <= VNStageIntLLROutputS1xD(243)(2);
  CNStageIntLLRInputS2xD(200)(3) <= VNStageIntLLROutputS1xD(243)(3);
  CNStageIntLLRInputS2xD(252)(3) <= VNStageIntLLROutputS1xD(243)(4);
  CNStageIntLLRInputS2xD(312)(3) <= VNStageIntLLROutputS1xD(243)(5);
  CNStageIntLLRInputS2xD(337)(3) <= VNStageIntLLROutputS1xD(243)(6);
  CNStageIntLLRInputS2xD(147)(3) <= VNStageIntLLROutputS1xD(244)(0);
  CNStageIntLLRInputS2xD(266)(3) <= VNStageIntLLROutputS1xD(244)(1);
  CNStageIntLLRInputS2xD(3)(3) <= VNStageIntLLROutputS1xD(245)(0);
  CNStageIntLLRInputS2xD(66)(3) <= VNStageIntLLROutputS1xD(245)(1);
  CNStageIntLLRInputS2xD(136)(3) <= VNStageIntLLROutputS1xD(245)(2);
  CNStageIntLLRInputS2xD(207)(3) <= VNStageIntLLROutputS1xD(245)(3);
  CNStageIntLLRInputS2xD(262)(3) <= VNStageIntLLROutputS1xD(245)(4);
  CNStageIntLLRInputS2xD(313)(3) <= VNStageIntLLROutputS1xD(245)(5);
  CNStageIntLLRInputS2xD(370)(3) <= VNStageIntLLROutputS1xD(245)(6);
  CNStageIntLLRInputS2xD(2)(3) <= VNStageIntLLROutputS1xD(246)(0);
  CNStageIntLLRInputS2xD(69)(3) <= VNStageIntLLROutputS1xD(246)(1);
  CNStageIntLLRInputS2xD(161)(3) <= VNStageIntLLROutputS1xD(246)(2);
  CNStageIntLLRInputS2xD(185)(3) <= VNStageIntLLROutputS1xD(246)(3);
  CNStageIntLLRInputS2xD(226)(3) <= VNStageIntLLROutputS1xD(246)(4);
  CNStageIntLLRInputS2xD(302)(3) <= VNStageIntLLROutputS1xD(246)(5);
  CNStageIntLLRInputS2xD(1)(3) <= VNStageIntLLROutputS1xD(247)(0);
  CNStageIntLLRInputS2xD(109)(3) <= VNStageIntLLROutputS1xD(247)(1);
  CNStageIntLLRInputS2xD(168)(3) <= VNStageIntLLROutputS1xD(247)(2);
  CNStageIntLLRInputS2xD(194)(3) <= VNStageIntLLROutputS1xD(247)(3);
  CNStageIntLLRInputS2xD(247)(3) <= VNStageIntLLROutputS1xD(247)(4);
  CNStageIntLLRInputS2xD(327)(3) <= VNStageIntLLROutputS1xD(247)(5);
  CNStageIntLLRInputS2xD(349)(3) <= VNStageIntLLROutputS1xD(247)(6);
  CNStageIntLLRInputS2xD(0)(3) <= VNStageIntLLROutputS1xD(248)(0);
  CNStageIntLLRInputS2xD(87)(3) <= VNStageIntLLROutputS1xD(248)(1);
  CNStageIntLLRInputS2xD(151)(3) <= VNStageIntLLROutputS1xD(248)(2);
  CNStageIntLLRInputS2xD(189)(3) <= VNStageIntLLROutputS1xD(248)(3);
  CNStageIntLLRInputS2xD(248)(3) <= VNStageIntLLROutputS1xD(248)(4);
  CNStageIntLLRInputS2xD(280)(3) <= VNStageIntLLROutputS1xD(248)(5);
  CNStageIntLLRInputS2xD(357)(3) <= VNStageIntLLROutputS1xD(248)(6);
  CNStageIntLLRInputS2xD(152)(3) <= VNStageIntLLROutputS1xD(249)(0);
  CNStageIntLLRInputS2xD(192)(3) <= VNStageIntLLROutputS1xD(249)(1);
  CNStageIntLLRInputS2xD(225)(3) <= VNStageIntLLROutputS1xD(249)(2);
  CNStageIntLLRInputS2xD(317)(3) <= VNStageIntLLROutputS1xD(249)(3);
  CNStageIntLLRInputS2xD(353)(3) <= VNStageIntLLROutputS1xD(249)(4);
  CNStageIntLLRInputS2xD(79)(3) <= VNStageIntLLROutputS1xD(250)(0);
  CNStageIntLLRInputS2xD(120)(3) <= VNStageIntLLROutputS1xD(250)(1);
  CNStageIntLLRInputS2xD(184)(3) <= VNStageIntLLROutputS1xD(250)(2);
  CNStageIntLLRInputS2xD(319)(3) <= VNStageIntLLROutputS1xD(250)(3);
  CNStageIntLLRInputS2xD(358)(3) <= VNStageIntLLROutputS1xD(250)(4);
  CNStageIntLLRInputS2xD(62)(3) <= VNStageIntLLROutputS1xD(251)(0);
  CNStageIntLLRInputS2xD(159)(3) <= VNStageIntLLROutputS1xD(251)(1);
  CNStageIntLLRInputS2xD(215)(3) <= VNStageIntLLROutputS1xD(251)(2);
  CNStageIntLLRInputS2xD(289)(3) <= VNStageIntLLROutputS1xD(251)(3);
  CNStageIntLLRInputS2xD(348)(3) <= VNStageIntLLROutputS1xD(251)(4);
  CNStageIntLLRInputS2xD(89)(3) <= VNStageIntLLROutputS1xD(252)(0);
  CNStageIntLLRInputS2xD(112)(3) <= VNStageIntLLROutputS1xD(252)(1);
  CNStageIntLLRInputS2xD(199)(3) <= VNStageIntLLROutputS1xD(252)(2);
  CNStageIntLLRInputS2xD(239)(3) <= VNStageIntLLROutputS1xD(252)(3);
  CNStageIntLLRInputS2xD(325)(3) <= VNStageIntLLROutputS1xD(252)(4);
  CNStageIntLLRInputS2xD(373)(3) <= VNStageIntLLROutputS1xD(252)(5);
  CNStageIntLLRInputS2xD(80)(3) <= VNStageIntLLROutputS1xD(253)(0);
  CNStageIntLLRInputS2xD(121)(3) <= VNStageIntLLROutputS1xD(253)(1);
  CNStageIntLLRInputS2xD(211)(3) <= VNStageIntLLROutputS1xD(253)(2);
  CNStageIntLLRInputS2xD(279)(3) <= VNStageIntLLROutputS1xD(253)(3);
  CNStageIntLLRInputS2xD(283)(3) <= VNStageIntLLROutputS1xD(253)(4);
  CNStageIntLLRInputS2xD(380)(3) <= VNStageIntLLROutputS1xD(253)(5);
  CNStageIntLLRInputS2xD(67)(3) <= VNStageIntLLROutputS1xD(254)(0);
  CNStageIntLLRInputS2xD(222)(3) <= VNStageIntLLROutputS1xD(254)(1);
  CNStageIntLLRInputS2xD(238)(3) <= VNStageIntLLROutputS1xD(254)(2);
  CNStageIntLLRInputS2xD(290)(3) <= VNStageIntLLROutputS1xD(254)(3);
  CNStageIntLLRInputS2xD(362)(3) <= VNStageIntLLROutputS1xD(254)(4);
  CNStageIntLLRInputS2xD(52)(3) <= VNStageIntLLROutputS1xD(255)(0);
  CNStageIntLLRInputS2xD(86)(3) <= VNStageIntLLROutputS1xD(255)(1);
  CNStageIntLLRInputS2xD(167)(3) <= VNStageIntLLROutputS1xD(255)(2);
  CNStageIntLLRInputS2xD(195)(3) <= VNStageIntLLROutputS1xD(255)(3);
  CNStageIntLLRInputS2xD(233)(3) <= VNStageIntLLROutputS1xD(255)(4);
  CNStageIntLLRInputS2xD(318)(3) <= VNStageIntLLROutputS1xD(255)(5);
  CNStageIntLLRInputS2xD(364)(3) <= VNStageIntLLROutputS1xD(255)(6);
  CNStageIntLLRInputS2xD(53)(4) <= VNStageIntLLROutputS1xD(256)(0);
  CNStageIntLLRInputS2xD(106)(4) <= VNStageIntLLROutputS1xD(256)(1);
  CNStageIntLLRInputS2xD(127)(4) <= VNStageIntLLROutputS1xD(256)(2);
  CNStageIntLLRInputS2xD(242)(4) <= VNStageIntLLROutputS1xD(256)(3);
  CNStageIntLLRInputS2xD(296)(4) <= VNStageIntLLROutputS1xD(256)(4);
  CNStageIntLLRInputS2xD(339)(4) <= VNStageIntLLROutputS1xD(256)(5);
  CNStageIntLLRInputS2xD(51)(4) <= VNStageIntLLROutputS1xD(257)(0);
  CNStageIntLLRInputS2xD(85)(4) <= VNStageIntLLROutputS1xD(257)(1);
  CNStageIntLLRInputS2xD(166)(4) <= VNStageIntLLROutputS1xD(257)(2);
  CNStageIntLLRInputS2xD(194)(4) <= VNStageIntLLROutputS1xD(257)(3);
  CNStageIntLLRInputS2xD(232)(4) <= VNStageIntLLROutputS1xD(257)(4);
  CNStageIntLLRInputS2xD(317)(4) <= VNStageIntLLROutputS1xD(257)(5);
  CNStageIntLLRInputS2xD(363)(4) <= VNStageIntLLROutputS1xD(257)(6);
  CNStageIntLLRInputS2xD(50)(4) <= VNStageIntLLROutputS1xD(258)(0);
  CNStageIntLLRInputS2xD(57)(4) <= VNStageIntLLROutputS1xD(258)(1);
  CNStageIntLLRInputS2xD(331)(4) <= VNStageIntLLROutputS1xD(258)(2);
  CNStageIntLLRInputS2xD(54)(4) <= VNStageIntLLROutputS1xD(259)(0);
  CNStageIntLLRInputS2xD(114)(4) <= VNStageIntLLROutputS1xD(259)(1);
  CNStageIntLLRInputS2xD(274)(4) <= VNStageIntLLROutputS1xD(259)(2);
  CNStageIntLLRInputS2xD(303)(4) <= VNStageIntLLROutputS1xD(259)(3);
  CNStageIntLLRInputS2xD(370)(4) <= VNStageIntLLROutputS1xD(259)(4);
  CNStageIntLLRInputS2xD(49)(4) <= VNStageIntLLROutputS1xD(260)(0);
  CNStageIntLLRInputS2xD(71)(4) <= VNStageIntLLROutputS1xD(260)(1);
  CNStageIntLLRInputS2xD(138)(4) <= VNStageIntLLROutputS1xD(260)(2);
  CNStageIntLLRInputS2xD(186)(4) <= VNStageIntLLROutputS1xD(260)(3);
  CNStageIntLLRInputS2xD(243)(4) <= VNStageIntLLROutputS1xD(260)(4);
  CNStageIntLLRInputS2xD(383)(4) <= VNStageIntLLROutputS1xD(260)(5);
  CNStageIntLLRInputS2xD(48)(4) <= VNStageIntLLROutputS1xD(261)(0);
  CNStageIntLLRInputS2xD(63)(4) <= VNStageIntLLROutputS1xD(261)(1);
  CNStageIntLLRInputS2xD(152)(4) <= VNStageIntLLROutputS1xD(261)(2);
  CNStageIntLLRInputS2xD(204)(4) <= VNStageIntLLROutputS1xD(261)(3);
  CNStageIntLLRInputS2xD(305)(4) <= VNStageIntLLROutputS1xD(261)(4);
  CNStageIntLLRInputS2xD(333)(4) <= VNStageIntLLROutputS1xD(261)(5);
  CNStageIntLLRInputS2xD(47)(4) <= VNStageIntLLROutputS1xD(262)(0);
  CNStageIntLLRInputS2xD(95)(4) <= VNStageIntLLROutputS1xD(262)(1);
  CNStageIntLLRInputS2xD(149)(4) <= VNStageIntLLROutputS1xD(262)(2);
  CNStageIntLLRInputS2xD(212)(4) <= VNStageIntLLROutputS1xD(262)(3);
  CNStageIntLLRInputS2xD(319)(4) <= VNStageIntLLROutputS1xD(262)(4);
  CNStageIntLLRInputS2xD(362)(4) <= VNStageIntLLROutputS1xD(262)(5);
  CNStageIntLLRInputS2xD(46)(4) <= VNStageIntLLROutputS1xD(263)(0);
  CNStageIntLLRInputS2xD(104)(4) <= VNStageIntLLROutputS1xD(263)(1);
  CNStageIntLLRInputS2xD(169)(4) <= VNStageIntLLROutputS1xD(263)(2);
  CNStageIntLLRInputS2xD(207)(4) <= VNStageIntLLROutputS1xD(263)(3);
  CNStageIntLLRInputS2xD(253)(4) <= VNStageIntLLROutputS1xD(263)(4);
  CNStageIntLLRInputS2xD(315)(4) <= VNStageIntLLROutputS1xD(263)(5);
  CNStageIntLLRInputS2xD(378)(4) <= VNStageIntLLROutputS1xD(263)(6);
  CNStageIntLLRInputS2xD(45)(4) <= VNStageIntLLROutputS1xD(264)(0);
  CNStageIntLLRInputS2xD(98)(4) <= VNStageIntLLROutputS1xD(264)(1);
  CNStageIntLLRInputS2xD(132)(4) <= VNStageIntLLROutputS1xD(264)(2);
  CNStageIntLLRInputS2xD(213)(4) <= VNStageIntLLROutputS1xD(264)(3);
  CNStageIntLLRInputS2xD(256)(4) <= VNStageIntLLROutputS1xD(264)(4);
  CNStageIntLLRInputS2xD(281)(4) <= VNStageIntLLROutputS1xD(264)(5);
  CNStageIntLLRInputS2xD(349)(4) <= VNStageIntLLROutputS1xD(264)(6);
  CNStageIntLLRInputS2xD(44)(4) <= VNStageIntLLROutputS1xD(265)(0);
  CNStageIntLLRInputS2xD(133)(4) <= VNStageIntLLROutputS1xD(265)(1);
  CNStageIntLLRInputS2xD(203)(4) <= VNStageIntLLROutputS1xD(265)(2);
  CNStageIntLLRInputS2xD(244)(4) <= VNStageIntLLROutputS1xD(265)(3);
  CNStageIntLLRInputS2xD(43)(4) <= VNStageIntLLROutputS1xD(266)(0);
  CNStageIntLLRInputS2xD(168)(4) <= VNStageIntLLROutputS1xD(266)(1);
  CNStageIntLLRInputS2xD(173)(4) <= VNStageIntLLROutputS1xD(266)(2);
  CNStageIntLLRInputS2xD(273)(4) <= VNStageIntLLROutputS1xD(266)(3);
  CNStageIntLLRInputS2xD(300)(4) <= VNStageIntLLROutputS1xD(266)(4);
  CNStageIntLLRInputS2xD(42)(4) <= VNStageIntLLROutputS1xD(267)(0);
  CNStageIntLLRInputS2xD(72)(4) <= VNStageIntLLROutputS1xD(267)(1);
  CNStageIntLLRInputS2xD(159)(4) <= VNStageIntLLROutputS1xD(267)(2);
  CNStageIntLLRInputS2xD(180)(4) <= VNStageIntLLROutputS1xD(267)(3);
  CNStageIntLLRInputS2xD(241)(4) <= VNStageIntLLROutputS1xD(267)(4);
  CNStageIntLLRInputS2xD(280)(4) <= VNStageIntLLROutputS1xD(267)(5);
  CNStageIntLLRInputS2xD(364)(4) <= VNStageIntLLROutputS1xD(267)(6);
  CNStageIntLLRInputS2xD(41)(4) <= VNStageIntLLROutputS1xD(268)(0);
  CNStageIntLLRInputS2xD(109)(4) <= VNStageIntLLROutputS1xD(268)(1);
  CNStageIntLLRInputS2xD(118)(4) <= VNStageIntLLROutputS1xD(268)(2);
  CNStageIntLLRInputS2xD(216)(4) <= VNStageIntLLROutputS1xD(268)(3);
  CNStageIntLLRInputS2xD(266)(4) <= VNStageIntLLROutputS1xD(268)(4);
  CNStageIntLLRInputS2xD(325)(4) <= VNStageIntLLROutputS1xD(268)(5);
  CNStageIntLLRInputS2xD(360)(4) <= VNStageIntLLROutputS1xD(268)(6);
  CNStageIntLLRInputS2xD(67)(4) <= VNStageIntLLROutputS1xD(269)(0);
  CNStageIntLLRInputS2xD(122)(4) <= VNStageIntLLROutputS1xD(269)(1);
  CNStageIntLLRInputS2xD(218)(4) <= VNStageIntLLROutputS1xD(269)(2);
  CNStageIntLLRInputS2xD(250)(4) <= VNStageIntLLROutputS1xD(269)(3);
  CNStageIntLLRInputS2xD(287)(4) <= VNStageIntLLROutputS1xD(269)(4);
  CNStageIntLLRInputS2xD(381)(4) <= VNStageIntLLROutputS1xD(269)(5);
  CNStageIntLLRInputS2xD(40)(4) <= VNStageIntLLROutputS1xD(270)(0);
  CNStageIntLLRInputS2xD(79)(4) <= VNStageIntLLROutputS1xD(270)(1);
  CNStageIntLLRInputS2xD(170)(4) <= VNStageIntLLROutputS1xD(270)(2);
  CNStageIntLLRInputS2xD(190)(4) <= VNStageIntLLROutputS1xD(270)(3);
  CNStageIntLLRInputS2xD(275)(4) <= VNStageIntLLROutputS1xD(270)(4);
  CNStageIntLLRInputS2xD(292)(4) <= VNStageIntLLROutputS1xD(270)(5);
  CNStageIntLLRInputS2xD(344)(4) <= VNStageIntLLROutputS1xD(270)(6);
  CNStageIntLLRInputS2xD(39)(4) <= VNStageIntLLROutputS1xD(271)(0);
  CNStageIntLLRInputS2xD(105)(4) <= VNStageIntLLROutputS1xD(271)(1);
  CNStageIntLLRInputS2xD(171)(4) <= VNStageIntLLROutputS1xD(271)(2);
  CNStageIntLLRInputS2xD(268)(4) <= VNStageIntLLROutputS1xD(271)(3);
  CNStageIntLLRInputS2xD(332)(4) <= VNStageIntLLROutputS1xD(271)(4);
  CNStageIntLLRInputS2xD(345)(4) <= VNStageIntLLROutputS1xD(271)(5);
  CNStageIntLLRInputS2xD(38)(4) <= VNStageIntLLROutputS1xD(272)(0);
  CNStageIntLLRInputS2xD(94)(4) <= VNStageIntLLROutputS1xD(272)(1);
  CNStageIntLLRInputS2xD(116)(4) <= VNStageIntLLROutputS1xD(272)(2);
  CNStageIntLLRInputS2xD(184)(4) <= VNStageIntLLROutputS1xD(272)(3);
  CNStageIntLLRInputS2xD(254)(4) <= VNStageIntLLROutputS1xD(272)(4);
  CNStageIntLLRInputS2xD(291)(4) <= VNStageIntLLROutputS1xD(272)(5);
  CNStageIntLLRInputS2xD(380)(4) <= VNStageIntLLROutputS1xD(272)(6);
  CNStageIntLLRInputS2xD(37)(4) <= VNStageIntLLROutputS1xD(273)(0);
  CNStageIntLLRInputS2xD(81)(4) <= VNStageIntLLROutputS1xD(273)(1);
  CNStageIntLLRInputS2xD(156)(4) <= VNStageIntLLROutputS1xD(273)(2);
  CNStageIntLLRInputS2xD(272)(4) <= VNStageIntLLROutputS1xD(273)(3);
  CNStageIntLLRInputS2xD(285)(4) <= VNStageIntLLROutputS1xD(273)(4);
  CNStageIntLLRInputS2xD(371)(4) <= VNStageIntLLROutputS1xD(273)(5);
  CNStageIntLLRInputS2xD(36)(4) <= VNStageIntLLROutputS1xD(274)(0);
  CNStageIntLLRInputS2xD(164)(4) <= VNStageIntLLROutputS1xD(274)(1);
  CNStageIntLLRInputS2xD(217)(4) <= VNStageIntLLROutputS1xD(274)(2);
  CNStageIntLLRInputS2xD(248)(4) <= VNStageIntLLROutputS1xD(274)(3);
  CNStageIntLLRInputS2xD(35)(4) <= VNStageIntLLROutputS1xD(275)(0);
  CNStageIntLLRInputS2xD(59)(4) <= VNStageIntLLROutputS1xD(275)(1);
  CNStageIntLLRInputS2xD(128)(4) <= VNStageIntLLROutputS1xD(275)(2);
  CNStageIntLLRInputS2xD(179)(4) <= VNStageIntLLROutputS1xD(275)(3);
  CNStageIntLLRInputS2xD(329)(4) <= VNStageIntLLROutputS1xD(275)(4);
  CNStageIntLLRInputS2xD(34)(4) <= VNStageIntLLROutputS1xD(276)(0);
  CNStageIntLLRInputS2xD(69)(4) <= VNStageIntLLROutputS1xD(276)(1);
  CNStageIntLLRInputS2xD(126)(4) <= VNStageIntLLROutputS1xD(276)(2);
  CNStageIntLLRInputS2xD(205)(4) <= VNStageIntLLROutputS1xD(276)(3);
  CNStageIntLLRInputS2xD(259)(4) <= VNStageIntLLROutputS1xD(276)(4);
  CNStageIntLLRInputS2xD(297)(4) <= VNStageIntLLROutputS1xD(276)(5);
  CNStageIntLLRInputS2xD(33)(4) <= VNStageIntLLROutputS1xD(277)(0);
  CNStageIntLLRInputS2xD(64)(4) <= VNStageIntLLROutputS1xD(277)(1);
  CNStageIntLLRInputS2xD(162)(4) <= VNStageIntLLROutputS1xD(277)(2);
  CNStageIntLLRInputS2xD(185)(4) <= VNStageIntLLROutputS1xD(277)(3);
  CNStageIntLLRInputS2xD(252)(4) <= VNStageIntLLROutputS1xD(277)(4);
  CNStageIntLLRInputS2xD(295)(4) <= VNStageIntLLROutputS1xD(277)(5);
  CNStageIntLLRInputS2xD(334)(4) <= VNStageIntLLROutputS1xD(277)(6);
  CNStageIntLLRInputS2xD(32)(4) <= VNStageIntLLROutputS1xD(278)(0);
  CNStageIntLLRInputS2xD(70)(4) <= VNStageIntLLROutputS1xD(278)(1);
  CNStageIntLLRInputS2xD(141)(4) <= VNStageIntLLROutputS1xD(278)(2);
  CNStageIntLLRInputS2xD(229)(4) <= VNStageIntLLROutputS1xD(278)(3);
  CNStageIntLLRInputS2xD(328)(4) <= VNStageIntLLROutputS1xD(278)(4);
  CNStageIntLLRInputS2xD(31)(4) <= VNStageIntLLROutputS1xD(279)(0);
  CNStageIntLLRInputS2xD(58)(4) <= VNStageIntLLROutputS1xD(279)(1);
  CNStageIntLLRInputS2xD(144)(4) <= VNStageIntLLROutputS1xD(279)(2);
  CNStageIntLLRInputS2xD(219)(4) <= VNStageIntLLROutputS1xD(279)(3);
  CNStageIntLLRInputS2xD(239)(4) <= VNStageIntLLROutputS1xD(279)(4);
  CNStageIntLLRInputS2xD(368)(4) <= VNStageIntLLROutputS1xD(279)(5);
  CNStageIntLLRInputS2xD(30)(4) <= VNStageIntLLROutputS1xD(280)(0);
  CNStageIntLLRInputS2xD(84)(4) <= VNStageIntLLROutputS1xD(280)(1);
  CNStageIntLLRInputS2xD(129)(4) <= VNStageIntLLROutputS1xD(280)(2);
  CNStageIntLLRInputS2xD(215)(4) <= VNStageIntLLROutputS1xD(280)(3);
  CNStageIntLLRInputS2xD(233)(4) <= VNStageIntLLROutputS1xD(280)(4);
  CNStageIntLLRInputS2xD(310)(4) <= VNStageIntLLROutputS1xD(280)(5);
  CNStageIntLLRInputS2xD(376)(4) <= VNStageIntLLROutputS1xD(280)(6);
  CNStageIntLLRInputS2xD(29)(4) <= VNStageIntLLROutputS1xD(281)(0);
  CNStageIntLLRInputS2xD(90)(4) <= VNStageIntLLROutputS1xD(281)(1);
  CNStageIntLLRInputS2xD(163)(4) <= VNStageIntLLROutputS1xD(281)(2);
  CNStageIntLLRInputS2xD(182)(4) <= VNStageIntLLROutputS1xD(281)(3);
  CNStageIntLLRInputS2xD(236)(4) <= VNStageIntLLROutputS1xD(281)(4);
  CNStageIntLLRInputS2xD(298)(4) <= VNStageIntLLROutputS1xD(281)(5);
  CNStageIntLLRInputS2xD(340)(4) <= VNStageIntLLROutputS1xD(281)(6);
  CNStageIntLLRInputS2xD(28)(4) <= VNStageIntLLROutputS1xD(282)(0);
  CNStageIntLLRInputS2xD(74)(4) <= VNStageIntLLROutputS1xD(282)(1);
  CNStageIntLLRInputS2xD(125)(4) <= VNStageIntLLROutputS1xD(282)(2);
  CNStageIntLLRInputS2xD(200)(4) <= VNStageIntLLROutputS1xD(282)(3);
  CNStageIntLLRInputS2xD(226)(4) <= VNStageIntLLROutputS1xD(282)(4);
  CNStageIntLLRInputS2xD(338)(4) <= VNStageIntLLROutputS1xD(282)(5);
  CNStageIntLLRInputS2xD(27)(4) <= VNStageIntLLROutputS1xD(283)(0);
  CNStageIntLLRInputS2xD(76)(4) <= VNStageIntLLROutputS1xD(283)(1);
  CNStageIntLLRInputS2xD(153)(4) <= VNStageIntLLROutputS1xD(283)(2);
  CNStageIntLLRInputS2xD(201)(4) <= VNStageIntLLROutputS1xD(283)(3);
  CNStageIntLLRInputS2xD(260)(4) <= VNStageIntLLROutputS1xD(283)(4);
  CNStageIntLLRInputS2xD(294)(4) <= VNStageIntLLROutputS1xD(283)(5);
  CNStageIntLLRInputS2xD(374)(4) <= VNStageIntLLROutputS1xD(283)(6);
  CNStageIntLLRInputS2xD(26)(4) <= VNStageIntLLROutputS1xD(284)(0);
  CNStageIntLLRInputS2xD(100)(4) <= VNStageIntLLROutputS1xD(284)(1);
  CNStageIntLLRInputS2xD(137)(4) <= VNStageIntLLROutputS1xD(284)(2);
  CNStageIntLLRInputS2xD(181)(4) <= VNStageIntLLROutputS1xD(284)(3);
  CNStageIntLLRInputS2xD(245)(4) <= VNStageIntLLROutputS1xD(284)(4);
  CNStageIntLLRInputS2xD(320)(4) <= VNStageIntLLROutputS1xD(284)(5);
  CNStageIntLLRInputS2xD(353)(4) <= VNStageIntLLROutputS1xD(284)(6);
  CNStageIntLLRInputS2xD(25)(4) <= VNStageIntLLROutputS1xD(285)(0);
  CNStageIntLLRInputS2xD(82)(4) <= VNStageIntLLROutputS1xD(285)(1);
  CNStageIntLLRInputS2xD(165)(4) <= VNStageIntLLROutputS1xD(285)(2);
  CNStageIntLLRInputS2xD(172)(4) <= VNStageIntLLROutputS1xD(285)(3);
  CNStageIntLLRInputS2xD(255)(4) <= VNStageIntLLROutputS1xD(285)(4);
  CNStageIntLLRInputS2xD(304)(4) <= VNStageIntLLROutputS1xD(285)(5);
  CNStageIntLLRInputS2xD(355)(4) <= VNStageIntLLROutputS1xD(285)(6);
  CNStageIntLLRInputS2xD(24)(4) <= VNStageIntLLROutputS1xD(286)(0);
  CNStageIntLLRInputS2xD(93)(4) <= VNStageIntLLROutputS1xD(286)(1);
  CNStageIntLLRInputS2xD(155)(4) <= VNStageIntLLROutputS1xD(286)(2);
  CNStageIntLLRInputS2xD(189)(4) <= VNStageIntLLROutputS1xD(286)(3);
  CNStageIntLLRInputS2xD(267)(4) <= VNStageIntLLROutputS1xD(286)(4);
  CNStageIntLLRInputS2xD(330)(4) <= VNStageIntLLROutputS1xD(286)(5);
  CNStageIntLLRInputS2xD(341)(4) <= VNStageIntLLROutputS1xD(286)(6);
  CNStageIntLLRInputS2xD(23)(4) <= VNStageIntLLROutputS1xD(287)(0);
  CNStageIntLLRInputS2xD(101)(4) <= VNStageIntLLROutputS1xD(287)(1);
  CNStageIntLLRInputS2xD(142)(4) <= VNStageIntLLROutputS1xD(287)(2);
  CNStageIntLLRInputS2xD(193)(4) <= VNStageIntLLROutputS1xD(287)(3);
  CNStageIntLLRInputS2xD(240)(4) <= VNStageIntLLROutputS1xD(287)(4);
  CNStageIntLLRInputS2xD(322)(4) <= VNStageIntLLROutputS1xD(287)(5);
  CNStageIntLLRInputS2xD(375)(4) <= VNStageIntLLROutputS1xD(287)(6);
  CNStageIntLLRInputS2xD(22)(4) <= VNStageIntLLROutputS1xD(288)(0);
  CNStageIntLLRInputS2xD(75)(4) <= VNStageIntLLROutputS1xD(288)(1);
  CNStageIntLLRInputS2xD(161)(4) <= VNStageIntLLROutputS1xD(288)(2);
  CNStageIntLLRInputS2xD(224)(4) <= VNStageIntLLROutputS1xD(288)(3);
  CNStageIntLLRInputS2xD(228)(4) <= VNStageIntLLROutputS1xD(288)(4);
  CNStageIntLLRInputS2xD(308)(4) <= VNStageIntLLROutputS1xD(288)(5);
  CNStageIntLLRInputS2xD(337)(4) <= VNStageIntLLROutputS1xD(288)(6);
  CNStageIntLLRInputS2xD(21)(4) <= VNStageIntLLROutputS1xD(289)(0);
  CNStageIntLLRInputS2xD(89)(4) <= VNStageIntLLROutputS1xD(289)(1);
  CNStageIntLLRInputS2xD(134)(4) <= VNStageIntLLROutputS1xD(289)(2);
  CNStageIntLLRInputS2xD(192)(4) <= VNStageIntLLROutputS1xD(289)(3);
  CNStageIntLLRInputS2xD(269)(4) <= VNStageIntLLROutputS1xD(289)(4);
  CNStageIntLLRInputS2xD(327)(4) <= VNStageIntLLROutputS1xD(289)(5);
  CNStageIntLLRInputS2xD(365)(4) <= VNStageIntLLROutputS1xD(289)(6);
  CNStageIntLLRInputS2xD(20)(4) <= VNStageIntLLROutputS1xD(290)(0);
  CNStageIntLLRInputS2xD(60)(4) <= VNStageIntLLROutputS1xD(290)(1);
  CNStageIntLLRInputS2xD(131)(4) <= VNStageIntLLROutputS1xD(290)(2);
  CNStageIntLLRInputS2xD(187)(4) <= VNStageIntLLROutputS1xD(290)(3);
  CNStageIntLLRInputS2xD(231)(4) <= VNStageIntLLROutputS1xD(290)(4);
  CNStageIntLLRInputS2xD(350)(4) <= VNStageIntLLROutputS1xD(290)(5);
  CNStageIntLLRInputS2xD(19)(4) <= VNStageIntLLROutputS1xD(291)(0);
  CNStageIntLLRInputS2xD(96)(4) <= VNStageIntLLROutputS1xD(291)(1);
  CNStageIntLLRInputS2xD(147)(4) <= VNStageIntLLROutputS1xD(291)(2);
  CNStageIntLLRInputS2xD(223)(4) <= VNStageIntLLROutputS1xD(291)(3);
  CNStageIntLLRInputS2xD(249)(4) <= VNStageIntLLROutputS1xD(291)(4);
  CNStageIntLLRInputS2xD(377)(4) <= VNStageIntLLROutputS1xD(291)(5);
  CNStageIntLLRInputS2xD(18)(4) <= VNStageIntLLROutputS1xD(292)(0);
  CNStageIntLLRInputS2xD(62)(4) <= VNStageIntLLROutputS1xD(292)(1);
  CNStageIntLLRInputS2xD(139)(4) <= VNStageIntLLROutputS1xD(292)(2);
  CNStageIntLLRInputS2xD(177)(4) <= VNStageIntLLROutputS1xD(292)(3);
  CNStageIntLLRInputS2xD(257)(4) <= VNStageIntLLROutputS1xD(292)(4);
  CNStageIntLLRInputS2xD(313)(4) <= VNStageIntLLROutputS1xD(292)(5);
  CNStageIntLLRInputS2xD(367)(4) <= VNStageIntLLROutputS1xD(292)(6);
  CNStageIntLLRInputS2xD(17)(4) <= VNStageIntLLROutputS1xD(293)(0);
  CNStageIntLLRInputS2xD(77)(4) <= VNStageIntLLROutputS1xD(293)(1);
  CNStageIntLLRInputS2xD(113)(4) <= VNStageIntLLROutputS1xD(293)(2);
  CNStageIntLLRInputS2xD(197)(4) <= VNStageIntLLROutputS1xD(293)(3);
  CNStageIntLLRInputS2xD(306)(4) <= VNStageIntLLROutputS1xD(293)(4);
  CNStageIntLLRInputS2xD(354)(4) <= VNStageIntLLROutputS1xD(293)(5);
  CNStageIntLLRInputS2xD(16)(4) <= VNStageIntLLROutputS1xD(294)(0);
  CNStageIntLLRInputS2xD(73)(4) <= VNStageIntLLROutputS1xD(294)(1);
  CNStageIntLLRInputS2xD(123)(4) <= VNStageIntLLROutputS1xD(294)(2);
  CNStageIntLLRInputS2xD(196)(4) <= VNStageIntLLROutputS1xD(294)(3);
  CNStageIntLLRInputS2xD(258)(4) <= VNStageIntLLROutputS1xD(294)(4);
  CNStageIntLLRInputS2xD(284)(4) <= VNStageIntLLROutputS1xD(294)(5);
  CNStageIntLLRInputS2xD(373)(4) <= VNStageIntLLROutputS1xD(294)(6);
  CNStageIntLLRInputS2xD(15)(4) <= VNStageIntLLROutputS1xD(295)(0);
  CNStageIntLLRInputS2xD(92)(4) <= VNStageIntLLROutputS1xD(295)(1);
  CNStageIntLLRInputS2xD(117)(4) <= VNStageIntLLROutputS1xD(295)(2);
  CNStageIntLLRInputS2xD(175)(4) <= VNStageIntLLROutputS1xD(295)(3);
  CNStageIntLLRInputS2xD(346)(4) <= VNStageIntLLROutputS1xD(295)(4);
  CNStageIntLLRInputS2xD(14)(4) <= VNStageIntLLROutputS1xD(296)(0);
  CNStageIntLLRInputS2xD(55)(4) <= VNStageIntLLROutputS1xD(296)(1);
  CNStageIntLLRInputS2xD(121)(4) <= VNStageIntLLROutputS1xD(296)(2);
  CNStageIntLLRInputS2xD(208)(4) <= VNStageIntLLROutputS1xD(296)(3);
  CNStageIntLLRInputS2xD(286)(4) <= VNStageIntLLROutputS1xD(296)(4);
  CNStageIntLLRInputS2xD(343)(4) <= VNStageIntLLROutputS1xD(296)(5);
  CNStageIntLLRInputS2xD(13)(4) <= VNStageIntLLROutputS1xD(297)(0);
  CNStageIntLLRInputS2xD(56)(4) <= VNStageIntLLROutputS1xD(297)(1);
  CNStageIntLLRInputS2xD(111)(4) <= VNStageIntLLROutputS1xD(297)(2);
  CNStageIntLLRInputS2xD(211)(4) <= VNStageIntLLROutputS1xD(297)(3);
  CNStageIntLLRInputS2xD(277)(4) <= VNStageIntLLROutputS1xD(297)(4);
  CNStageIntLLRInputS2xD(290)(4) <= VNStageIntLLROutputS1xD(297)(5);
  CNStageIntLLRInputS2xD(358)(4) <= VNStageIntLLROutputS1xD(297)(6);
  CNStageIntLLRInputS2xD(12)(4) <= VNStageIntLLROutputS1xD(298)(0);
  CNStageIntLLRInputS2xD(91)(4) <= VNStageIntLLROutputS1xD(298)(1);
  CNStageIntLLRInputS2xD(148)(4) <= VNStageIntLLROutputS1xD(298)(2);
  CNStageIntLLRInputS2xD(198)(4) <= VNStageIntLLROutputS1xD(298)(3);
  CNStageIntLLRInputS2xD(262)(4) <= VNStageIntLLROutputS1xD(298)(4);
  CNStageIntLLRInputS2xD(282)(4) <= VNStageIntLLROutputS1xD(298)(5);
  CNStageIntLLRInputS2xD(351)(4) <= VNStageIntLLROutputS1xD(298)(6);
  CNStageIntLLRInputS2xD(83)(4) <= VNStageIntLLROutputS1xD(299)(0);
  CNStageIntLLRInputS2xD(130)(4) <= VNStageIntLLROutputS1xD(299)(1);
  CNStageIntLLRInputS2xD(176)(4) <= VNStageIntLLROutputS1xD(299)(2);
  CNStageIntLLRInputS2xD(264)(4) <= VNStageIntLLROutputS1xD(299)(3);
  CNStageIntLLRInputS2xD(314)(4) <= VNStageIntLLROutputS1xD(299)(4);
  CNStageIntLLRInputS2xD(11)(4) <= VNStageIntLLROutputS1xD(300)(0);
  CNStageIntLLRInputS2xD(99)(4) <= VNStageIntLLROutputS1xD(300)(1);
  CNStageIntLLRInputS2xD(143)(4) <= VNStageIntLLROutputS1xD(300)(2);
  CNStageIntLLRInputS2xD(195)(4) <= VNStageIntLLROutputS1xD(300)(3);
  CNStageIntLLRInputS2xD(299)(4) <= VNStageIntLLROutputS1xD(300)(4);
  CNStageIntLLRInputS2xD(335)(4) <= VNStageIntLLROutputS1xD(300)(5);
  CNStageIntLLRInputS2xD(10)(4) <= VNStageIntLLROutputS1xD(301)(0);
  CNStageIntLLRInputS2xD(103)(4) <= VNStageIntLLROutputS1xD(301)(1);
  CNStageIntLLRInputS2xD(154)(4) <= VNStageIntLLROutputS1xD(301)(2);
  CNStageIntLLRInputS2xD(220)(4) <= VNStageIntLLROutputS1xD(301)(3);
  CNStageIntLLRInputS2xD(270)(4) <= VNStageIntLLROutputS1xD(301)(4);
  CNStageIntLLRInputS2xD(309)(4) <= VNStageIntLLROutputS1xD(301)(5);
  CNStageIntLLRInputS2xD(9)(4) <= VNStageIntLLROutputS1xD(302)(0);
  CNStageIntLLRInputS2xD(110)(4) <= VNStageIntLLROutputS1xD(302)(1);
  CNStageIntLLRInputS2xD(124)(4) <= VNStageIntLLROutputS1xD(302)(2);
  CNStageIntLLRInputS2xD(206)(4) <= VNStageIntLLROutputS1xD(302)(3);
  CNStageIntLLRInputS2xD(227)(4) <= VNStageIntLLROutputS1xD(302)(4);
  CNStageIntLLRInputS2xD(321)(4) <= VNStageIntLLROutputS1xD(302)(5);
  CNStageIntLLRInputS2xD(8)(4) <= VNStageIntLLROutputS1xD(303)(0);
  CNStageIntLLRInputS2xD(102)(4) <= VNStageIntLLROutputS1xD(303)(1);
  CNStageIntLLRInputS2xD(112)(4) <= VNStageIntLLROutputS1xD(303)(2);
  CNStageIntLLRInputS2xD(178)(4) <= VNStageIntLLROutputS1xD(303)(3);
  CNStageIntLLRInputS2xD(235)(4) <= VNStageIntLLROutputS1xD(303)(4);
  CNStageIntLLRInputS2xD(293)(4) <= VNStageIntLLROutputS1xD(303)(5);
  CNStageIntLLRInputS2xD(382)(4) <= VNStageIntLLROutputS1xD(303)(6);
  CNStageIntLLRInputS2xD(7)(4) <= VNStageIntLLROutputS1xD(304)(0);
  CNStageIntLLRInputS2xD(97)(4) <= VNStageIntLLROutputS1xD(304)(1);
  CNStageIntLLRInputS2xD(157)(4) <= VNStageIntLLROutputS1xD(304)(2);
  CNStageIntLLRInputS2xD(222)(4) <= VNStageIntLLROutputS1xD(304)(3);
  CNStageIntLLRInputS2xD(263)(4) <= VNStageIntLLROutputS1xD(304)(4);
  CNStageIntLLRInputS2xD(283)(4) <= VNStageIntLLROutputS1xD(304)(5);
  CNStageIntLLRInputS2xD(359)(4) <= VNStageIntLLROutputS1xD(304)(6);
  CNStageIntLLRInputS2xD(6)(4) <= VNStageIntLLROutputS1xD(305)(0);
  CNStageIntLLRInputS2xD(80)(4) <= VNStageIntLLROutputS1xD(305)(1);
  CNStageIntLLRInputS2xD(115)(4) <= VNStageIntLLROutputS1xD(305)(2);
  CNStageIntLLRInputS2xD(209)(4) <= VNStageIntLLROutputS1xD(305)(3);
  CNStageIntLLRInputS2xD(276)(4) <= VNStageIntLLROutputS1xD(305)(4);
  CNStageIntLLRInputS2xD(323)(4) <= VNStageIntLLROutputS1xD(305)(5);
  CNStageIntLLRInputS2xD(342)(4) <= VNStageIntLLROutputS1xD(305)(6);
  CNStageIntLLRInputS2xD(5)(4) <= VNStageIntLLROutputS1xD(306)(0);
  CNStageIntLLRInputS2xD(87)(4) <= VNStageIntLLROutputS1xD(306)(1);
  CNStageIntLLRInputS2xD(136)(4) <= VNStageIntLLROutputS1xD(306)(2);
  CNStageIntLLRInputS2xD(174)(4) <= VNStageIntLLROutputS1xD(306)(3);
  CNStageIntLLRInputS2xD(4)(4) <= VNStageIntLLROutputS1xD(307)(0);
  CNStageIntLLRInputS2xD(107)(4) <= VNStageIntLLROutputS1xD(307)(1);
  CNStageIntLLRInputS2xD(145)(4) <= VNStageIntLLROutputS1xD(307)(2);
  CNStageIntLLRInputS2xD(202)(4) <= VNStageIntLLROutputS1xD(307)(3);
  CNStageIntLLRInputS2xD(230)(4) <= VNStageIntLLROutputS1xD(307)(4);
  CNStageIntLLRInputS2xD(302)(4) <= VNStageIntLLROutputS1xD(307)(5);
  CNStageIntLLRInputS2xD(366)(4) <= VNStageIntLLROutputS1xD(307)(6);
  CNStageIntLLRInputS2xD(140)(4) <= VNStageIntLLROutputS1xD(308)(0);
  CNStageIntLLRInputS2xD(199)(4) <= VNStageIntLLROutputS1xD(308)(1);
  CNStageIntLLRInputS2xD(251)(4) <= VNStageIntLLROutputS1xD(308)(2);
  CNStageIntLLRInputS2xD(311)(4) <= VNStageIntLLROutputS1xD(308)(3);
  CNStageIntLLRInputS2xD(336)(4) <= VNStageIntLLROutputS1xD(308)(4);
  CNStageIntLLRInputS2xD(3)(4) <= VNStageIntLLROutputS1xD(309)(0);
  CNStageIntLLRInputS2xD(86)(4) <= VNStageIntLLROutputS1xD(309)(1);
  CNStageIntLLRInputS2xD(146)(4) <= VNStageIntLLROutputS1xD(309)(2);
  CNStageIntLLRInputS2xD(214)(4) <= VNStageIntLLROutputS1xD(309)(3);
  CNStageIntLLRInputS2xD(265)(4) <= VNStageIntLLROutputS1xD(309)(4);
  CNStageIntLLRInputS2xD(307)(4) <= VNStageIntLLROutputS1xD(309)(5);
  CNStageIntLLRInputS2xD(2)(4) <= VNStageIntLLROutputS1xD(310)(0);
  CNStageIntLLRInputS2xD(65)(4) <= VNStageIntLLROutputS1xD(310)(1);
  CNStageIntLLRInputS2xD(135)(4) <= VNStageIntLLROutputS1xD(310)(2);
  CNStageIntLLRInputS2xD(261)(4) <= VNStageIntLLROutputS1xD(310)(3);
  CNStageIntLLRInputS2xD(312)(4) <= VNStageIntLLROutputS1xD(310)(4);
  CNStageIntLLRInputS2xD(369)(4) <= VNStageIntLLROutputS1xD(310)(5);
  CNStageIntLLRInputS2xD(1)(4) <= VNStageIntLLROutputS1xD(311)(0);
  CNStageIntLLRInputS2xD(68)(4) <= VNStageIntLLROutputS1xD(311)(1);
  CNStageIntLLRInputS2xD(160)(4) <= VNStageIntLLROutputS1xD(311)(2);
  CNStageIntLLRInputS2xD(225)(4) <= VNStageIntLLROutputS1xD(311)(3);
  CNStageIntLLRInputS2xD(301)(4) <= VNStageIntLLROutputS1xD(311)(4);
  CNStageIntLLRInputS2xD(0)(4) <= VNStageIntLLROutputS1xD(312)(0);
  CNStageIntLLRInputS2xD(108)(4) <= VNStageIntLLROutputS1xD(312)(1);
  CNStageIntLLRInputS2xD(167)(4) <= VNStageIntLLROutputS1xD(312)(2);
  CNStageIntLLRInputS2xD(246)(4) <= VNStageIntLLROutputS1xD(312)(3);
  CNStageIntLLRInputS2xD(326)(4) <= VNStageIntLLROutputS1xD(312)(4);
  CNStageIntLLRInputS2xD(348)(4) <= VNStageIntLLROutputS1xD(312)(5);
  CNStageIntLLRInputS2xD(150)(4) <= VNStageIntLLROutputS1xD(313)(0);
  CNStageIntLLRInputS2xD(188)(4) <= VNStageIntLLROutputS1xD(313)(1);
  CNStageIntLLRInputS2xD(247)(4) <= VNStageIntLLROutputS1xD(313)(2);
  CNStageIntLLRInputS2xD(356)(4) <= VNStageIntLLROutputS1xD(313)(3);
  CNStageIntLLRInputS2xD(191)(4) <= VNStageIntLLROutputS1xD(314)(0);
  CNStageIntLLRInputS2xD(278)(4) <= VNStageIntLLROutputS1xD(314)(1);
  CNStageIntLLRInputS2xD(316)(4) <= VNStageIntLLROutputS1xD(314)(2);
  CNStageIntLLRInputS2xD(352)(4) <= VNStageIntLLROutputS1xD(314)(3);
  CNStageIntLLRInputS2xD(78)(4) <= VNStageIntLLROutputS1xD(315)(0);
  CNStageIntLLRInputS2xD(119)(4) <= VNStageIntLLROutputS1xD(315)(1);
  CNStageIntLLRInputS2xD(183)(4) <= VNStageIntLLROutputS1xD(315)(2);
  CNStageIntLLRInputS2xD(271)(4) <= VNStageIntLLROutputS1xD(315)(3);
  CNStageIntLLRInputS2xD(318)(4) <= VNStageIntLLROutputS1xD(315)(4);
  CNStageIntLLRInputS2xD(357)(4) <= VNStageIntLLROutputS1xD(315)(5);
  CNStageIntLLRInputS2xD(61)(4) <= VNStageIntLLROutputS1xD(316)(0);
  CNStageIntLLRInputS2xD(158)(4) <= VNStageIntLLROutputS1xD(316)(1);
  CNStageIntLLRInputS2xD(234)(4) <= VNStageIntLLROutputS1xD(316)(2);
  CNStageIntLLRInputS2xD(288)(4) <= VNStageIntLLROutputS1xD(316)(3);
  CNStageIntLLRInputS2xD(347)(4) <= VNStageIntLLROutputS1xD(316)(4);
  CNStageIntLLRInputS2xD(88)(4) <= VNStageIntLLROutputS1xD(317)(0);
  CNStageIntLLRInputS2xD(238)(4) <= VNStageIntLLROutputS1xD(317)(1);
  CNStageIntLLRInputS2xD(324)(4) <= VNStageIntLLROutputS1xD(317)(2);
  CNStageIntLLRInputS2xD(372)(4) <= VNStageIntLLROutputS1xD(317)(3);
  CNStageIntLLRInputS2xD(120)(4) <= VNStageIntLLROutputS1xD(318)(0);
  CNStageIntLLRInputS2xD(210)(4) <= VNStageIntLLROutputS1xD(318)(1);
  CNStageIntLLRInputS2xD(279)(4) <= VNStageIntLLROutputS1xD(318)(2);
  CNStageIntLLRInputS2xD(379)(4) <= VNStageIntLLROutputS1xD(318)(3);
  CNStageIntLLRInputS2xD(52)(4) <= VNStageIntLLROutputS1xD(319)(0);
  CNStageIntLLRInputS2xD(66)(4) <= VNStageIntLLROutputS1xD(319)(1);
  CNStageIntLLRInputS2xD(151)(4) <= VNStageIntLLROutputS1xD(319)(2);
  CNStageIntLLRInputS2xD(221)(4) <= VNStageIntLLROutputS1xD(319)(3);
  CNStageIntLLRInputS2xD(237)(4) <= VNStageIntLLROutputS1xD(319)(4);
  CNStageIntLLRInputS2xD(289)(4) <= VNStageIntLLROutputS1xD(319)(5);
  CNStageIntLLRInputS2xD(361)(4) <= VNStageIntLLROutputS1xD(319)(6);
  CNStageIntLLRInputS2xD(53)(5) <= VNStageIntLLROutputS1xD(320)(0);
  CNStageIntLLRInputS2xD(126)(5) <= VNStageIntLLROutputS1xD(320)(1);
  CNStageIntLLRInputS2xD(196)(5) <= VNStageIntLLROutputS1xD(320)(2);
  CNStageIntLLRInputS2xD(295)(5) <= VNStageIntLLROutputS1xD(320)(3);
  CNStageIntLLRInputS2xD(338)(5) <= VNStageIntLLROutputS1xD(320)(4);
  CNStageIntLLRInputS2xD(51)(5) <= VNStageIntLLROutputS1xD(321)(0);
  CNStageIntLLRInputS2xD(65)(5) <= VNStageIntLLROutputS1xD(321)(1);
  CNStageIntLLRInputS2xD(150)(5) <= VNStageIntLLROutputS1xD(321)(2);
  CNStageIntLLRInputS2xD(220)(5) <= VNStageIntLLROutputS1xD(321)(3);
  CNStageIntLLRInputS2xD(236)(5) <= VNStageIntLLROutputS1xD(321)(4);
  CNStageIntLLRInputS2xD(288)(5) <= VNStageIntLLROutputS1xD(321)(5);
  CNStageIntLLRInputS2xD(360)(5) <= VNStageIntLLROutputS1xD(321)(6);
  CNStageIntLLRInputS2xD(50)(5) <= VNStageIntLLROutputS1xD(322)(0);
  CNStageIntLLRInputS2xD(84)(5) <= VNStageIntLLROutputS1xD(322)(1);
  CNStageIntLLRInputS2xD(165)(5) <= VNStageIntLLROutputS1xD(322)(2);
  CNStageIntLLRInputS2xD(231)(5) <= VNStageIntLLROutputS1xD(322)(3);
  CNStageIntLLRInputS2xD(316)(5) <= VNStageIntLLROutputS1xD(322)(4);
  CNStageIntLLRInputS2xD(362)(5) <= VNStageIntLLROutputS1xD(322)(5);
  CNStageIntLLRInputS2xD(56)(5) <= VNStageIntLLROutputS1xD(323)(0);
  CNStageIntLLRInputS2xD(136)(5) <= VNStageIntLLROutputS1xD(323)(1);
  CNStageIntLLRInputS2xD(184)(5) <= VNStageIntLLROutputS1xD(323)(2);
  CNStageIntLLRInputS2xD(268)(5) <= VNStageIntLLROutputS1xD(323)(3);
  CNStageIntLLRInputS2xD(330)(5) <= VNStageIntLLROutputS1xD(323)(4);
  CNStageIntLLRInputS2xD(49)(5) <= VNStageIntLLROutputS1xD(324)(0);
  CNStageIntLLRInputS2xD(109)(5) <= VNStageIntLLROutputS1xD(324)(1);
  CNStageIntLLRInputS2xD(113)(5) <= VNStageIntLLROutputS1xD(324)(2);
  CNStageIntLLRInputS2xD(223)(5) <= VNStageIntLLROutputS1xD(324)(3);
  CNStageIntLLRInputS2xD(273)(5) <= VNStageIntLLROutputS1xD(324)(4);
  CNStageIntLLRInputS2xD(302)(5) <= VNStageIntLLROutputS1xD(324)(5);
  CNStageIntLLRInputS2xD(369)(5) <= VNStageIntLLROutputS1xD(324)(6);
  CNStageIntLLRInputS2xD(48)(5) <= VNStageIntLLROutputS1xD(325)(0);
  CNStageIntLLRInputS2xD(70)(5) <= VNStageIntLLROutputS1xD(325)(1);
  CNStageIntLLRInputS2xD(137)(5) <= VNStageIntLLROutputS1xD(325)(2);
  CNStageIntLLRInputS2xD(185)(5) <= VNStageIntLLROutputS1xD(325)(3);
  CNStageIntLLRInputS2xD(242)(5) <= VNStageIntLLROutputS1xD(325)(4);
  CNStageIntLLRInputS2xD(284)(5) <= VNStageIntLLROutputS1xD(325)(5);
  CNStageIntLLRInputS2xD(382)(5) <= VNStageIntLLROutputS1xD(325)(6);
  CNStageIntLLRInputS2xD(47)(5) <= VNStageIntLLROutputS1xD(326)(0);
  CNStageIntLLRInputS2xD(62)(5) <= VNStageIntLLROutputS1xD(326)(1);
  CNStageIntLLRInputS2xD(203)(5) <= VNStageIntLLROutputS1xD(326)(2);
  CNStageIntLLRInputS2xD(241)(5) <= VNStageIntLLROutputS1xD(326)(3);
  CNStageIntLLRInputS2xD(304)(5) <= VNStageIntLLROutputS1xD(326)(4);
  CNStageIntLLRInputS2xD(46)(5) <= VNStageIntLLROutputS1xD(327)(0);
  CNStageIntLLRInputS2xD(94)(5) <= VNStageIntLLROutputS1xD(327)(1);
  CNStageIntLLRInputS2xD(148)(5) <= VNStageIntLLROutputS1xD(327)(2);
  CNStageIntLLRInputS2xD(211)(5) <= VNStageIntLLROutputS1xD(327)(3);
  CNStageIntLLRInputS2xD(272)(5) <= VNStageIntLLROutputS1xD(327)(4);
  CNStageIntLLRInputS2xD(318)(5) <= VNStageIntLLROutputS1xD(327)(5);
  CNStageIntLLRInputS2xD(361)(5) <= VNStageIntLLROutputS1xD(327)(6);
  CNStageIntLLRInputS2xD(45)(5) <= VNStageIntLLROutputS1xD(328)(0);
  CNStageIntLLRInputS2xD(103)(5) <= VNStageIntLLROutputS1xD(328)(1);
  CNStageIntLLRInputS2xD(168)(5) <= VNStageIntLLROutputS1xD(328)(2);
  CNStageIntLLRInputS2xD(314)(5) <= VNStageIntLLROutputS1xD(328)(3);
  CNStageIntLLRInputS2xD(377)(5) <= VNStageIntLLROutputS1xD(328)(4);
  CNStageIntLLRInputS2xD(44)(5) <= VNStageIntLLROutputS1xD(329)(0);
  CNStageIntLLRInputS2xD(97)(5) <= VNStageIntLLROutputS1xD(329)(1);
  CNStageIntLLRInputS2xD(131)(5) <= VNStageIntLLROutputS1xD(329)(2);
  CNStageIntLLRInputS2xD(212)(5) <= VNStageIntLLROutputS1xD(329)(3);
  CNStageIntLLRInputS2xD(255)(5) <= VNStageIntLLROutputS1xD(329)(4);
  CNStageIntLLRInputS2xD(280)(5) <= VNStageIntLLROutputS1xD(329)(5);
  CNStageIntLLRInputS2xD(348)(5) <= VNStageIntLLROutputS1xD(329)(6);
  CNStageIntLLRInputS2xD(43)(5) <= VNStageIntLLROutputS1xD(330)(0);
  CNStageIntLLRInputS2xD(101)(5) <= VNStageIntLLROutputS1xD(330)(1);
  CNStageIntLLRInputS2xD(132)(5) <= VNStageIntLLROutputS1xD(330)(2);
  CNStageIntLLRInputS2xD(202)(5) <= VNStageIntLLROutputS1xD(330)(3);
  CNStageIntLLRInputS2xD(243)(5) <= VNStageIntLLROutputS1xD(330)(4);
  CNStageIntLLRInputS2xD(42)(5) <= VNStageIntLLROutputS1xD(331)(0);
  CNStageIntLLRInputS2xD(92)(5) <= VNStageIntLLROutputS1xD(331)(1);
  CNStageIntLLRInputS2xD(167)(5) <= VNStageIntLLROutputS1xD(331)(2);
  CNStageIntLLRInputS2xD(172)(5) <= VNStageIntLLROutputS1xD(331)(3);
  CNStageIntLLRInputS2xD(350)(5) <= VNStageIntLLROutputS1xD(331)(4);
  CNStageIntLLRInputS2xD(41)(5) <= VNStageIntLLROutputS1xD(332)(0);
  CNStageIntLLRInputS2xD(71)(5) <= VNStageIntLLROutputS1xD(332)(1);
  CNStageIntLLRInputS2xD(158)(5) <= VNStageIntLLROutputS1xD(332)(2);
  CNStageIntLLRInputS2xD(179)(5) <= VNStageIntLLROutputS1xD(332)(3);
  CNStageIntLLRInputS2xD(240)(5) <= VNStageIntLLROutputS1xD(332)(4);
  CNStageIntLLRInputS2xD(363)(5) <= VNStageIntLLROutputS1xD(332)(5);
  CNStageIntLLRInputS2xD(108)(5) <= VNStageIntLLROutputS1xD(333)(0);
  CNStageIntLLRInputS2xD(117)(5) <= VNStageIntLLROutputS1xD(333)(1);
  CNStageIntLLRInputS2xD(215)(5) <= VNStageIntLLROutputS1xD(333)(2);
  CNStageIntLLRInputS2xD(265)(5) <= VNStageIntLLROutputS1xD(333)(3);
  CNStageIntLLRInputS2xD(324)(5) <= VNStageIntLLROutputS1xD(333)(4);
  CNStageIntLLRInputS2xD(359)(5) <= VNStageIntLLROutputS1xD(333)(5);
  CNStageIntLLRInputS2xD(40)(5) <= VNStageIntLLROutputS1xD(334)(0);
  CNStageIntLLRInputS2xD(66)(5) <= VNStageIntLLROutputS1xD(334)(1);
  CNStageIntLLRInputS2xD(217)(5) <= VNStageIntLLROutputS1xD(334)(2);
  CNStageIntLLRInputS2xD(286)(5) <= VNStageIntLLROutputS1xD(334)(3);
  CNStageIntLLRInputS2xD(380)(5) <= VNStageIntLLROutputS1xD(334)(4);
  CNStageIntLLRInputS2xD(39)(5) <= VNStageIntLLROutputS1xD(335)(0);
  CNStageIntLLRInputS2xD(78)(5) <= VNStageIntLLROutputS1xD(335)(1);
  CNStageIntLLRInputS2xD(170)(5) <= VNStageIntLLROutputS1xD(335)(2);
  CNStageIntLLRInputS2xD(189)(5) <= VNStageIntLLROutputS1xD(335)(3);
  CNStageIntLLRInputS2xD(274)(5) <= VNStageIntLLROutputS1xD(335)(4);
  CNStageIntLLRInputS2xD(291)(5) <= VNStageIntLLROutputS1xD(335)(5);
  CNStageIntLLRInputS2xD(343)(5) <= VNStageIntLLROutputS1xD(335)(6);
  CNStageIntLLRInputS2xD(38)(5) <= VNStageIntLLROutputS1xD(336)(0);
  CNStageIntLLRInputS2xD(104)(5) <= VNStageIntLLROutputS1xD(336)(1);
  CNStageIntLLRInputS2xD(121)(5) <= VNStageIntLLROutputS1xD(336)(2);
  CNStageIntLLRInputS2xD(267)(5) <= VNStageIntLLROutputS1xD(336)(3);
  CNStageIntLLRInputS2xD(332)(5) <= VNStageIntLLROutputS1xD(336)(4);
  CNStageIntLLRInputS2xD(344)(5) <= VNStageIntLLROutputS1xD(336)(5);
  CNStageIntLLRInputS2xD(37)(5) <= VNStageIntLLROutputS1xD(337)(0);
  CNStageIntLLRInputS2xD(93)(5) <= VNStageIntLLROutputS1xD(337)(1);
  CNStageIntLLRInputS2xD(115)(5) <= VNStageIntLLROutputS1xD(337)(2);
  CNStageIntLLRInputS2xD(183)(5) <= VNStageIntLLROutputS1xD(337)(3);
  CNStageIntLLRInputS2xD(253)(5) <= VNStageIntLLROutputS1xD(337)(4);
  CNStageIntLLRInputS2xD(290)(5) <= VNStageIntLLROutputS1xD(337)(5);
  CNStageIntLLRInputS2xD(379)(5) <= VNStageIntLLROutputS1xD(337)(6);
  CNStageIntLLRInputS2xD(36)(5) <= VNStageIntLLROutputS1xD(338)(0);
  CNStageIntLLRInputS2xD(80)(5) <= VNStageIntLLROutputS1xD(338)(1);
  CNStageIntLLRInputS2xD(155)(5) <= VNStageIntLLROutputS1xD(338)(2);
  CNStageIntLLRInputS2xD(190)(5) <= VNStageIntLLROutputS1xD(338)(3);
  CNStageIntLLRInputS2xD(370)(5) <= VNStageIntLLROutputS1xD(338)(4);
  CNStageIntLLRInputS2xD(35)(5) <= VNStageIntLLROutputS1xD(339)(0);
  CNStageIntLLRInputS2xD(96)(5) <= VNStageIntLLROutputS1xD(339)(1);
  CNStageIntLLRInputS2xD(163)(5) <= VNStageIntLLROutputS1xD(339)(2);
  CNStageIntLLRInputS2xD(216)(5) <= VNStageIntLLROutputS1xD(339)(3);
  CNStageIntLLRInputS2xD(247)(5) <= VNStageIntLLROutputS1xD(339)(4);
  CNStageIntLLRInputS2xD(322)(5) <= VNStageIntLLROutputS1xD(339)(5);
  CNStageIntLLRInputS2xD(34)(5) <= VNStageIntLLROutputS1xD(340)(0);
  CNStageIntLLRInputS2xD(58)(5) <= VNStageIntLLROutputS1xD(340)(1);
  CNStageIntLLRInputS2xD(127)(5) <= VNStageIntLLROutputS1xD(340)(2);
  CNStageIntLLRInputS2xD(178)(5) <= VNStageIntLLROutputS1xD(340)(3);
  CNStageIntLLRInputS2xD(245)(5) <= VNStageIntLLROutputS1xD(340)(4);
  CNStageIntLLRInputS2xD(334)(5) <= VNStageIntLLROutputS1xD(340)(5);
  CNStageIntLLRInputS2xD(33)(5) <= VNStageIntLLROutputS1xD(341)(0);
  CNStageIntLLRInputS2xD(68)(5) <= VNStageIntLLROutputS1xD(341)(1);
  CNStageIntLLRInputS2xD(125)(5) <= VNStageIntLLROutputS1xD(341)(2);
  CNStageIntLLRInputS2xD(204)(5) <= VNStageIntLLROutputS1xD(341)(3);
  CNStageIntLLRInputS2xD(258)(5) <= VNStageIntLLROutputS1xD(341)(4);
  CNStageIntLLRInputS2xD(296)(5) <= VNStageIntLLROutputS1xD(341)(5);
  CNStageIntLLRInputS2xD(32)(5) <= VNStageIntLLROutputS1xD(342)(0);
  CNStageIntLLRInputS2xD(63)(5) <= VNStageIntLLROutputS1xD(342)(1);
  CNStageIntLLRInputS2xD(161)(5) <= VNStageIntLLROutputS1xD(342)(2);
  CNStageIntLLRInputS2xD(251)(5) <= VNStageIntLLROutputS1xD(342)(3);
  CNStageIntLLRInputS2xD(294)(5) <= VNStageIntLLROutputS1xD(342)(4);
  CNStageIntLLRInputS2xD(31)(5) <= VNStageIntLLROutputS1xD(343)(0);
  CNStageIntLLRInputS2xD(69)(5) <= VNStageIntLLROutputS1xD(343)(1);
  CNStageIntLLRInputS2xD(140)(5) <= VNStageIntLLROutputS1xD(343)(2);
  CNStageIntLLRInputS2xD(206)(5) <= VNStageIntLLROutputS1xD(343)(3);
  CNStageIntLLRInputS2xD(228)(5) <= VNStageIntLLROutputS1xD(343)(4);
  CNStageIntLLRInputS2xD(327)(5) <= VNStageIntLLROutputS1xD(343)(5);
  CNStageIntLLRInputS2xD(30)(5) <= VNStageIntLLROutputS1xD(344)(0);
  CNStageIntLLRInputS2xD(57)(5) <= VNStageIntLLROutputS1xD(344)(1);
  CNStageIntLLRInputS2xD(143)(5) <= VNStageIntLLROutputS1xD(344)(2);
  CNStageIntLLRInputS2xD(218)(5) <= VNStageIntLLROutputS1xD(344)(3);
  CNStageIntLLRInputS2xD(238)(5) <= VNStageIntLLROutputS1xD(344)(4);
  CNStageIntLLRInputS2xD(307)(5) <= VNStageIntLLROutputS1xD(344)(5);
  CNStageIntLLRInputS2xD(367)(5) <= VNStageIntLLROutputS1xD(344)(6);
  CNStageIntLLRInputS2xD(29)(5) <= VNStageIntLLROutputS1xD(345)(0);
  CNStageIntLLRInputS2xD(83)(5) <= VNStageIntLLROutputS1xD(345)(1);
  CNStageIntLLRInputS2xD(128)(5) <= VNStageIntLLROutputS1xD(345)(2);
  CNStageIntLLRInputS2xD(232)(5) <= VNStageIntLLROutputS1xD(345)(3);
  CNStageIntLLRInputS2xD(309)(5) <= VNStageIntLLROutputS1xD(345)(4);
  CNStageIntLLRInputS2xD(375)(5) <= VNStageIntLLROutputS1xD(345)(5);
  CNStageIntLLRInputS2xD(28)(5) <= VNStageIntLLROutputS1xD(346)(0);
  CNStageIntLLRInputS2xD(89)(5) <= VNStageIntLLROutputS1xD(346)(1);
  CNStageIntLLRInputS2xD(162)(5) <= VNStageIntLLROutputS1xD(346)(2);
  CNStageIntLLRInputS2xD(181)(5) <= VNStageIntLLROutputS1xD(346)(3);
  CNStageIntLLRInputS2xD(235)(5) <= VNStageIntLLROutputS1xD(346)(4);
  CNStageIntLLRInputS2xD(297)(5) <= VNStageIntLLROutputS1xD(346)(5);
  CNStageIntLLRInputS2xD(339)(5) <= VNStageIntLLROutputS1xD(346)(6);
  CNStageIntLLRInputS2xD(27)(5) <= VNStageIntLLROutputS1xD(347)(0);
  CNStageIntLLRInputS2xD(73)(5) <= VNStageIntLLROutputS1xD(347)(1);
  CNStageIntLLRInputS2xD(124)(5) <= VNStageIntLLROutputS1xD(347)(2);
  CNStageIntLLRInputS2xD(199)(5) <= VNStageIntLLROutputS1xD(347)(3);
  CNStageIntLLRInputS2xD(225)(5) <= VNStageIntLLROutputS1xD(347)(4);
  CNStageIntLLRInputS2xD(328)(5) <= VNStageIntLLROutputS1xD(347)(5);
  CNStageIntLLRInputS2xD(337)(5) <= VNStageIntLLROutputS1xD(347)(6);
  CNStageIntLLRInputS2xD(26)(5) <= VNStageIntLLROutputS1xD(348)(0);
  CNStageIntLLRInputS2xD(75)(5) <= VNStageIntLLROutputS1xD(348)(1);
  CNStageIntLLRInputS2xD(152)(5) <= VNStageIntLLROutputS1xD(348)(2);
  CNStageIntLLRInputS2xD(200)(5) <= VNStageIntLLROutputS1xD(348)(3);
  CNStageIntLLRInputS2xD(259)(5) <= VNStageIntLLROutputS1xD(348)(4);
  CNStageIntLLRInputS2xD(293)(5) <= VNStageIntLLROutputS1xD(348)(5);
  CNStageIntLLRInputS2xD(373)(5) <= VNStageIntLLROutputS1xD(348)(6);
  CNStageIntLLRInputS2xD(25)(5) <= VNStageIntLLROutputS1xD(349)(0);
  CNStageIntLLRInputS2xD(99)(5) <= VNStageIntLLROutputS1xD(349)(1);
  CNStageIntLLRInputS2xD(180)(5) <= VNStageIntLLROutputS1xD(349)(2);
  CNStageIntLLRInputS2xD(244)(5) <= VNStageIntLLROutputS1xD(349)(3);
  CNStageIntLLRInputS2xD(319)(5) <= VNStageIntLLROutputS1xD(349)(4);
  CNStageIntLLRInputS2xD(352)(5) <= VNStageIntLLROutputS1xD(349)(5);
  CNStageIntLLRInputS2xD(24)(5) <= VNStageIntLLROutputS1xD(350)(0);
  CNStageIntLLRInputS2xD(81)(5) <= VNStageIntLLROutputS1xD(350)(1);
  CNStageIntLLRInputS2xD(164)(5) <= VNStageIntLLROutputS1xD(350)(2);
  CNStageIntLLRInputS2xD(171)(5) <= VNStageIntLLROutputS1xD(350)(3);
  CNStageIntLLRInputS2xD(254)(5) <= VNStageIntLLROutputS1xD(350)(4);
  CNStageIntLLRInputS2xD(303)(5) <= VNStageIntLLROutputS1xD(350)(5);
  CNStageIntLLRInputS2xD(23)(5) <= VNStageIntLLROutputS1xD(351)(0);
  CNStageIntLLRInputS2xD(154)(5) <= VNStageIntLLROutputS1xD(351)(1);
  CNStageIntLLRInputS2xD(188)(5) <= VNStageIntLLROutputS1xD(351)(2);
  CNStageIntLLRInputS2xD(266)(5) <= VNStageIntLLROutputS1xD(351)(3);
  CNStageIntLLRInputS2xD(329)(5) <= VNStageIntLLROutputS1xD(351)(4);
  CNStageIntLLRInputS2xD(340)(5) <= VNStageIntLLROutputS1xD(351)(5);
  CNStageIntLLRInputS2xD(22)(5) <= VNStageIntLLROutputS1xD(352)(0);
  CNStageIntLLRInputS2xD(100)(5) <= VNStageIntLLROutputS1xD(352)(1);
  CNStageIntLLRInputS2xD(141)(5) <= VNStageIntLLROutputS1xD(352)(2);
  CNStageIntLLRInputS2xD(192)(5) <= VNStageIntLLROutputS1xD(352)(3);
  CNStageIntLLRInputS2xD(239)(5) <= VNStageIntLLROutputS1xD(352)(4);
  CNStageIntLLRInputS2xD(321)(5) <= VNStageIntLLROutputS1xD(352)(5);
  CNStageIntLLRInputS2xD(374)(5) <= VNStageIntLLROutputS1xD(352)(6);
  CNStageIntLLRInputS2xD(21)(5) <= VNStageIntLLROutputS1xD(353)(0);
  CNStageIntLLRInputS2xD(74)(5) <= VNStageIntLLROutputS1xD(353)(1);
  CNStageIntLLRInputS2xD(160)(5) <= VNStageIntLLROutputS1xD(353)(2);
  CNStageIntLLRInputS2xD(224)(5) <= VNStageIntLLROutputS1xD(353)(3);
  CNStageIntLLRInputS2xD(227)(5) <= VNStageIntLLROutputS1xD(353)(4);
  CNStageIntLLRInputS2xD(336)(5) <= VNStageIntLLROutputS1xD(353)(5);
  CNStageIntLLRInputS2xD(20)(5) <= VNStageIntLLROutputS1xD(354)(0);
  CNStageIntLLRInputS2xD(88)(5) <= VNStageIntLLROutputS1xD(354)(1);
  CNStageIntLLRInputS2xD(133)(5) <= VNStageIntLLROutputS1xD(354)(2);
  CNStageIntLLRInputS2xD(191)(5) <= VNStageIntLLROutputS1xD(354)(3);
  CNStageIntLLRInputS2xD(326)(5) <= VNStageIntLLROutputS1xD(354)(4);
  CNStageIntLLRInputS2xD(364)(5) <= VNStageIntLLROutputS1xD(354)(5);
  CNStageIntLLRInputS2xD(19)(5) <= VNStageIntLLROutputS1xD(355)(0);
  CNStageIntLLRInputS2xD(59)(5) <= VNStageIntLLROutputS1xD(355)(1);
  CNStageIntLLRInputS2xD(130)(5) <= VNStageIntLLROutputS1xD(355)(2);
  CNStageIntLLRInputS2xD(186)(5) <= VNStageIntLLROutputS1xD(355)(3);
  CNStageIntLLRInputS2xD(230)(5) <= VNStageIntLLROutputS1xD(355)(4);
  CNStageIntLLRInputS2xD(300)(5) <= VNStageIntLLROutputS1xD(355)(5);
  CNStageIntLLRInputS2xD(349)(5) <= VNStageIntLLROutputS1xD(355)(6);
  CNStageIntLLRInputS2xD(18)(5) <= VNStageIntLLROutputS1xD(356)(0);
  CNStageIntLLRInputS2xD(95)(5) <= VNStageIntLLROutputS1xD(356)(1);
  CNStageIntLLRInputS2xD(146)(5) <= VNStageIntLLROutputS1xD(356)(2);
  CNStageIntLLRInputS2xD(222)(5) <= VNStageIntLLROutputS1xD(356)(3);
  CNStageIntLLRInputS2xD(299)(5) <= VNStageIntLLROutputS1xD(356)(4);
  CNStageIntLLRInputS2xD(376)(5) <= VNStageIntLLROutputS1xD(356)(5);
  CNStageIntLLRInputS2xD(17)(5) <= VNStageIntLLROutputS1xD(357)(0);
  CNStageIntLLRInputS2xD(61)(5) <= VNStageIntLLROutputS1xD(357)(1);
  CNStageIntLLRInputS2xD(138)(5) <= VNStageIntLLROutputS1xD(357)(2);
  CNStageIntLLRInputS2xD(176)(5) <= VNStageIntLLROutputS1xD(357)(3);
  CNStageIntLLRInputS2xD(256)(5) <= VNStageIntLLROutputS1xD(357)(4);
  CNStageIntLLRInputS2xD(312)(5) <= VNStageIntLLROutputS1xD(357)(5);
  CNStageIntLLRInputS2xD(366)(5) <= VNStageIntLLROutputS1xD(357)(6);
  CNStageIntLLRInputS2xD(16)(5) <= VNStageIntLLROutputS1xD(358)(0);
  CNStageIntLLRInputS2xD(76)(5) <= VNStageIntLLROutputS1xD(358)(1);
  CNStageIntLLRInputS2xD(112)(5) <= VNStageIntLLROutputS1xD(358)(2);
  CNStageIntLLRInputS2xD(252)(5) <= VNStageIntLLROutputS1xD(358)(3);
  CNStageIntLLRInputS2xD(305)(5) <= VNStageIntLLROutputS1xD(358)(4);
  CNStageIntLLRInputS2xD(353)(5) <= VNStageIntLLROutputS1xD(358)(5);
  CNStageIntLLRInputS2xD(15)(5) <= VNStageIntLLROutputS1xD(359)(0);
  CNStageIntLLRInputS2xD(72)(5) <= VNStageIntLLROutputS1xD(359)(1);
  CNStageIntLLRInputS2xD(122)(5) <= VNStageIntLLROutputS1xD(359)(2);
  CNStageIntLLRInputS2xD(195)(5) <= VNStageIntLLROutputS1xD(359)(3);
  CNStageIntLLRInputS2xD(257)(5) <= VNStageIntLLROutputS1xD(359)(4);
  CNStageIntLLRInputS2xD(283)(5) <= VNStageIntLLROutputS1xD(359)(5);
  CNStageIntLLRInputS2xD(372)(5) <= VNStageIntLLROutputS1xD(359)(6);
  CNStageIntLLRInputS2xD(14)(5) <= VNStageIntLLROutputS1xD(360)(0);
  CNStageIntLLRInputS2xD(91)(5) <= VNStageIntLLROutputS1xD(360)(1);
  CNStageIntLLRInputS2xD(116)(5) <= VNStageIntLLROutputS1xD(360)(2);
  CNStageIntLLRInputS2xD(174)(5) <= VNStageIntLLROutputS1xD(360)(3);
  CNStageIntLLRInputS2xD(248)(5) <= VNStageIntLLROutputS1xD(360)(4);
  CNStageIntLLRInputS2xD(292)(5) <= VNStageIntLLROutputS1xD(360)(5);
  CNStageIntLLRInputS2xD(345)(5) <= VNStageIntLLROutputS1xD(360)(6);
  CNStageIntLLRInputS2xD(13)(5) <= VNStageIntLLROutputS1xD(361)(0);
  CNStageIntLLRInputS2xD(54)(5) <= VNStageIntLLROutputS1xD(361)(1);
  CNStageIntLLRInputS2xD(120)(5) <= VNStageIntLLROutputS1xD(361)(2);
  CNStageIntLLRInputS2xD(207)(5) <= VNStageIntLLROutputS1xD(361)(3);
  CNStageIntLLRInputS2xD(271)(5) <= VNStageIntLLROutputS1xD(361)(4);
  CNStageIntLLRInputS2xD(285)(5) <= VNStageIntLLROutputS1xD(361)(5);
  CNStageIntLLRInputS2xD(342)(5) <= VNStageIntLLROutputS1xD(361)(6);
  CNStageIntLLRInputS2xD(12)(5) <= VNStageIntLLROutputS1xD(362)(0);
  CNStageIntLLRInputS2xD(55)(5) <= VNStageIntLLROutputS1xD(362)(1);
  CNStageIntLLRInputS2xD(169)(5) <= VNStageIntLLROutputS1xD(362)(2);
  CNStageIntLLRInputS2xD(210)(5) <= VNStageIntLLROutputS1xD(362)(3);
  CNStageIntLLRInputS2xD(276)(5) <= VNStageIntLLROutputS1xD(362)(4);
  CNStageIntLLRInputS2xD(289)(5) <= VNStageIntLLROutputS1xD(362)(5);
  CNStageIntLLRInputS2xD(357)(5) <= VNStageIntLLROutputS1xD(362)(6);
  CNStageIntLLRInputS2xD(90)(5) <= VNStageIntLLROutputS1xD(363)(0);
  CNStageIntLLRInputS2xD(147)(5) <= VNStageIntLLROutputS1xD(363)(1);
  CNStageIntLLRInputS2xD(197)(5) <= VNStageIntLLROutputS1xD(363)(2);
  CNStageIntLLRInputS2xD(261)(5) <= VNStageIntLLROutputS1xD(363)(3);
  CNStageIntLLRInputS2xD(281)(5) <= VNStageIntLLROutputS1xD(363)(4);
  CNStageIntLLRInputS2xD(11)(5) <= VNStageIntLLROutputS1xD(364)(0);
  CNStageIntLLRInputS2xD(82)(5) <= VNStageIntLLROutputS1xD(364)(1);
  CNStageIntLLRInputS2xD(129)(5) <= VNStageIntLLROutputS1xD(364)(2);
  CNStageIntLLRInputS2xD(175)(5) <= VNStageIntLLROutputS1xD(364)(3);
  CNStageIntLLRInputS2xD(263)(5) <= VNStageIntLLROutputS1xD(364)(4);
  CNStageIntLLRInputS2xD(313)(5) <= VNStageIntLLROutputS1xD(364)(5);
  CNStageIntLLRInputS2xD(10)(5) <= VNStageIntLLROutputS1xD(365)(0);
  CNStageIntLLRInputS2xD(98)(5) <= VNStageIntLLROutputS1xD(365)(1);
  CNStageIntLLRInputS2xD(142)(5) <= VNStageIntLLROutputS1xD(365)(2);
  CNStageIntLLRInputS2xD(194)(5) <= VNStageIntLLROutputS1xD(365)(3);
  CNStageIntLLRInputS2xD(234)(5) <= VNStageIntLLROutputS1xD(365)(4);
  CNStageIntLLRInputS2xD(298)(5) <= VNStageIntLLROutputS1xD(365)(5);
  CNStageIntLLRInputS2xD(9)(5) <= VNStageIntLLROutputS1xD(366)(0);
  CNStageIntLLRInputS2xD(102)(5) <= VNStageIntLLROutputS1xD(366)(1);
  CNStageIntLLRInputS2xD(153)(5) <= VNStageIntLLROutputS1xD(366)(2);
  CNStageIntLLRInputS2xD(219)(5) <= VNStageIntLLROutputS1xD(366)(3);
  CNStageIntLLRInputS2xD(269)(5) <= VNStageIntLLROutputS1xD(366)(4);
  CNStageIntLLRInputS2xD(308)(5) <= VNStageIntLLROutputS1xD(366)(5);
  CNStageIntLLRInputS2xD(8)(5) <= VNStageIntLLROutputS1xD(367)(0);
  CNStageIntLLRInputS2xD(110)(5) <= VNStageIntLLROutputS1xD(367)(1);
  CNStageIntLLRInputS2xD(123)(5) <= VNStageIntLLROutputS1xD(367)(2);
  CNStageIntLLRInputS2xD(205)(5) <= VNStageIntLLROutputS1xD(367)(3);
  CNStageIntLLRInputS2xD(226)(5) <= VNStageIntLLROutputS1xD(367)(4);
  CNStageIntLLRInputS2xD(320)(5) <= VNStageIntLLROutputS1xD(367)(5);
  CNStageIntLLRInputS2xD(333)(5) <= VNStageIntLLROutputS1xD(367)(6);
  CNStageIntLLRInputS2xD(7)(5) <= VNStageIntLLROutputS1xD(368)(0);
  CNStageIntLLRInputS2xD(177)(5) <= VNStageIntLLROutputS1xD(368)(1);
  CNStageIntLLRInputS2xD(381)(5) <= VNStageIntLLROutputS1xD(368)(2);
  CNStageIntLLRInputS2xD(6)(5) <= VNStageIntLLROutputS1xD(369)(0);
  CNStageIntLLRInputS2xD(156)(5) <= VNStageIntLLROutputS1xD(369)(1);
  CNStageIntLLRInputS2xD(221)(5) <= VNStageIntLLROutputS1xD(369)(2);
  CNStageIntLLRInputS2xD(262)(5) <= VNStageIntLLROutputS1xD(369)(3);
  CNStageIntLLRInputS2xD(358)(5) <= VNStageIntLLROutputS1xD(369)(4);
  CNStageIntLLRInputS2xD(5)(5) <= VNStageIntLLROutputS1xD(370)(0);
  CNStageIntLLRInputS2xD(114)(5) <= VNStageIntLLROutputS1xD(370)(1);
  CNStageIntLLRInputS2xD(208)(5) <= VNStageIntLLROutputS1xD(370)(2);
  CNStageIntLLRInputS2xD(275)(5) <= VNStageIntLLROutputS1xD(370)(3);
  CNStageIntLLRInputS2xD(341)(5) <= VNStageIntLLROutputS1xD(370)(4);
  CNStageIntLLRInputS2xD(4)(5) <= VNStageIntLLROutputS1xD(371)(0);
  CNStageIntLLRInputS2xD(135)(5) <= VNStageIntLLROutputS1xD(371)(1);
  CNStageIntLLRInputS2xD(173)(5) <= VNStageIntLLROutputS1xD(371)(2);
  CNStageIntLLRInputS2xD(249)(5) <= VNStageIntLLROutputS1xD(371)(3);
  CNStageIntLLRInputS2xD(354)(5) <= VNStageIntLLROutputS1xD(371)(4);
  CNStageIntLLRInputS2xD(106)(5) <= VNStageIntLLROutputS1xD(372)(0);
  CNStageIntLLRInputS2xD(144)(5) <= VNStageIntLLROutputS1xD(372)(1);
  CNStageIntLLRInputS2xD(201)(5) <= VNStageIntLLROutputS1xD(372)(2);
  CNStageIntLLRInputS2xD(229)(5) <= VNStageIntLLROutputS1xD(372)(3);
  CNStageIntLLRInputS2xD(301)(5) <= VNStageIntLLROutputS1xD(372)(4);
  CNStageIntLLRInputS2xD(365)(5) <= VNStageIntLLROutputS1xD(372)(5);
  CNStageIntLLRInputS2xD(3)(5) <= VNStageIntLLROutputS1xD(373)(0);
  CNStageIntLLRInputS2xD(139)(5) <= VNStageIntLLROutputS1xD(373)(1);
  CNStageIntLLRInputS2xD(250)(5) <= VNStageIntLLROutputS1xD(373)(2);
  CNStageIntLLRInputS2xD(310)(5) <= VNStageIntLLROutputS1xD(373)(3);
  CNStageIntLLRInputS2xD(335)(5) <= VNStageIntLLROutputS1xD(373)(4);
  CNStageIntLLRInputS2xD(2)(5) <= VNStageIntLLROutputS1xD(374)(0);
  CNStageIntLLRInputS2xD(85)(5) <= VNStageIntLLROutputS1xD(374)(1);
  CNStageIntLLRInputS2xD(145)(5) <= VNStageIntLLROutputS1xD(374)(2);
  CNStageIntLLRInputS2xD(213)(5) <= VNStageIntLLROutputS1xD(374)(3);
  CNStageIntLLRInputS2xD(264)(5) <= VNStageIntLLROutputS1xD(374)(4);
  CNStageIntLLRInputS2xD(306)(5) <= VNStageIntLLROutputS1xD(374)(5);
  CNStageIntLLRInputS2xD(383)(5) <= VNStageIntLLROutputS1xD(374)(6);
  CNStageIntLLRInputS2xD(1)(5) <= VNStageIntLLROutputS1xD(375)(0);
  CNStageIntLLRInputS2xD(64)(5) <= VNStageIntLLROutputS1xD(375)(1);
  CNStageIntLLRInputS2xD(134)(5) <= VNStageIntLLROutputS1xD(375)(2);
  CNStageIntLLRInputS2xD(260)(5) <= VNStageIntLLROutputS1xD(375)(3);
  CNStageIntLLRInputS2xD(311)(5) <= VNStageIntLLROutputS1xD(375)(4);
  CNStageIntLLRInputS2xD(368)(5) <= VNStageIntLLROutputS1xD(375)(5);
  CNStageIntLLRInputS2xD(0)(5) <= VNStageIntLLROutputS1xD(376)(0);
  CNStageIntLLRInputS2xD(67)(5) <= VNStageIntLLROutputS1xD(376)(1);
  CNStageIntLLRInputS2xD(159)(5) <= VNStageIntLLROutputS1xD(376)(2);
  CNStageIntLLRInputS2xD(278)(5) <= VNStageIntLLROutputS1xD(376)(3);
  CNStageIntLLRInputS2xD(107)(5) <= VNStageIntLLROutputS1xD(377)(0);
  CNStageIntLLRInputS2xD(166)(5) <= VNStageIntLLROutputS1xD(377)(1);
  CNStageIntLLRInputS2xD(193)(5) <= VNStageIntLLROutputS1xD(377)(2);
  CNStageIntLLRInputS2xD(325)(5) <= VNStageIntLLROutputS1xD(377)(3);
  CNStageIntLLRInputS2xD(347)(5) <= VNStageIntLLROutputS1xD(377)(4);
  CNStageIntLLRInputS2xD(86)(5) <= VNStageIntLLROutputS1xD(378)(0);
  CNStageIntLLRInputS2xD(149)(5) <= VNStageIntLLROutputS1xD(378)(1);
  CNStageIntLLRInputS2xD(187)(5) <= VNStageIntLLROutputS1xD(378)(2);
  CNStageIntLLRInputS2xD(246)(5) <= VNStageIntLLROutputS1xD(378)(3);
  CNStageIntLLRInputS2xD(331)(5) <= VNStageIntLLROutputS1xD(378)(4);
  CNStageIntLLRInputS2xD(355)(5) <= VNStageIntLLROutputS1xD(378)(5);
  CNStageIntLLRInputS2xD(105)(5) <= VNStageIntLLROutputS1xD(379)(0);
  CNStageIntLLRInputS2xD(151)(5) <= VNStageIntLLROutputS1xD(379)(1);
  CNStageIntLLRInputS2xD(277)(5) <= VNStageIntLLROutputS1xD(379)(2);
  CNStageIntLLRInputS2xD(315)(5) <= VNStageIntLLROutputS1xD(379)(3);
  CNStageIntLLRInputS2xD(351)(5) <= VNStageIntLLROutputS1xD(379)(4);
  CNStageIntLLRInputS2xD(77)(5) <= VNStageIntLLROutputS1xD(380)(0);
  CNStageIntLLRInputS2xD(118)(5) <= VNStageIntLLROutputS1xD(380)(1);
  CNStageIntLLRInputS2xD(182)(5) <= VNStageIntLLROutputS1xD(380)(2);
  CNStageIntLLRInputS2xD(270)(5) <= VNStageIntLLROutputS1xD(380)(3);
  CNStageIntLLRInputS2xD(317)(5) <= VNStageIntLLROutputS1xD(380)(4);
  CNStageIntLLRInputS2xD(356)(5) <= VNStageIntLLROutputS1xD(380)(5);
  CNStageIntLLRInputS2xD(60)(5) <= VNStageIntLLROutputS1xD(381)(0);
  CNStageIntLLRInputS2xD(157)(5) <= VNStageIntLLROutputS1xD(381)(1);
  CNStageIntLLRInputS2xD(214)(5) <= VNStageIntLLROutputS1xD(381)(2);
  CNStageIntLLRInputS2xD(233)(5) <= VNStageIntLLROutputS1xD(381)(3);
  CNStageIntLLRInputS2xD(287)(5) <= VNStageIntLLROutputS1xD(381)(4);
  CNStageIntLLRInputS2xD(346)(5) <= VNStageIntLLROutputS1xD(381)(5);
  CNStageIntLLRInputS2xD(87)(5) <= VNStageIntLLROutputS1xD(382)(0);
  CNStageIntLLRInputS2xD(111)(5) <= VNStageIntLLROutputS1xD(382)(1);
  CNStageIntLLRInputS2xD(198)(5) <= VNStageIntLLROutputS1xD(382)(2);
  CNStageIntLLRInputS2xD(237)(5) <= VNStageIntLLROutputS1xD(382)(3);
  CNStageIntLLRInputS2xD(323)(5) <= VNStageIntLLROutputS1xD(382)(4);
  CNStageIntLLRInputS2xD(371)(5) <= VNStageIntLLROutputS1xD(382)(5);
  CNStageIntLLRInputS2xD(52)(5) <= VNStageIntLLROutputS1xD(383)(0);
  CNStageIntLLRInputS2xD(79)(5) <= VNStageIntLLROutputS1xD(383)(1);
  CNStageIntLLRInputS2xD(119)(5) <= VNStageIntLLROutputS1xD(383)(2);
  CNStageIntLLRInputS2xD(209)(5) <= VNStageIntLLROutputS1xD(383)(3);
  CNStageIntLLRInputS2xD(279)(5) <= VNStageIntLLROutputS1xD(383)(4);
  CNStageIntLLRInputS2xD(282)(5) <= VNStageIntLLROutputS1xD(383)(5);
  CNStageIntLLRInputS2xD(378)(5) <= VNStageIntLLROutputS1xD(383)(6);

  -- Variable Nodes (Iteration 2)
  VNStageIntLLRInputS2xD(56)(0) <= CNStageIntLLROutputS2xD(0)(0);
  VNStageIntLLRInputS2xD(120)(0) <= CNStageIntLLROutputS2xD(0)(1);
  VNStageIntLLRInputS2xD(184)(0) <= CNStageIntLLROutputS2xD(0)(2);
  VNStageIntLLRInputS2xD(248)(0) <= CNStageIntLLROutputS2xD(0)(3);
  VNStageIntLLRInputS2xD(312)(0) <= CNStageIntLLROutputS2xD(0)(4);
  VNStageIntLLRInputS2xD(376)(0) <= CNStageIntLLROutputS2xD(0)(5);
  VNStageIntLLRInputS2xD(55)(0) <= CNStageIntLLROutputS2xD(1)(0);
  VNStageIntLLRInputS2xD(119)(0) <= CNStageIntLLROutputS2xD(1)(1);
  VNStageIntLLRInputS2xD(183)(0) <= CNStageIntLLROutputS2xD(1)(2);
  VNStageIntLLRInputS2xD(247)(0) <= CNStageIntLLROutputS2xD(1)(3);
  VNStageIntLLRInputS2xD(311)(0) <= CNStageIntLLROutputS2xD(1)(4);
  VNStageIntLLRInputS2xD(375)(0) <= CNStageIntLLROutputS2xD(1)(5);
  VNStageIntLLRInputS2xD(54)(0) <= CNStageIntLLROutputS2xD(2)(0);
  VNStageIntLLRInputS2xD(118)(0) <= CNStageIntLLROutputS2xD(2)(1);
  VNStageIntLLRInputS2xD(182)(0) <= CNStageIntLLROutputS2xD(2)(2);
  VNStageIntLLRInputS2xD(246)(0) <= CNStageIntLLROutputS2xD(2)(3);
  VNStageIntLLRInputS2xD(310)(0) <= CNStageIntLLROutputS2xD(2)(4);
  VNStageIntLLRInputS2xD(374)(0) <= CNStageIntLLROutputS2xD(2)(5);
  VNStageIntLLRInputS2xD(53)(0) <= CNStageIntLLROutputS2xD(3)(0);
  VNStageIntLLRInputS2xD(117)(0) <= CNStageIntLLROutputS2xD(3)(1);
  VNStageIntLLRInputS2xD(181)(0) <= CNStageIntLLROutputS2xD(3)(2);
  VNStageIntLLRInputS2xD(245)(0) <= CNStageIntLLROutputS2xD(3)(3);
  VNStageIntLLRInputS2xD(309)(0) <= CNStageIntLLROutputS2xD(3)(4);
  VNStageIntLLRInputS2xD(373)(0) <= CNStageIntLLROutputS2xD(3)(5);
  VNStageIntLLRInputS2xD(51)(0) <= CNStageIntLLROutputS2xD(4)(0);
  VNStageIntLLRInputS2xD(115)(0) <= CNStageIntLLROutputS2xD(4)(1);
  VNStageIntLLRInputS2xD(179)(0) <= CNStageIntLLROutputS2xD(4)(2);
  VNStageIntLLRInputS2xD(243)(0) <= CNStageIntLLROutputS2xD(4)(3);
  VNStageIntLLRInputS2xD(307)(0) <= CNStageIntLLROutputS2xD(4)(4);
  VNStageIntLLRInputS2xD(371)(0) <= CNStageIntLLROutputS2xD(4)(5);
  VNStageIntLLRInputS2xD(50)(0) <= CNStageIntLLROutputS2xD(5)(0);
  VNStageIntLLRInputS2xD(114)(0) <= CNStageIntLLROutputS2xD(5)(1);
  VNStageIntLLRInputS2xD(178)(0) <= CNStageIntLLROutputS2xD(5)(2);
  VNStageIntLLRInputS2xD(242)(0) <= CNStageIntLLROutputS2xD(5)(3);
  VNStageIntLLRInputS2xD(306)(0) <= CNStageIntLLROutputS2xD(5)(4);
  VNStageIntLLRInputS2xD(370)(0) <= CNStageIntLLROutputS2xD(5)(5);
  VNStageIntLLRInputS2xD(49)(0) <= CNStageIntLLROutputS2xD(6)(0);
  VNStageIntLLRInputS2xD(113)(0) <= CNStageIntLLROutputS2xD(6)(1);
  VNStageIntLLRInputS2xD(177)(0) <= CNStageIntLLROutputS2xD(6)(2);
  VNStageIntLLRInputS2xD(241)(0) <= CNStageIntLLROutputS2xD(6)(3);
  VNStageIntLLRInputS2xD(305)(0) <= CNStageIntLLROutputS2xD(6)(4);
  VNStageIntLLRInputS2xD(369)(0) <= CNStageIntLLROutputS2xD(6)(5);
  VNStageIntLLRInputS2xD(48)(0) <= CNStageIntLLROutputS2xD(7)(0);
  VNStageIntLLRInputS2xD(112)(0) <= CNStageIntLLROutputS2xD(7)(1);
  VNStageIntLLRInputS2xD(176)(0) <= CNStageIntLLROutputS2xD(7)(2);
  VNStageIntLLRInputS2xD(240)(0) <= CNStageIntLLROutputS2xD(7)(3);
  VNStageIntLLRInputS2xD(304)(0) <= CNStageIntLLROutputS2xD(7)(4);
  VNStageIntLLRInputS2xD(368)(0) <= CNStageIntLLROutputS2xD(7)(5);
  VNStageIntLLRInputS2xD(47)(0) <= CNStageIntLLROutputS2xD(8)(0);
  VNStageIntLLRInputS2xD(111)(0) <= CNStageIntLLROutputS2xD(8)(1);
  VNStageIntLLRInputS2xD(175)(0) <= CNStageIntLLROutputS2xD(8)(2);
  VNStageIntLLRInputS2xD(239)(0) <= CNStageIntLLROutputS2xD(8)(3);
  VNStageIntLLRInputS2xD(303)(0) <= CNStageIntLLROutputS2xD(8)(4);
  VNStageIntLLRInputS2xD(367)(0) <= CNStageIntLLROutputS2xD(8)(5);
  VNStageIntLLRInputS2xD(46)(0) <= CNStageIntLLROutputS2xD(9)(0);
  VNStageIntLLRInputS2xD(110)(0) <= CNStageIntLLROutputS2xD(9)(1);
  VNStageIntLLRInputS2xD(174)(0) <= CNStageIntLLROutputS2xD(9)(2);
  VNStageIntLLRInputS2xD(238)(0) <= CNStageIntLLROutputS2xD(9)(3);
  VNStageIntLLRInputS2xD(302)(0) <= CNStageIntLLROutputS2xD(9)(4);
  VNStageIntLLRInputS2xD(366)(0) <= CNStageIntLLROutputS2xD(9)(5);
  VNStageIntLLRInputS2xD(45)(0) <= CNStageIntLLROutputS2xD(10)(0);
  VNStageIntLLRInputS2xD(109)(0) <= CNStageIntLLROutputS2xD(10)(1);
  VNStageIntLLRInputS2xD(173)(0) <= CNStageIntLLROutputS2xD(10)(2);
  VNStageIntLLRInputS2xD(237)(0) <= CNStageIntLLROutputS2xD(10)(3);
  VNStageIntLLRInputS2xD(301)(0) <= CNStageIntLLROutputS2xD(10)(4);
  VNStageIntLLRInputS2xD(365)(0) <= CNStageIntLLROutputS2xD(10)(5);
  VNStageIntLLRInputS2xD(44)(0) <= CNStageIntLLROutputS2xD(11)(0);
  VNStageIntLLRInputS2xD(108)(0) <= CNStageIntLLROutputS2xD(11)(1);
  VNStageIntLLRInputS2xD(172)(0) <= CNStageIntLLROutputS2xD(11)(2);
  VNStageIntLLRInputS2xD(236)(0) <= CNStageIntLLROutputS2xD(11)(3);
  VNStageIntLLRInputS2xD(300)(0) <= CNStageIntLLROutputS2xD(11)(4);
  VNStageIntLLRInputS2xD(364)(0) <= CNStageIntLLROutputS2xD(11)(5);
  VNStageIntLLRInputS2xD(42)(0) <= CNStageIntLLROutputS2xD(12)(0);
  VNStageIntLLRInputS2xD(106)(0) <= CNStageIntLLROutputS2xD(12)(1);
  VNStageIntLLRInputS2xD(170)(0) <= CNStageIntLLROutputS2xD(12)(2);
  VNStageIntLLRInputS2xD(234)(0) <= CNStageIntLLROutputS2xD(12)(3);
  VNStageIntLLRInputS2xD(298)(0) <= CNStageIntLLROutputS2xD(12)(4);
  VNStageIntLLRInputS2xD(362)(0) <= CNStageIntLLROutputS2xD(12)(5);
  VNStageIntLLRInputS2xD(41)(0) <= CNStageIntLLROutputS2xD(13)(0);
  VNStageIntLLRInputS2xD(105)(0) <= CNStageIntLLROutputS2xD(13)(1);
  VNStageIntLLRInputS2xD(169)(0) <= CNStageIntLLROutputS2xD(13)(2);
  VNStageIntLLRInputS2xD(233)(0) <= CNStageIntLLROutputS2xD(13)(3);
  VNStageIntLLRInputS2xD(297)(0) <= CNStageIntLLROutputS2xD(13)(4);
  VNStageIntLLRInputS2xD(361)(0) <= CNStageIntLLROutputS2xD(13)(5);
  VNStageIntLLRInputS2xD(40)(0) <= CNStageIntLLROutputS2xD(14)(0);
  VNStageIntLLRInputS2xD(104)(0) <= CNStageIntLLROutputS2xD(14)(1);
  VNStageIntLLRInputS2xD(168)(0) <= CNStageIntLLROutputS2xD(14)(2);
  VNStageIntLLRInputS2xD(232)(0) <= CNStageIntLLROutputS2xD(14)(3);
  VNStageIntLLRInputS2xD(296)(0) <= CNStageIntLLROutputS2xD(14)(4);
  VNStageIntLLRInputS2xD(360)(0) <= CNStageIntLLROutputS2xD(14)(5);
  VNStageIntLLRInputS2xD(39)(0) <= CNStageIntLLROutputS2xD(15)(0);
  VNStageIntLLRInputS2xD(103)(0) <= CNStageIntLLROutputS2xD(15)(1);
  VNStageIntLLRInputS2xD(167)(0) <= CNStageIntLLROutputS2xD(15)(2);
  VNStageIntLLRInputS2xD(231)(0) <= CNStageIntLLROutputS2xD(15)(3);
  VNStageIntLLRInputS2xD(295)(0) <= CNStageIntLLROutputS2xD(15)(4);
  VNStageIntLLRInputS2xD(359)(0) <= CNStageIntLLROutputS2xD(15)(5);
  VNStageIntLLRInputS2xD(38)(0) <= CNStageIntLLROutputS2xD(16)(0);
  VNStageIntLLRInputS2xD(102)(0) <= CNStageIntLLROutputS2xD(16)(1);
  VNStageIntLLRInputS2xD(166)(0) <= CNStageIntLLROutputS2xD(16)(2);
  VNStageIntLLRInputS2xD(230)(0) <= CNStageIntLLROutputS2xD(16)(3);
  VNStageIntLLRInputS2xD(294)(0) <= CNStageIntLLROutputS2xD(16)(4);
  VNStageIntLLRInputS2xD(358)(0) <= CNStageIntLLROutputS2xD(16)(5);
  VNStageIntLLRInputS2xD(37)(0) <= CNStageIntLLROutputS2xD(17)(0);
  VNStageIntLLRInputS2xD(101)(0) <= CNStageIntLLROutputS2xD(17)(1);
  VNStageIntLLRInputS2xD(165)(0) <= CNStageIntLLROutputS2xD(17)(2);
  VNStageIntLLRInputS2xD(229)(0) <= CNStageIntLLROutputS2xD(17)(3);
  VNStageIntLLRInputS2xD(293)(0) <= CNStageIntLLROutputS2xD(17)(4);
  VNStageIntLLRInputS2xD(357)(0) <= CNStageIntLLROutputS2xD(17)(5);
  VNStageIntLLRInputS2xD(36)(0) <= CNStageIntLLROutputS2xD(18)(0);
  VNStageIntLLRInputS2xD(100)(0) <= CNStageIntLLROutputS2xD(18)(1);
  VNStageIntLLRInputS2xD(164)(0) <= CNStageIntLLROutputS2xD(18)(2);
  VNStageIntLLRInputS2xD(228)(0) <= CNStageIntLLROutputS2xD(18)(3);
  VNStageIntLLRInputS2xD(292)(0) <= CNStageIntLLROutputS2xD(18)(4);
  VNStageIntLLRInputS2xD(356)(0) <= CNStageIntLLROutputS2xD(18)(5);
  VNStageIntLLRInputS2xD(35)(0) <= CNStageIntLLROutputS2xD(19)(0);
  VNStageIntLLRInputS2xD(99)(0) <= CNStageIntLLROutputS2xD(19)(1);
  VNStageIntLLRInputS2xD(163)(0) <= CNStageIntLLROutputS2xD(19)(2);
  VNStageIntLLRInputS2xD(227)(0) <= CNStageIntLLROutputS2xD(19)(3);
  VNStageIntLLRInputS2xD(291)(0) <= CNStageIntLLROutputS2xD(19)(4);
  VNStageIntLLRInputS2xD(355)(0) <= CNStageIntLLROutputS2xD(19)(5);
  VNStageIntLLRInputS2xD(34)(0) <= CNStageIntLLROutputS2xD(20)(0);
  VNStageIntLLRInputS2xD(98)(0) <= CNStageIntLLROutputS2xD(20)(1);
  VNStageIntLLRInputS2xD(162)(0) <= CNStageIntLLROutputS2xD(20)(2);
  VNStageIntLLRInputS2xD(226)(0) <= CNStageIntLLROutputS2xD(20)(3);
  VNStageIntLLRInputS2xD(290)(0) <= CNStageIntLLROutputS2xD(20)(4);
  VNStageIntLLRInputS2xD(354)(0) <= CNStageIntLLROutputS2xD(20)(5);
  VNStageIntLLRInputS2xD(33)(0) <= CNStageIntLLROutputS2xD(21)(0);
  VNStageIntLLRInputS2xD(97)(0) <= CNStageIntLLROutputS2xD(21)(1);
  VNStageIntLLRInputS2xD(161)(0) <= CNStageIntLLROutputS2xD(21)(2);
  VNStageIntLLRInputS2xD(225)(0) <= CNStageIntLLROutputS2xD(21)(3);
  VNStageIntLLRInputS2xD(289)(0) <= CNStageIntLLROutputS2xD(21)(4);
  VNStageIntLLRInputS2xD(353)(0) <= CNStageIntLLROutputS2xD(21)(5);
  VNStageIntLLRInputS2xD(32)(0) <= CNStageIntLLROutputS2xD(22)(0);
  VNStageIntLLRInputS2xD(96)(0) <= CNStageIntLLROutputS2xD(22)(1);
  VNStageIntLLRInputS2xD(160)(0) <= CNStageIntLLROutputS2xD(22)(2);
  VNStageIntLLRInputS2xD(224)(0) <= CNStageIntLLROutputS2xD(22)(3);
  VNStageIntLLRInputS2xD(288)(0) <= CNStageIntLLROutputS2xD(22)(4);
  VNStageIntLLRInputS2xD(352)(0) <= CNStageIntLLROutputS2xD(22)(5);
  VNStageIntLLRInputS2xD(31)(0) <= CNStageIntLLROutputS2xD(23)(0);
  VNStageIntLLRInputS2xD(95)(0) <= CNStageIntLLROutputS2xD(23)(1);
  VNStageIntLLRInputS2xD(159)(0) <= CNStageIntLLROutputS2xD(23)(2);
  VNStageIntLLRInputS2xD(223)(0) <= CNStageIntLLROutputS2xD(23)(3);
  VNStageIntLLRInputS2xD(287)(0) <= CNStageIntLLROutputS2xD(23)(4);
  VNStageIntLLRInputS2xD(351)(0) <= CNStageIntLLROutputS2xD(23)(5);
  VNStageIntLLRInputS2xD(30)(0) <= CNStageIntLLROutputS2xD(24)(0);
  VNStageIntLLRInputS2xD(94)(0) <= CNStageIntLLROutputS2xD(24)(1);
  VNStageIntLLRInputS2xD(158)(0) <= CNStageIntLLROutputS2xD(24)(2);
  VNStageIntLLRInputS2xD(222)(0) <= CNStageIntLLROutputS2xD(24)(3);
  VNStageIntLLRInputS2xD(286)(0) <= CNStageIntLLROutputS2xD(24)(4);
  VNStageIntLLRInputS2xD(350)(0) <= CNStageIntLLROutputS2xD(24)(5);
  VNStageIntLLRInputS2xD(29)(0) <= CNStageIntLLROutputS2xD(25)(0);
  VNStageIntLLRInputS2xD(93)(0) <= CNStageIntLLROutputS2xD(25)(1);
  VNStageIntLLRInputS2xD(157)(0) <= CNStageIntLLROutputS2xD(25)(2);
  VNStageIntLLRInputS2xD(221)(0) <= CNStageIntLLROutputS2xD(25)(3);
  VNStageIntLLRInputS2xD(285)(0) <= CNStageIntLLROutputS2xD(25)(4);
  VNStageIntLLRInputS2xD(349)(0) <= CNStageIntLLROutputS2xD(25)(5);
  VNStageIntLLRInputS2xD(28)(0) <= CNStageIntLLROutputS2xD(26)(0);
  VNStageIntLLRInputS2xD(92)(0) <= CNStageIntLLROutputS2xD(26)(1);
  VNStageIntLLRInputS2xD(156)(0) <= CNStageIntLLROutputS2xD(26)(2);
  VNStageIntLLRInputS2xD(220)(0) <= CNStageIntLLROutputS2xD(26)(3);
  VNStageIntLLRInputS2xD(284)(0) <= CNStageIntLLROutputS2xD(26)(4);
  VNStageIntLLRInputS2xD(348)(0) <= CNStageIntLLROutputS2xD(26)(5);
  VNStageIntLLRInputS2xD(27)(0) <= CNStageIntLLROutputS2xD(27)(0);
  VNStageIntLLRInputS2xD(91)(0) <= CNStageIntLLROutputS2xD(27)(1);
  VNStageIntLLRInputS2xD(155)(0) <= CNStageIntLLROutputS2xD(27)(2);
  VNStageIntLLRInputS2xD(219)(0) <= CNStageIntLLROutputS2xD(27)(3);
  VNStageIntLLRInputS2xD(283)(0) <= CNStageIntLLROutputS2xD(27)(4);
  VNStageIntLLRInputS2xD(347)(0) <= CNStageIntLLROutputS2xD(27)(5);
  VNStageIntLLRInputS2xD(26)(0) <= CNStageIntLLROutputS2xD(28)(0);
  VNStageIntLLRInputS2xD(90)(0) <= CNStageIntLLROutputS2xD(28)(1);
  VNStageIntLLRInputS2xD(154)(0) <= CNStageIntLLROutputS2xD(28)(2);
  VNStageIntLLRInputS2xD(218)(0) <= CNStageIntLLROutputS2xD(28)(3);
  VNStageIntLLRInputS2xD(282)(0) <= CNStageIntLLROutputS2xD(28)(4);
  VNStageIntLLRInputS2xD(346)(0) <= CNStageIntLLROutputS2xD(28)(5);
  VNStageIntLLRInputS2xD(25)(0) <= CNStageIntLLROutputS2xD(29)(0);
  VNStageIntLLRInputS2xD(89)(0) <= CNStageIntLLROutputS2xD(29)(1);
  VNStageIntLLRInputS2xD(153)(0) <= CNStageIntLLROutputS2xD(29)(2);
  VNStageIntLLRInputS2xD(217)(0) <= CNStageIntLLROutputS2xD(29)(3);
  VNStageIntLLRInputS2xD(281)(0) <= CNStageIntLLROutputS2xD(29)(4);
  VNStageIntLLRInputS2xD(345)(0) <= CNStageIntLLROutputS2xD(29)(5);
  VNStageIntLLRInputS2xD(24)(0) <= CNStageIntLLROutputS2xD(30)(0);
  VNStageIntLLRInputS2xD(88)(0) <= CNStageIntLLROutputS2xD(30)(1);
  VNStageIntLLRInputS2xD(152)(0) <= CNStageIntLLROutputS2xD(30)(2);
  VNStageIntLLRInputS2xD(216)(0) <= CNStageIntLLROutputS2xD(30)(3);
  VNStageIntLLRInputS2xD(280)(0) <= CNStageIntLLROutputS2xD(30)(4);
  VNStageIntLLRInputS2xD(344)(0) <= CNStageIntLLROutputS2xD(30)(5);
  VNStageIntLLRInputS2xD(23)(0) <= CNStageIntLLROutputS2xD(31)(0);
  VNStageIntLLRInputS2xD(87)(0) <= CNStageIntLLROutputS2xD(31)(1);
  VNStageIntLLRInputS2xD(151)(0) <= CNStageIntLLROutputS2xD(31)(2);
  VNStageIntLLRInputS2xD(215)(0) <= CNStageIntLLROutputS2xD(31)(3);
  VNStageIntLLRInputS2xD(279)(0) <= CNStageIntLLROutputS2xD(31)(4);
  VNStageIntLLRInputS2xD(343)(0) <= CNStageIntLLROutputS2xD(31)(5);
  VNStageIntLLRInputS2xD(22)(0) <= CNStageIntLLROutputS2xD(32)(0);
  VNStageIntLLRInputS2xD(86)(0) <= CNStageIntLLROutputS2xD(32)(1);
  VNStageIntLLRInputS2xD(150)(0) <= CNStageIntLLROutputS2xD(32)(2);
  VNStageIntLLRInputS2xD(214)(0) <= CNStageIntLLROutputS2xD(32)(3);
  VNStageIntLLRInputS2xD(278)(0) <= CNStageIntLLROutputS2xD(32)(4);
  VNStageIntLLRInputS2xD(342)(0) <= CNStageIntLLROutputS2xD(32)(5);
  VNStageIntLLRInputS2xD(21)(0) <= CNStageIntLLROutputS2xD(33)(0);
  VNStageIntLLRInputS2xD(85)(0) <= CNStageIntLLROutputS2xD(33)(1);
  VNStageIntLLRInputS2xD(149)(0) <= CNStageIntLLROutputS2xD(33)(2);
  VNStageIntLLRInputS2xD(213)(0) <= CNStageIntLLROutputS2xD(33)(3);
  VNStageIntLLRInputS2xD(277)(0) <= CNStageIntLLROutputS2xD(33)(4);
  VNStageIntLLRInputS2xD(341)(0) <= CNStageIntLLROutputS2xD(33)(5);
  VNStageIntLLRInputS2xD(20)(0) <= CNStageIntLLROutputS2xD(34)(0);
  VNStageIntLLRInputS2xD(84)(0) <= CNStageIntLLROutputS2xD(34)(1);
  VNStageIntLLRInputS2xD(148)(0) <= CNStageIntLLROutputS2xD(34)(2);
  VNStageIntLLRInputS2xD(212)(0) <= CNStageIntLLROutputS2xD(34)(3);
  VNStageIntLLRInputS2xD(276)(0) <= CNStageIntLLROutputS2xD(34)(4);
  VNStageIntLLRInputS2xD(340)(0) <= CNStageIntLLROutputS2xD(34)(5);
  VNStageIntLLRInputS2xD(19)(0) <= CNStageIntLLROutputS2xD(35)(0);
  VNStageIntLLRInputS2xD(83)(0) <= CNStageIntLLROutputS2xD(35)(1);
  VNStageIntLLRInputS2xD(147)(0) <= CNStageIntLLROutputS2xD(35)(2);
  VNStageIntLLRInputS2xD(211)(0) <= CNStageIntLLROutputS2xD(35)(3);
  VNStageIntLLRInputS2xD(275)(0) <= CNStageIntLLROutputS2xD(35)(4);
  VNStageIntLLRInputS2xD(339)(0) <= CNStageIntLLROutputS2xD(35)(5);
  VNStageIntLLRInputS2xD(18)(0) <= CNStageIntLLROutputS2xD(36)(0);
  VNStageIntLLRInputS2xD(82)(0) <= CNStageIntLLROutputS2xD(36)(1);
  VNStageIntLLRInputS2xD(146)(0) <= CNStageIntLLROutputS2xD(36)(2);
  VNStageIntLLRInputS2xD(210)(0) <= CNStageIntLLROutputS2xD(36)(3);
  VNStageIntLLRInputS2xD(274)(0) <= CNStageIntLLROutputS2xD(36)(4);
  VNStageIntLLRInputS2xD(338)(0) <= CNStageIntLLROutputS2xD(36)(5);
  VNStageIntLLRInputS2xD(17)(0) <= CNStageIntLLROutputS2xD(37)(0);
  VNStageIntLLRInputS2xD(81)(0) <= CNStageIntLLROutputS2xD(37)(1);
  VNStageIntLLRInputS2xD(145)(0) <= CNStageIntLLROutputS2xD(37)(2);
  VNStageIntLLRInputS2xD(209)(0) <= CNStageIntLLROutputS2xD(37)(3);
  VNStageIntLLRInputS2xD(273)(0) <= CNStageIntLLROutputS2xD(37)(4);
  VNStageIntLLRInputS2xD(337)(0) <= CNStageIntLLROutputS2xD(37)(5);
  VNStageIntLLRInputS2xD(16)(0) <= CNStageIntLLROutputS2xD(38)(0);
  VNStageIntLLRInputS2xD(80)(0) <= CNStageIntLLROutputS2xD(38)(1);
  VNStageIntLLRInputS2xD(144)(0) <= CNStageIntLLROutputS2xD(38)(2);
  VNStageIntLLRInputS2xD(208)(0) <= CNStageIntLLROutputS2xD(38)(3);
  VNStageIntLLRInputS2xD(272)(0) <= CNStageIntLLROutputS2xD(38)(4);
  VNStageIntLLRInputS2xD(336)(0) <= CNStageIntLLROutputS2xD(38)(5);
  VNStageIntLLRInputS2xD(15)(0) <= CNStageIntLLROutputS2xD(39)(0);
  VNStageIntLLRInputS2xD(79)(0) <= CNStageIntLLROutputS2xD(39)(1);
  VNStageIntLLRInputS2xD(143)(0) <= CNStageIntLLROutputS2xD(39)(2);
  VNStageIntLLRInputS2xD(207)(0) <= CNStageIntLLROutputS2xD(39)(3);
  VNStageIntLLRInputS2xD(271)(0) <= CNStageIntLLROutputS2xD(39)(4);
  VNStageIntLLRInputS2xD(335)(0) <= CNStageIntLLROutputS2xD(39)(5);
  VNStageIntLLRInputS2xD(14)(0) <= CNStageIntLLROutputS2xD(40)(0);
  VNStageIntLLRInputS2xD(78)(0) <= CNStageIntLLROutputS2xD(40)(1);
  VNStageIntLLRInputS2xD(142)(0) <= CNStageIntLLROutputS2xD(40)(2);
  VNStageIntLLRInputS2xD(206)(0) <= CNStageIntLLROutputS2xD(40)(3);
  VNStageIntLLRInputS2xD(270)(0) <= CNStageIntLLROutputS2xD(40)(4);
  VNStageIntLLRInputS2xD(334)(0) <= CNStageIntLLROutputS2xD(40)(5);
  VNStageIntLLRInputS2xD(12)(0) <= CNStageIntLLROutputS2xD(41)(0);
  VNStageIntLLRInputS2xD(76)(0) <= CNStageIntLLROutputS2xD(41)(1);
  VNStageIntLLRInputS2xD(140)(0) <= CNStageIntLLROutputS2xD(41)(2);
  VNStageIntLLRInputS2xD(204)(0) <= CNStageIntLLROutputS2xD(41)(3);
  VNStageIntLLRInputS2xD(268)(0) <= CNStageIntLLROutputS2xD(41)(4);
  VNStageIntLLRInputS2xD(332)(0) <= CNStageIntLLROutputS2xD(41)(5);
  VNStageIntLLRInputS2xD(11)(0) <= CNStageIntLLROutputS2xD(42)(0);
  VNStageIntLLRInputS2xD(75)(0) <= CNStageIntLLROutputS2xD(42)(1);
  VNStageIntLLRInputS2xD(139)(0) <= CNStageIntLLROutputS2xD(42)(2);
  VNStageIntLLRInputS2xD(203)(0) <= CNStageIntLLROutputS2xD(42)(3);
  VNStageIntLLRInputS2xD(267)(0) <= CNStageIntLLROutputS2xD(42)(4);
  VNStageIntLLRInputS2xD(331)(0) <= CNStageIntLLROutputS2xD(42)(5);
  VNStageIntLLRInputS2xD(10)(0) <= CNStageIntLLROutputS2xD(43)(0);
  VNStageIntLLRInputS2xD(74)(0) <= CNStageIntLLROutputS2xD(43)(1);
  VNStageIntLLRInputS2xD(138)(0) <= CNStageIntLLROutputS2xD(43)(2);
  VNStageIntLLRInputS2xD(202)(0) <= CNStageIntLLROutputS2xD(43)(3);
  VNStageIntLLRInputS2xD(266)(0) <= CNStageIntLLROutputS2xD(43)(4);
  VNStageIntLLRInputS2xD(330)(0) <= CNStageIntLLROutputS2xD(43)(5);
  VNStageIntLLRInputS2xD(9)(0) <= CNStageIntLLROutputS2xD(44)(0);
  VNStageIntLLRInputS2xD(73)(0) <= CNStageIntLLROutputS2xD(44)(1);
  VNStageIntLLRInputS2xD(137)(0) <= CNStageIntLLROutputS2xD(44)(2);
  VNStageIntLLRInputS2xD(201)(0) <= CNStageIntLLROutputS2xD(44)(3);
  VNStageIntLLRInputS2xD(265)(0) <= CNStageIntLLROutputS2xD(44)(4);
  VNStageIntLLRInputS2xD(329)(0) <= CNStageIntLLROutputS2xD(44)(5);
  VNStageIntLLRInputS2xD(8)(0) <= CNStageIntLLROutputS2xD(45)(0);
  VNStageIntLLRInputS2xD(72)(0) <= CNStageIntLLROutputS2xD(45)(1);
  VNStageIntLLRInputS2xD(136)(0) <= CNStageIntLLROutputS2xD(45)(2);
  VNStageIntLLRInputS2xD(200)(0) <= CNStageIntLLROutputS2xD(45)(3);
  VNStageIntLLRInputS2xD(264)(0) <= CNStageIntLLROutputS2xD(45)(4);
  VNStageIntLLRInputS2xD(328)(0) <= CNStageIntLLROutputS2xD(45)(5);
  VNStageIntLLRInputS2xD(7)(0) <= CNStageIntLLROutputS2xD(46)(0);
  VNStageIntLLRInputS2xD(71)(0) <= CNStageIntLLROutputS2xD(46)(1);
  VNStageIntLLRInputS2xD(135)(0) <= CNStageIntLLROutputS2xD(46)(2);
  VNStageIntLLRInputS2xD(199)(0) <= CNStageIntLLROutputS2xD(46)(3);
  VNStageIntLLRInputS2xD(263)(0) <= CNStageIntLLROutputS2xD(46)(4);
  VNStageIntLLRInputS2xD(327)(0) <= CNStageIntLLROutputS2xD(46)(5);
  VNStageIntLLRInputS2xD(6)(0) <= CNStageIntLLROutputS2xD(47)(0);
  VNStageIntLLRInputS2xD(70)(0) <= CNStageIntLLROutputS2xD(47)(1);
  VNStageIntLLRInputS2xD(134)(0) <= CNStageIntLLROutputS2xD(47)(2);
  VNStageIntLLRInputS2xD(198)(0) <= CNStageIntLLROutputS2xD(47)(3);
  VNStageIntLLRInputS2xD(262)(0) <= CNStageIntLLROutputS2xD(47)(4);
  VNStageIntLLRInputS2xD(326)(0) <= CNStageIntLLROutputS2xD(47)(5);
  VNStageIntLLRInputS2xD(5)(0) <= CNStageIntLLROutputS2xD(48)(0);
  VNStageIntLLRInputS2xD(69)(0) <= CNStageIntLLROutputS2xD(48)(1);
  VNStageIntLLRInputS2xD(133)(0) <= CNStageIntLLROutputS2xD(48)(2);
  VNStageIntLLRInputS2xD(197)(0) <= CNStageIntLLROutputS2xD(48)(3);
  VNStageIntLLRInputS2xD(261)(0) <= CNStageIntLLROutputS2xD(48)(4);
  VNStageIntLLRInputS2xD(325)(0) <= CNStageIntLLROutputS2xD(48)(5);
  VNStageIntLLRInputS2xD(4)(0) <= CNStageIntLLROutputS2xD(49)(0);
  VNStageIntLLRInputS2xD(68)(0) <= CNStageIntLLROutputS2xD(49)(1);
  VNStageIntLLRInputS2xD(132)(0) <= CNStageIntLLROutputS2xD(49)(2);
  VNStageIntLLRInputS2xD(196)(0) <= CNStageIntLLROutputS2xD(49)(3);
  VNStageIntLLRInputS2xD(260)(0) <= CNStageIntLLROutputS2xD(49)(4);
  VNStageIntLLRInputS2xD(324)(0) <= CNStageIntLLROutputS2xD(49)(5);
  VNStageIntLLRInputS2xD(2)(0) <= CNStageIntLLROutputS2xD(50)(0);
  VNStageIntLLRInputS2xD(66)(0) <= CNStageIntLLROutputS2xD(50)(1);
  VNStageIntLLRInputS2xD(130)(0) <= CNStageIntLLROutputS2xD(50)(2);
  VNStageIntLLRInputS2xD(194)(0) <= CNStageIntLLROutputS2xD(50)(3);
  VNStageIntLLRInputS2xD(258)(0) <= CNStageIntLLROutputS2xD(50)(4);
  VNStageIntLLRInputS2xD(322)(0) <= CNStageIntLLROutputS2xD(50)(5);
  VNStageIntLLRInputS2xD(1)(0) <= CNStageIntLLROutputS2xD(51)(0);
  VNStageIntLLRInputS2xD(65)(0) <= CNStageIntLLROutputS2xD(51)(1);
  VNStageIntLLRInputS2xD(129)(0) <= CNStageIntLLROutputS2xD(51)(2);
  VNStageIntLLRInputS2xD(193)(0) <= CNStageIntLLROutputS2xD(51)(3);
  VNStageIntLLRInputS2xD(257)(0) <= CNStageIntLLROutputS2xD(51)(4);
  VNStageIntLLRInputS2xD(321)(0) <= CNStageIntLLROutputS2xD(51)(5);
  VNStageIntLLRInputS2xD(63)(0) <= CNStageIntLLROutputS2xD(52)(0);
  VNStageIntLLRInputS2xD(127)(0) <= CNStageIntLLROutputS2xD(52)(1);
  VNStageIntLLRInputS2xD(191)(0) <= CNStageIntLLROutputS2xD(52)(2);
  VNStageIntLLRInputS2xD(255)(0) <= CNStageIntLLROutputS2xD(52)(3);
  VNStageIntLLRInputS2xD(319)(0) <= CNStageIntLLROutputS2xD(52)(4);
  VNStageIntLLRInputS2xD(383)(0) <= CNStageIntLLROutputS2xD(52)(5);
  VNStageIntLLRInputS2xD(0)(0) <= CNStageIntLLROutputS2xD(53)(0);
  VNStageIntLLRInputS2xD(64)(0) <= CNStageIntLLROutputS2xD(53)(1);
  VNStageIntLLRInputS2xD(128)(0) <= CNStageIntLLROutputS2xD(53)(2);
  VNStageIntLLRInputS2xD(192)(0) <= CNStageIntLLROutputS2xD(53)(3);
  VNStageIntLLRInputS2xD(256)(0) <= CNStageIntLLROutputS2xD(53)(4);
  VNStageIntLLRInputS2xD(320)(0) <= CNStageIntLLROutputS2xD(53)(5);
  VNStageIntLLRInputS2xD(42)(1) <= CNStageIntLLROutputS2xD(54)(0);
  VNStageIntLLRInputS2xD(112)(1) <= CNStageIntLLROutputS2xD(54)(1);
  VNStageIntLLRInputS2xD(182)(1) <= CNStageIntLLROutputS2xD(54)(2);
  VNStageIntLLRInputS2xD(203)(1) <= CNStageIntLLROutputS2xD(54)(3);
  VNStageIntLLRInputS2xD(259)(0) <= CNStageIntLLROutputS2xD(54)(4);
  VNStageIntLLRInputS2xD(361)(1) <= CNStageIntLLROutputS2xD(54)(5);
  VNStageIntLLRInputS2xD(41)(1) <= CNStageIntLLROutputS2xD(55)(0);
  VNStageIntLLRInputS2xD(117)(1) <= CNStageIntLLROutputS2xD(55)(1);
  VNStageIntLLRInputS2xD(138)(1) <= CNStageIntLLROutputS2xD(55)(2);
  VNStageIntLLRInputS2xD(194)(1) <= CNStageIntLLROutputS2xD(55)(3);
  VNStageIntLLRInputS2xD(296)(1) <= CNStageIntLLROutputS2xD(55)(4);
  VNStageIntLLRInputS2xD(362)(1) <= CNStageIntLLROutputS2xD(55)(5);
  VNStageIntLLRInputS2xD(40)(1) <= CNStageIntLLROutputS2xD(56)(0);
  VNStageIntLLRInputS2xD(73)(1) <= CNStageIntLLROutputS2xD(56)(1);
  VNStageIntLLRInputS2xD(129)(1) <= CNStageIntLLROutputS2xD(56)(2);
  VNStageIntLLRInputS2xD(231)(1) <= CNStageIntLLROutputS2xD(56)(3);
  VNStageIntLLRInputS2xD(297)(1) <= CNStageIntLLROutputS2xD(56)(4);
  VNStageIntLLRInputS2xD(323)(0) <= CNStageIntLLROutputS2xD(56)(5);
  VNStageIntLLRInputS2xD(39)(1) <= CNStageIntLLROutputS2xD(57)(0);
  VNStageIntLLRInputS2xD(127)(1) <= CNStageIntLLROutputS2xD(57)(1);
  VNStageIntLLRInputS2xD(166)(1) <= CNStageIntLLROutputS2xD(57)(2);
  VNStageIntLLRInputS2xD(232)(1) <= CNStageIntLLROutputS2xD(57)(3);
  VNStageIntLLRInputS2xD(258)(1) <= CNStageIntLLROutputS2xD(57)(4);
  VNStageIntLLRInputS2xD(344)(1) <= CNStageIntLLROutputS2xD(57)(5);
  VNStageIntLLRInputS2xD(38)(1) <= CNStageIntLLROutputS2xD(58)(0);
  VNStageIntLLRInputS2xD(101)(1) <= CNStageIntLLROutputS2xD(58)(1);
  VNStageIntLLRInputS2xD(167)(1) <= CNStageIntLLROutputS2xD(58)(2);
  VNStageIntLLRInputS2xD(193)(1) <= CNStageIntLLROutputS2xD(58)(3);
  VNStageIntLLRInputS2xD(279)(1) <= CNStageIntLLROutputS2xD(58)(4);
  VNStageIntLLRInputS2xD(340)(1) <= CNStageIntLLROutputS2xD(58)(5);
  VNStageIntLLRInputS2xD(37)(1) <= CNStageIntLLROutputS2xD(59)(0);
  VNStageIntLLRInputS2xD(102)(1) <= CNStageIntLLROutputS2xD(59)(1);
  VNStageIntLLRInputS2xD(191)(1) <= CNStageIntLLROutputS2xD(59)(2);
  VNStageIntLLRInputS2xD(214)(1) <= CNStageIntLLROutputS2xD(59)(3);
  VNStageIntLLRInputS2xD(275)(1) <= CNStageIntLLROutputS2xD(59)(4);
  VNStageIntLLRInputS2xD(355)(1) <= CNStageIntLLROutputS2xD(59)(5);
  VNStageIntLLRInputS2xD(36)(1) <= CNStageIntLLROutputS2xD(60)(0);
  VNStageIntLLRInputS2xD(126)(0) <= CNStageIntLLROutputS2xD(60)(1);
  VNStageIntLLRInputS2xD(149)(1) <= CNStageIntLLROutputS2xD(60)(2);
  VNStageIntLLRInputS2xD(210)(1) <= CNStageIntLLROutputS2xD(60)(3);
  VNStageIntLLRInputS2xD(290)(1) <= CNStageIntLLROutputS2xD(60)(4);
  VNStageIntLLRInputS2xD(381)(0) <= CNStageIntLLROutputS2xD(60)(5);
  VNStageIntLLRInputS2xD(35)(1) <= CNStageIntLLROutputS2xD(61)(0);
  VNStageIntLLRInputS2xD(84)(1) <= CNStageIntLLROutputS2xD(61)(1);
  VNStageIntLLRInputS2xD(145)(1) <= CNStageIntLLROutputS2xD(61)(2);
  VNStageIntLLRInputS2xD(225)(1) <= CNStageIntLLROutputS2xD(61)(3);
  VNStageIntLLRInputS2xD(316)(0) <= CNStageIntLLROutputS2xD(61)(4);
  VNStageIntLLRInputS2xD(357)(1) <= CNStageIntLLROutputS2xD(61)(5);
  VNStageIntLLRInputS2xD(34)(1) <= CNStageIntLLROutputS2xD(62)(0);
  VNStageIntLLRInputS2xD(80)(1) <= CNStageIntLLROutputS2xD(62)(1);
  VNStageIntLLRInputS2xD(160)(1) <= CNStageIntLLROutputS2xD(62)(2);
  VNStageIntLLRInputS2xD(251)(0) <= CNStageIntLLROutputS2xD(62)(3);
  VNStageIntLLRInputS2xD(292)(1) <= CNStageIntLLROutputS2xD(62)(4);
  VNStageIntLLRInputS2xD(326)(1) <= CNStageIntLLROutputS2xD(62)(5);
  VNStageIntLLRInputS2xD(33)(1) <= CNStageIntLLROutputS2xD(63)(0);
  VNStageIntLLRInputS2xD(95)(1) <= CNStageIntLLROutputS2xD(63)(1);
  VNStageIntLLRInputS2xD(186)(0) <= CNStageIntLLROutputS2xD(63)(2);
  VNStageIntLLRInputS2xD(227)(1) <= CNStageIntLLROutputS2xD(63)(3);
  VNStageIntLLRInputS2xD(261)(1) <= CNStageIntLLROutputS2xD(63)(4);
  VNStageIntLLRInputS2xD(342)(1) <= CNStageIntLLROutputS2xD(63)(5);
  VNStageIntLLRInputS2xD(32)(1) <= CNStageIntLLROutputS2xD(64)(0);
  VNStageIntLLRInputS2xD(121)(0) <= CNStageIntLLROutputS2xD(64)(1);
  VNStageIntLLRInputS2xD(162)(1) <= CNStageIntLLROutputS2xD(64)(2);
  VNStageIntLLRInputS2xD(196)(1) <= CNStageIntLLROutputS2xD(64)(3);
  VNStageIntLLRInputS2xD(277)(1) <= CNStageIntLLROutputS2xD(64)(4);
  VNStageIntLLRInputS2xD(375)(1) <= CNStageIntLLROutputS2xD(64)(5);
  VNStageIntLLRInputS2xD(31)(1) <= CNStageIntLLROutputS2xD(65)(0);
  VNStageIntLLRInputS2xD(97)(1) <= CNStageIntLLROutputS2xD(65)(1);
  VNStageIntLLRInputS2xD(131)(0) <= CNStageIntLLROutputS2xD(65)(2);
  VNStageIntLLRInputS2xD(212)(1) <= CNStageIntLLROutputS2xD(65)(3);
  VNStageIntLLRInputS2xD(310)(1) <= CNStageIntLLROutputS2xD(65)(4);
  VNStageIntLLRInputS2xD(321)(1) <= CNStageIntLLROutputS2xD(65)(5);
  VNStageIntLLRInputS2xD(30)(1) <= CNStageIntLLROutputS2xD(66)(0);
  VNStageIntLLRInputS2xD(66)(1) <= CNStageIntLLROutputS2xD(66)(1);
  VNStageIntLLRInputS2xD(147)(1) <= CNStageIntLLROutputS2xD(66)(2);
  VNStageIntLLRInputS2xD(245)(1) <= CNStageIntLLROutputS2xD(66)(3);
  VNStageIntLLRInputS2xD(319)(1) <= CNStageIntLLROutputS2xD(66)(4);
  VNStageIntLLRInputS2xD(334)(1) <= CNStageIntLLROutputS2xD(66)(5);
  VNStageIntLLRInputS2xD(29)(1) <= CNStageIntLLROutputS2xD(67)(0);
  VNStageIntLLRInputS2xD(82)(1) <= CNStageIntLLROutputS2xD(67)(1);
  VNStageIntLLRInputS2xD(180)(0) <= CNStageIntLLROutputS2xD(67)(2);
  VNStageIntLLRInputS2xD(254)(0) <= CNStageIntLLROutputS2xD(67)(3);
  VNStageIntLLRInputS2xD(269)(0) <= CNStageIntLLROutputS2xD(67)(4);
  VNStageIntLLRInputS2xD(376)(1) <= CNStageIntLLROutputS2xD(67)(5);
  VNStageIntLLRInputS2xD(28)(1) <= CNStageIntLLROutputS2xD(68)(0);
  VNStageIntLLRInputS2xD(115)(1) <= CNStageIntLLROutputS2xD(68)(1);
  VNStageIntLLRInputS2xD(189)(0) <= CNStageIntLLROutputS2xD(68)(2);
  VNStageIntLLRInputS2xD(204)(1) <= CNStageIntLLROutputS2xD(68)(3);
  VNStageIntLLRInputS2xD(311)(1) <= CNStageIntLLROutputS2xD(68)(4);
  VNStageIntLLRInputS2xD(341)(1) <= CNStageIntLLROutputS2xD(68)(5);
  VNStageIntLLRInputS2xD(27)(1) <= CNStageIntLLROutputS2xD(69)(0);
  VNStageIntLLRInputS2xD(124)(0) <= CNStageIntLLROutputS2xD(69)(1);
  VNStageIntLLRInputS2xD(139)(1) <= CNStageIntLLROutputS2xD(69)(2);
  VNStageIntLLRInputS2xD(246)(1) <= CNStageIntLLROutputS2xD(69)(3);
  VNStageIntLLRInputS2xD(276)(1) <= CNStageIntLLROutputS2xD(69)(4);
  VNStageIntLLRInputS2xD(343)(1) <= CNStageIntLLROutputS2xD(69)(5);
  VNStageIntLLRInputS2xD(26)(1) <= CNStageIntLLROutputS2xD(70)(0);
  VNStageIntLLRInputS2xD(74)(1) <= CNStageIntLLROutputS2xD(70)(1);
  VNStageIntLLRInputS2xD(181)(1) <= CNStageIntLLROutputS2xD(70)(2);
  VNStageIntLLRInputS2xD(211)(1) <= CNStageIntLLROutputS2xD(70)(3);
  VNStageIntLLRInputS2xD(278)(1) <= CNStageIntLLROutputS2xD(70)(4);
  VNStageIntLLRInputS2xD(325)(1) <= CNStageIntLLROutputS2xD(70)(5);
  VNStageIntLLRInputS2xD(25)(1) <= CNStageIntLLROutputS2xD(71)(0);
  VNStageIntLLRInputS2xD(116)(0) <= CNStageIntLLROutputS2xD(71)(1);
  VNStageIntLLRInputS2xD(146)(1) <= CNStageIntLLROutputS2xD(71)(2);
  VNStageIntLLRInputS2xD(213)(1) <= CNStageIntLLROutputS2xD(71)(3);
  VNStageIntLLRInputS2xD(260)(1) <= CNStageIntLLROutputS2xD(71)(4);
  VNStageIntLLRInputS2xD(332)(1) <= CNStageIntLLROutputS2xD(71)(5);
  VNStageIntLLRInputS2xD(24)(1) <= CNStageIntLLROutputS2xD(72)(0);
  VNStageIntLLRInputS2xD(81)(1) <= CNStageIntLLROutputS2xD(72)(1);
  VNStageIntLLRInputS2xD(148)(1) <= CNStageIntLLROutputS2xD(72)(2);
  VNStageIntLLRInputS2xD(195)(0) <= CNStageIntLLROutputS2xD(72)(3);
  VNStageIntLLRInputS2xD(267)(1) <= CNStageIntLLROutputS2xD(72)(4);
  VNStageIntLLRInputS2xD(359)(1) <= CNStageIntLLROutputS2xD(72)(5);
  VNStageIntLLRInputS2xD(23)(1) <= CNStageIntLLROutputS2xD(73)(0);
  VNStageIntLLRInputS2xD(83)(1) <= CNStageIntLLROutputS2xD(73)(1);
  VNStageIntLLRInputS2xD(130)(1) <= CNStageIntLLROutputS2xD(73)(2);
  VNStageIntLLRInputS2xD(202)(1) <= CNStageIntLLROutputS2xD(73)(3);
  VNStageIntLLRInputS2xD(294)(1) <= CNStageIntLLROutputS2xD(73)(4);
  VNStageIntLLRInputS2xD(347)(1) <= CNStageIntLLROutputS2xD(73)(5);
  VNStageIntLLRInputS2xD(22)(1) <= CNStageIntLLROutputS2xD(74)(0);
  VNStageIntLLRInputS2xD(65)(1) <= CNStageIntLLROutputS2xD(74)(1);
  VNStageIntLLRInputS2xD(137)(1) <= CNStageIntLLROutputS2xD(74)(2);
  VNStageIntLLRInputS2xD(229)(1) <= CNStageIntLLROutputS2xD(74)(3);
  VNStageIntLLRInputS2xD(282)(1) <= CNStageIntLLROutputS2xD(74)(4);
  VNStageIntLLRInputS2xD(353)(1) <= CNStageIntLLROutputS2xD(74)(5);
  VNStageIntLLRInputS2xD(21)(1) <= CNStageIntLLROutputS2xD(75)(0);
  VNStageIntLLRInputS2xD(72)(1) <= CNStageIntLLROutputS2xD(75)(1);
  VNStageIntLLRInputS2xD(164)(1) <= CNStageIntLLROutputS2xD(75)(2);
  VNStageIntLLRInputS2xD(217)(1) <= CNStageIntLLROutputS2xD(75)(3);
  VNStageIntLLRInputS2xD(288)(1) <= CNStageIntLLROutputS2xD(75)(4);
  VNStageIntLLRInputS2xD(348)(1) <= CNStageIntLLROutputS2xD(75)(5);
  VNStageIntLLRInputS2xD(20)(1) <= CNStageIntLLROutputS2xD(76)(0);
  VNStageIntLLRInputS2xD(99)(1) <= CNStageIntLLROutputS2xD(76)(1);
  VNStageIntLLRInputS2xD(152)(1) <= CNStageIntLLROutputS2xD(76)(2);
  VNStageIntLLRInputS2xD(223)(1) <= CNStageIntLLROutputS2xD(76)(3);
  VNStageIntLLRInputS2xD(283)(1) <= CNStageIntLLROutputS2xD(76)(4);
  VNStageIntLLRInputS2xD(358)(1) <= CNStageIntLLROutputS2xD(76)(5);
  VNStageIntLLRInputS2xD(19)(1) <= CNStageIntLLROutputS2xD(77)(0);
  VNStageIntLLRInputS2xD(87)(1) <= CNStageIntLLROutputS2xD(77)(1);
  VNStageIntLLRInputS2xD(158)(1) <= CNStageIntLLROutputS2xD(77)(2);
  VNStageIntLLRInputS2xD(218)(1) <= CNStageIntLLROutputS2xD(77)(3);
  VNStageIntLLRInputS2xD(293)(1) <= CNStageIntLLROutputS2xD(77)(4);
  VNStageIntLLRInputS2xD(380)(0) <= CNStageIntLLROutputS2xD(77)(5);
  VNStageIntLLRInputS2xD(18)(1) <= CNStageIntLLROutputS2xD(78)(0);
  VNStageIntLLRInputS2xD(93)(1) <= CNStageIntLLROutputS2xD(78)(1);
  VNStageIntLLRInputS2xD(153)(1) <= CNStageIntLLROutputS2xD(78)(2);
  VNStageIntLLRInputS2xD(228)(1) <= CNStageIntLLROutputS2xD(78)(3);
  VNStageIntLLRInputS2xD(315)(0) <= CNStageIntLLROutputS2xD(78)(4);
  VNStageIntLLRInputS2xD(335)(1) <= CNStageIntLLROutputS2xD(78)(5);
  VNStageIntLLRInputS2xD(17)(1) <= CNStageIntLLROutputS2xD(79)(0);
  VNStageIntLLRInputS2xD(88)(1) <= CNStageIntLLROutputS2xD(79)(1);
  VNStageIntLLRInputS2xD(163)(1) <= CNStageIntLLROutputS2xD(79)(2);
  VNStageIntLLRInputS2xD(250)(0) <= CNStageIntLLROutputS2xD(79)(3);
  VNStageIntLLRInputS2xD(270)(1) <= CNStageIntLLROutputS2xD(79)(4);
  VNStageIntLLRInputS2xD(383)(1) <= CNStageIntLLROutputS2xD(79)(5);
  VNStageIntLLRInputS2xD(15)(1) <= CNStageIntLLROutputS2xD(80)(0);
  VNStageIntLLRInputS2xD(120)(1) <= CNStageIntLLROutputS2xD(80)(1);
  VNStageIntLLRInputS2xD(140)(1) <= CNStageIntLLROutputS2xD(80)(2);
  VNStageIntLLRInputS2xD(253)(0) <= CNStageIntLLROutputS2xD(80)(3);
  VNStageIntLLRInputS2xD(305)(1) <= CNStageIntLLROutputS2xD(80)(4);
  VNStageIntLLRInputS2xD(338)(1) <= CNStageIntLLROutputS2xD(80)(5);
  VNStageIntLLRInputS2xD(14)(1) <= CNStageIntLLROutputS2xD(81)(0);
  VNStageIntLLRInputS2xD(75)(1) <= CNStageIntLLROutputS2xD(81)(1);
  VNStageIntLLRInputS2xD(188)(0) <= CNStageIntLLROutputS2xD(81)(2);
  VNStageIntLLRInputS2xD(240)(1) <= CNStageIntLLROutputS2xD(81)(3);
  VNStageIntLLRInputS2xD(273)(1) <= CNStageIntLLROutputS2xD(81)(4);
  VNStageIntLLRInputS2xD(350)(1) <= CNStageIntLLROutputS2xD(81)(5);
  VNStageIntLLRInputS2xD(13)(0) <= CNStageIntLLROutputS2xD(82)(0);
  VNStageIntLLRInputS2xD(123)(0) <= CNStageIntLLROutputS2xD(82)(1);
  VNStageIntLLRInputS2xD(175)(1) <= CNStageIntLLROutputS2xD(82)(2);
  VNStageIntLLRInputS2xD(208)(1) <= CNStageIntLLROutputS2xD(82)(3);
  VNStageIntLLRInputS2xD(285)(1) <= CNStageIntLLROutputS2xD(82)(4);
  VNStageIntLLRInputS2xD(364)(1) <= CNStageIntLLROutputS2xD(82)(5);
  VNStageIntLLRInputS2xD(12)(1) <= CNStageIntLLROutputS2xD(83)(0);
  VNStageIntLLRInputS2xD(110)(1) <= CNStageIntLLROutputS2xD(83)(1);
  VNStageIntLLRInputS2xD(143)(1) <= CNStageIntLLROutputS2xD(83)(2);
  VNStageIntLLRInputS2xD(220)(1) <= CNStageIntLLROutputS2xD(83)(3);
  VNStageIntLLRInputS2xD(299)(0) <= CNStageIntLLROutputS2xD(83)(4);
  VNStageIntLLRInputS2xD(345)(1) <= CNStageIntLLROutputS2xD(83)(5);
  VNStageIntLLRInputS2xD(11)(1) <= CNStageIntLLROutputS2xD(84)(0);
  VNStageIntLLRInputS2xD(78)(1) <= CNStageIntLLROutputS2xD(84)(1);
  VNStageIntLLRInputS2xD(155)(1) <= CNStageIntLLROutputS2xD(84)(2);
  VNStageIntLLRInputS2xD(234)(1) <= CNStageIntLLROutputS2xD(84)(3);
  VNStageIntLLRInputS2xD(280)(1) <= CNStageIntLLROutputS2xD(84)(4);
  VNStageIntLLRInputS2xD(322)(1) <= CNStageIntLLROutputS2xD(84)(5);
  VNStageIntLLRInputS2xD(10)(1) <= CNStageIntLLROutputS2xD(85)(0);
  VNStageIntLLRInputS2xD(90)(1) <= CNStageIntLLROutputS2xD(85)(1);
  VNStageIntLLRInputS2xD(169)(1) <= CNStageIntLLROutputS2xD(85)(2);
  VNStageIntLLRInputS2xD(215)(1) <= CNStageIntLLROutputS2xD(85)(3);
  VNStageIntLLRInputS2xD(257)(1) <= CNStageIntLLROutputS2xD(85)(4);
  VNStageIntLLRInputS2xD(374)(1) <= CNStageIntLLROutputS2xD(85)(5);
  VNStageIntLLRInputS2xD(9)(1) <= CNStageIntLLROutputS2xD(86)(0);
  VNStageIntLLRInputS2xD(104)(1) <= CNStageIntLLROutputS2xD(86)(1);
  VNStageIntLLRInputS2xD(150)(1) <= CNStageIntLLROutputS2xD(86)(2);
  VNStageIntLLRInputS2xD(255)(1) <= CNStageIntLLROutputS2xD(86)(3);
  VNStageIntLLRInputS2xD(309)(1) <= CNStageIntLLROutputS2xD(86)(4);
  VNStageIntLLRInputS2xD(378)(0) <= CNStageIntLLROutputS2xD(86)(5);
  VNStageIntLLRInputS2xD(7)(1) <= CNStageIntLLROutputS2xD(87)(0);
  VNStageIntLLRInputS2xD(125)(0) <= CNStageIntLLROutputS2xD(87)(1);
  VNStageIntLLRInputS2xD(179)(1) <= CNStageIntLLROutputS2xD(87)(2);
  VNStageIntLLRInputS2xD(248)(1) <= CNStageIntLLROutputS2xD(87)(3);
  VNStageIntLLRInputS2xD(306)(1) <= CNStageIntLLROutputS2xD(87)(4);
  VNStageIntLLRInputS2xD(382)(0) <= CNStageIntLLROutputS2xD(87)(5);
  VNStageIntLLRInputS2xD(6)(1) <= CNStageIntLLROutputS2xD(88)(0);
  VNStageIntLLRInputS2xD(114)(1) <= CNStageIntLLROutputS2xD(88)(1);
  VNStageIntLLRInputS2xD(183)(1) <= CNStageIntLLROutputS2xD(88)(2);
  VNStageIntLLRInputS2xD(241)(1) <= CNStageIntLLROutputS2xD(88)(3);
  VNStageIntLLRInputS2xD(317)(0) <= CNStageIntLLROutputS2xD(88)(4);
  VNStageIntLLRInputS2xD(354)(1) <= CNStageIntLLROutputS2xD(88)(5);
  VNStageIntLLRInputS2xD(5)(1) <= CNStageIntLLROutputS2xD(89)(0);
  VNStageIntLLRInputS2xD(118)(1) <= CNStageIntLLROutputS2xD(89)(1);
  VNStageIntLLRInputS2xD(176)(1) <= CNStageIntLLROutputS2xD(89)(2);
  VNStageIntLLRInputS2xD(252)(0) <= CNStageIntLLROutputS2xD(89)(3);
  VNStageIntLLRInputS2xD(289)(1) <= CNStageIntLLROutputS2xD(89)(4);
  VNStageIntLLRInputS2xD(346)(1) <= CNStageIntLLROutputS2xD(89)(5);
  VNStageIntLLRInputS2xD(4)(1) <= CNStageIntLLROutputS2xD(90)(0);
  VNStageIntLLRInputS2xD(111)(1) <= CNStageIntLLROutputS2xD(90)(1);
  VNStageIntLLRInputS2xD(187)(0) <= CNStageIntLLROutputS2xD(90)(2);
  VNStageIntLLRInputS2xD(224)(1) <= CNStageIntLLROutputS2xD(90)(3);
  VNStageIntLLRInputS2xD(281)(1) <= CNStageIntLLROutputS2xD(90)(4);
  VNStageIntLLRInputS2xD(363)(0) <= CNStageIntLLROutputS2xD(90)(5);
  VNStageIntLLRInputS2xD(3)(0) <= CNStageIntLLROutputS2xD(91)(0);
  VNStageIntLLRInputS2xD(122)(0) <= CNStageIntLLROutputS2xD(91)(1);
  VNStageIntLLRInputS2xD(159)(1) <= CNStageIntLLROutputS2xD(91)(2);
  VNStageIntLLRInputS2xD(216)(1) <= CNStageIntLLROutputS2xD(91)(3);
  VNStageIntLLRInputS2xD(298)(1) <= CNStageIntLLROutputS2xD(91)(4);
  VNStageIntLLRInputS2xD(360)(1) <= CNStageIntLLROutputS2xD(91)(5);
  VNStageIntLLRInputS2xD(2)(1) <= CNStageIntLLROutputS2xD(92)(0);
  VNStageIntLLRInputS2xD(94)(1) <= CNStageIntLLROutputS2xD(92)(1);
  VNStageIntLLRInputS2xD(151)(1) <= CNStageIntLLROutputS2xD(92)(2);
  VNStageIntLLRInputS2xD(233)(1) <= CNStageIntLLROutputS2xD(92)(3);
  VNStageIntLLRInputS2xD(295)(1) <= CNStageIntLLROutputS2xD(92)(4);
  VNStageIntLLRInputS2xD(331)(1) <= CNStageIntLLROutputS2xD(92)(5);
  VNStageIntLLRInputS2xD(63)(1) <= CNStageIntLLROutputS2xD(93)(0);
  VNStageIntLLRInputS2xD(103)(1) <= CNStageIntLLROutputS2xD(93)(1);
  VNStageIntLLRInputS2xD(165)(1) <= CNStageIntLLROutputS2xD(93)(2);
  VNStageIntLLRInputS2xD(201)(1) <= CNStageIntLLROutputS2xD(93)(3);
  VNStageIntLLRInputS2xD(286)(1) <= CNStageIntLLROutputS2xD(93)(4);
  VNStageIntLLRInputS2xD(337)(1) <= CNStageIntLLROutputS2xD(93)(5);
  VNStageIntLLRInputS2xD(62)(0) <= CNStageIntLLROutputS2xD(94)(0);
  VNStageIntLLRInputS2xD(100)(1) <= CNStageIntLLROutputS2xD(94)(1);
  VNStageIntLLRInputS2xD(136)(1) <= CNStageIntLLROutputS2xD(94)(2);
  VNStageIntLLRInputS2xD(221)(1) <= CNStageIntLLROutputS2xD(94)(3);
  VNStageIntLLRInputS2xD(272)(1) <= CNStageIntLLROutputS2xD(94)(4);
  VNStageIntLLRInputS2xD(327)(1) <= CNStageIntLLROutputS2xD(94)(5);
  VNStageIntLLRInputS2xD(61)(0) <= CNStageIntLLROutputS2xD(95)(0);
  VNStageIntLLRInputS2xD(71)(1) <= CNStageIntLLROutputS2xD(95)(1);
  VNStageIntLLRInputS2xD(156)(1) <= CNStageIntLLROutputS2xD(95)(2);
  VNStageIntLLRInputS2xD(207)(1) <= CNStageIntLLROutputS2xD(95)(3);
  VNStageIntLLRInputS2xD(262)(1) <= CNStageIntLLROutputS2xD(95)(4);
  VNStageIntLLRInputS2xD(356)(1) <= CNStageIntLLROutputS2xD(95)(5);
  VNStageIntLLRInputS2xD(60)(0) <= CNStageIntLLROutputS2xD(96)(0);
  VNStageIntLLRInputS2xD(91)(1) <= CNStageIntLLROutputS2xD(96)(1);
  VNStageIntLLRInputS2xD(142)(1) <= CNStageIntLLROutputS2xD(96)(2);
  VNStageIntLLRInputS2xD(197)(1) <= CNStageIntLLROutputS2xD(96)(3);
  VNStageIntLLRInputS2xD(291)(1) <= CNStageIntLLROutputS2xD(96)(4);
  VNStageIntLLRInputS2xD(339)(1) <= CNStageIntLLROutputS2xD(96)(5);
  VNStageIntLLRInputS2xD(58)(0) <= CNStageIntLLROutputS2xD(97)(0);
  VNStageIntLLRInputS2xD(67)(0) <= CNStageIntLLROutputS2xD(97)(1);
  VNStageIntLLRInputS2xD(161)(1) <= CNStageIntLLROutputS2xD(97)(2);
  VNStageIntLLRInputS2xD(209)(1) <= CNStageIntLLROutputS2xD(97)(3);
  VNStageIntLLRInputS2xD(304)(1) <= CNStageIntLLROutputS2xD(97)(4);
  VNStageIntLLRInputS2xD(329)(1) <= CNStageIntLLROutputS2xD(97)(5);
  VNStageIntLLRInputS2xD(57)(0) <= CNStageIntLLROutputS2xD(98)(0);
  VNStageIntLLRInputS2xD(96)(1) <= CNStageIntLLROutputS2xD(98)(1);
  VNStageIntLLRInputS2xD(144)(1) <= CNStageIntLLROutputS2xD(98)(2);
  VNStageIntLLRInputS2xD(239)(1) <= CNStageIntLLROutputS2xD(98)(3);
  VNStageIntLLRInputS2xD(264)(1) <= CNStageIntLLROutputS2xD(98)(4);
  VNStageIntLLRInputS2xD(365)(1) <= CNStageIntLLROutputS2xD(98)(5);
  VNStageIntLLRInputS2xD(56)(1) <= CNStageIntLLROutputS2xD(99)(0);
  VNStageIntLLRInputS2xD(79)(1) <= CNStageIntLLROutputS2xD(99)(1);
  VNStageIntLLRInputS2xD(174)(1) <= CNStageIntLLROutputS2xD(99)(2);
  VNStageIntLLRInputS2xD(199)(1) <= CNStageIntLLROutputS2xD(99)(3);
  VNStageIntLLRInputS2xD(300)(1) <= CNStageIntLLROutputS2xD(99)(4);
  VNStageIntLLRInputS2xD(349)(1) <= CNStageIntLLROutputS2xD(99)(5);
  VNStageIntLLRInputS2xD(55)(1) <= CNStageIntLLROutputS2xD(100)(0);
  VNStageIntLLRInputS2xD(109)(1) <= CNStageIntLLROutputS2xD(100)(1);
  VNStageIntLLRInputS2xD(134)(1) <= CNStageIntLLROutputS2xD(100)(2);
  VNStageIntLLRInputS2xD(235)(0) <= CNStageIntLLROutputS2xD(100)(3);
  VNStageIntLLRInputS2xD(284)(1) <= CNStageIntLLROutputS2xD(100)(4);
  VNStageIntLLRInputS2xD(352)(1) <= CNStageIntLLROutputS2xD(100)(5);
  VNStageIntLLRInputS2xD(54)(1) <= CNStageIntLLROutputS2xD(101)(0);
  VNStageIntLLRInputS2xD(69)(1) <= CNStageIntLLROutputS2xD(101)(1);
  VNStageIntLLRInputS2xD(170)(1) <= CNStageIntLLROutputS2xD(101)(2);
  VNStageIntLLRInputS2xD(219)(1) <= CNStageIntLLROutputS2xD(101)(3);
  VNStageIntLLRInputS2xD(287)(1) <= CNStageIntLLROutputS2xD(101)(4);
  VNStageIntLLRInputS2xD(330)(1) <= CNStageIntLLROutputS2xD(101)(5);
  VNStageIntLLRInputS2xD(52)(0) <= CNStageIntLLROutputS2xD(102)(0);
  VNStageIntLLRInputS2xD(89)(1) <= CNStageIntLLROutputS2xD(102)(1);
  VNStageIntLLRInputS2xD(157)(1) <= CNStageIntLLROutputS2xD(102)(2);
  VNStageIntLLRInputS2xD(200)(1) <= CNStageIntLLROutputS2xD(102)(3);
  VNStageIntLLRInputS2xD(303)(1) <= CNStageIntLLROutputS2xD(102)(4);
  VNStageIntLLRInputS2xD(366)(1) <= CNStageIntLLROutputS2xD(102)(5);
  VNStageIntLLRInputS2xD(51)(1) <= CNStageIntLLROutputS2xD(103)(0);
  VNStageIntLLRInputS2xD(92)(1) <= CNStageIntLLROutputS2xD(103)(1);
  VNStageIntLLRInputS2xD(135)(1) <= CNStageIntLLROutputS2xD(103)(2);
  VNStageIntLLRInputS2xD(238)(1) <= CNStageIntLLROutputS2xD(103)(3);
  VNStageIntLLRInputS2xD(301)(1) <= CNStageIntLLROutputS2xD(103)(4);
  VNStageIntLLRInputS2xD(328)(1) <= CNStageIntLLROutputS2xD(103)(5);
  VNStageIntLLRInputS2xD(50)(1) <= CNStageIntLLROutputS2xD(104)(0);
  VNStageIntLLRInputS2xD(70)(1) <= CNStageIntLLROutputS2xD(104)(1);
  VNStageIntLLRInputS2xD(173)(1) <= CNStageIntLLROutputS2xD(104)(2);
  VNStageIntLLRInputS2xD(236)(1) <= CNStageIntLLROutputS2xD(104)(3);
  VNStageIntLLRInputS2xD(263)(1) <= CNStageIntLLROutputS2xD(104)(4);
  VNStageIntLLRInputS2xD(336)(1) <= CNStageIntLLROutputS2xD(104)(5);
  VNStageIntLLRInputS2xD(49)(1) <= CNStageIntLLROutputS2xD(105)(0);
  VNStageIntLLRInputS2xD(108)(1) <= CNStageIntLLROutputS2xD(105)(1);
  VNStageIntLLRInputS2xD(171)(0) <= CNStageIntLLROutputS2xD(105)(2);
  VNStageIntLLRInputS2xD(198)(1) <= CNStageIntLLROutputS2xD(105)(3);
  VNStageIntLLRInputS2xD(271)(1) <= CNStageIntLLROutputS2xD(105)(4);
  VNStageIntLLRInputS2xD(379)(0) <= CNStageIntLLROutputS2xD(105)(5);
  VNStageIntLLRInputS2xD(46)(1) <= CNStageIntLLROutputS2xD(106)(0);
  VNStageIntLLRInputS2xD(76)(1) <= CNStageIntLLROutputS2xD(106)(1);
  VNStageIntLLRInputS2xD(184)(1) <= CNStageIntLLROutputS2xD(106)(2);
  VNStageIntLLRInputS2xD(243)(1) <= CNStageIntLLROutputS2xD(106)(3);
  VNStageIntLLRInputS2xD(256)(1) <= CNStageIntLLROutputS2xD(106)(4);
  VNStageIntLLRInputS2xD(372)(0) <= CNStageIntLLROutputS2xD(106)(5);
  VNStageIntLLRInputS2xD(45)(1) <= CNStageIntLLROutputS2xD(107)(0);
  VNStageIntLLRInputS2xD(119)(1) <= CNStageIntLLROutputS2xD(107)(1);
  VNStageIntLLRInputS2xD(178)(1) <= CNStageIntLLROutputS2xD(107)(2);
  VNStageIntLLRInputS2xD(192)(1) <= CNStageIntLLROutputS2xD(107)(3);
  VNStageIntLLRInputS2xD(307)(1) <= CNStageIntLLROutputS2xD(107)(4);
  VNStageIntLLRInputS2xD(377)(0) <= CNStageIntLLROutputS2xD(107)(5);
  VNStageIntLLRInputS2xD(44)(1) <= CNStageIntLLROutputS2xD(108)(0);
  VNStageIntLLRInputS2xD(113)(1) <= CNStageIntLLROutputS2xD(108)(1);
  VNStageIntLLRInputS2xD(128)(1) <= CNStageIntLLROutputS2xD(108)(2);
  VNStageIntLLRInputS2xD(242)(1) <= CNStageIntLLROutputS2xD(108)(3);
  VNStageIntLLRInputS2xD(312)(1) <= CNStageIntLLROutputS2xD(108)(4);
  VNStageIntLLRInputS2xD(333)(0) <= CNStageIntLLROutputS2xD(108)(5);
  VNStageIntLLRInputS2xD(43)(0) <= CNStageIntLLROutputS2xD(109)(0);
  VNStageIntLLRInputS2xD(64)(1) <= CNStageIntLLROutputS2xD(109)(1);
  VNStageIntLLRInputS2xD(177)(1) <= CNStageIntLLROutputS2xD(109)(2);
  VNStageIntLLRInputS2xD(247)(1) <= CNStageIntLLROutputS2xD(109)(3);
  VNStageIntLLRInputS2xD(268)(1) <= CNStageIntLLROutputS2xD(109)(4);
  VNStageIntLLRInputS2xD(324)(1) <= CNStageIntLLROutputS2xD(109)(5);
  VNStageIntLLRInputS2xD(0)(1) <= CNStageIntLLROutputS2xD(110)(0);
  VNStageIntLLRInputS2xD(107)(0) <= CNStageIntLLROutputS2xD(110)(1);
  VNStageIntLLRInputS2xD(172)(1) <= CNStageIntLLROutputS2xD(110)(2);
  VNStageIntLLRInputS2xD(237)(1) <= CNStageIntLLROutputS2xD(110)(3);
  VNStageIntLLRInputS2xD(302)(1) <= CNStageIntLLROutputS2xD(110)(4);
  VNStageIntLLRInputS2xD(367)(1) <= CNStageIntLLROutputS2xD(110)(5);
  VNStageIntLLRInputS2xD(32)(2) <= CNStageIntLLROutputS2xD(111)(0);
  VNStageIntLLRInputS2xD(117)(2) <= CNStageIntLLROutputS2xD(111)(1);
  VNStageIntLLRInputS2xD(136)(2) <= CNStageIntLLROutputS2xD(111)(2);
  VNStageIntLLRInputS2xD(198)(2) <= CNStageIntLLROutputS2xD(111)(3);
  VNStageIntLLRInputS2xD(297)(2) <= CNStageIntLLROutputS2xD(111)(4);
  VNStageIntLLRInputS2xD(382)(1) <= CNStageIntLLROutputS2xD(111)(5);
  VNStageIntLLRInputS2xD(30)(2) <= CNStageIntLLROutputS2xD(112)(0);
  VNStageIntLLRInputS2xD(68)(1) <= CNStageIntLLROutputS2xD(112)(1);
  VNStageIntLLRInputS2xD(167)(2) <= CNStageIntLLROutputS2xD(112)(2);
  VNStageIntLLRInputS2xD(252)(1) <= CNStageIntLLROutputS2xD(112)(3);
  VNStageIntLLRInputS2xD(303)(2) <= CNStageIntLLROutputS2xD(112)(4);
  VNStageIntLLRInputS2xD(358)(2) <= CNStageIntLLROutputS2xD(112)(5);
  VNStageIntLLRInputS2xD(29)(2) <= CNStageIntLLROutputS2xD(113)(0);
  VNStageIntLLRInputS2xD(102)(2) <= CNStageIntLLROutputS2xD(113)(1);
  VNStageIntLLRInputS2xD(187)(1) <= CNStageIntLLROutputS2xD(113)(2);
  VNStageIntLLRInputS2xD(238)(2) <= CNStageIntLLROutputS2xD(113)(3);
  VNStageIntLLRInputS2xD(293)(2) <= CNStageIntLLROutputS2xD(113)(4);
  VNStageIntLLRInputS2xD(324)(2) <= CNStageIntLLROutputS2xD(113)(5);
  VNStageIntLLRInputS2xD(28)(2) <= CNStageIntLLROutputS2xD(114)(0);
  VNStageIntLLRInputS2xD(122)(1) <= CNStageIntLLROutputS2xD(114)(1);
  VNStageIntLLRInputS2xD(173)(2) <= CNStageIntLLROutputS2xD(114)(2);
  VNStageIntLLRInputS2xD(228)(2) <= CNStageIntLLROutputS2xD(114)(3);
  VNStageIntLLRInputS2xD(259)(1) <= CNStageIntLLROutputS2xD(114)(4);
  VNStageIntLLRInputS2xD(370)(1) <= CNStageIntLLROutputS2xD(114)(5);
  VNStageIntLLRInputS2xD(27)(2) <= CNStageIntLLROutputS2xD(115)(0);
  VNStageIntLLRInputS2xD(108)(2) <= CNStageIntLLROutputS2xD(115)(1);
  VNStageIntLLRInputS2xD(163)(2) <= CNStageIntLLROutputS2xD(115)(2);
  VNStageIntLLRInputS2xD(194)(2) <= CNStageIntLLROutputS2xD(115)(3);
  VNStageIntLLRInputS2xD(305)(2) <= CNStageIntLLROutputS2xD(115)(4);
  VNStageIntLLRInputS2xD(337)(2) <= CNStageIntLLROutputS2xD(115)(5);
  VNStageIntLLRInputS2xD(26)(2) <= CNStageIntLLROutputS2xD(116)(0);
  VNStageIntLLRInputS2xD(98)(1) <= CNStageIntLLROutputS2xD(116)(1);
  VNStageIntLLRInputS2xD(129)(2) <= CNStageIntLLROutputS2xD(116)(2);
  VNStageIntLLRInputS2xD(240)(2) <= CNStageIntLLROutputS2xD(116)(3);
  VNStageIntLLRInputS2xD(272)(2) <= CNStageIntLLROutputS2xD(116)(4);
  VNStageIntLLRInputS2xD(360)(2) <= CNStageIntLLROutputS2xD(116)(5);
  VNStageIntLLRInputS2xD(25)(2) <= CNStageIntLLROutputS2xD(117)(0);
  VNStageIntLLRInputS2xD(127)(2) <= CNStageIntLLROutputS2xD(117)(1);
  VNStageIntLLRInputS2xD(175)(2) <= CNStageIntLLROutputS2xD(117)(2);
  VNStageIntLLRInputS2xD(207)(2) <= CNStageIntLLROutputS2xD(117)(3);
  VNStageIntLLRInputS2xD(295)(2) <= CNStageIntLLROutputS2xD(117)(4);
  VNStageIntLLRInputS2xD(333)(1) <= CNStageIntLLROutputS2xD(117)(5);
  VNStageIntLLRInputS2xD(24)(2) <= CNStageIntLLROutputS2xD(118)(0);
  VNStageIntLLRInputS2xD(110)(2) <= CNStageIntLLROutputS2xD(118)(1);
  VNStageIntLLRInputS2xD(142)(2) <= CNStageIntLLROutputS2xD(118)(2);
  VNStageIntLLRInputS2xD(230)(1) <= CNStageIntLLROutputS2xD(118)(3);
  VNStageIntLLRInputS2xD(268)(2) <= CNStageIntLLROutputS2xD(118)(4);
  VNStageIntLLRInputS2xD(380)(1) <= CNStageIntLLROutputS2xD(118)(5);
  VNStageIntLLRInputS2xD(23)(2) <= CNStageIntLLROutputS2xD(119)(0);
  VNStageIntLLRInputS2xD(77)(0) <= CNStageIntLLROutputS2xD(119)(1);
  VNStageIntLLRInputS2xD(165)(2) <= CNStageIntLLROutputS2xD(119)(2);
  VNStageIntLLRInputS2xD(203)(2) <= CNStageIntLLROutputS2xD(119)(3);
  VNStageIntLLRInputS2xD(315)(1) <= CNStageIntLLROutputS2xD(119)(4);
  VNStageIntLLRInputS2xD(383)(2) <= CNStageIntLLROutputS2xD(119)(5);
  VNStageIntLLRInputS2xD(22)(2) <= CNStageIntLLROutputS2xD(120)(0);
  VNStageIntLLRInputS2xD(100)(2) <= CNStageIntLLROutputS2xD(120)(1);
  VNStageIntLLRInputS2xD(138)(2) <= CNStageIntLLROutputS2xD(120)(2);
  VNStageIntLLRInputS2xD(250)(1) <= CNStageIntLLROutputS2xD(120)(3);
  VNStageIntLLRInputS2xD(318)(0) <= CNStageIntLLROutputS2xD(120)(4);
  VNStageIntLLRInputS2xD(361)(2) <= CNStageIntLLROutputS2xD(120)(5);
  VNStageIntLLRInputS2xD(21)(2) <= CNStageIntLLROutputS2xD(121)(0);
  VNStageIntLLRInputS2xD(73)(2) <= CNStageIntLLROutputS2xD(121)(1);
  VNStageIntLLRInputS2xD(185)(0) <= CNStageIntLLROutputS2xD(121)(2);
  VNStageIntLLRInputS2xD(253)(1) <= CNStageIntLLROutputS2xD(121)(3);
  VNStageIntLLRInputS2xD(296)(2) <= CNStageIntLLROutputS2xD(121)(4);
  VNStageIntLLRInputS2xD(336)(2) <= CNStageIntLLROutputS2xD(121)(5);
  VNStageIntLLRInputS2xD(19)(2) <= CNStageIntLLROutputS2xD(122)(0);
  VNStageIntLLRInputS2xD(123)(1) <= CNStageIntLLROutputS2xD(122)(1);
  VNStageIntLLRInputS2xD(166)(2) <= CNStageIntLLROutputS2xD(122)(2);
  VNStageIntLLRInputS2xD(206)(1) <= CNStageIntLLROutputS2xD(122)(3);
  VNStageIntLLRInputS2xD(269)(1) <= CNStageIntLLROutputS2xD(122)(4);
  VNStageIntLLRInputS2xD(359)(2) <= CNStageIntLLROutputS2xD(122)(5);
  VNStageIntLLRInputS2xD(18)(2) <= CNStageIntLLROutputS2xD(123)(0);
  VNStageIntLLRInputS2xD(101)(2) <= CNStageIntLLROutputS2xD(123)(1);
  VNStageIntLLRInputS2xD(141)(0) <= CNStageIntLLROutputS2xD(123)(2);
  VNStageIntLLRInputS2xD(204)(2) <= CNStageIntLLROutputS2xD(123)(3);
  VNStageIntLLRInputS2xD(294)(2) <= CNStageIntLLROutputS2xD(123)(4);
  VNStageIntLLRInputS2xD(367)(2) <= CNStageIntLLROutputS2xD(123)(5);
  VNStageIntLLRInputS2xD(17)(2) <= CNStageIntLLROutputS2xD(124)(0);
  VNStageIntLLRInputS2xD(76)(2) <= CNStageIntLLROutputS2xD(124)(1);
  VNStageIntLLRInputS2xD(139)(2) <= CNStageIntLLROutputS2xD(124)(2);
  VNStageIntLLRInputS2xD(229)(2) <= CNStageIntLLROutputS2xD(124)(3);
  VNStageIntLLRInputS2xD(302)(2) <= CNStageIntLLROutputS2xD(124)(4);
  VNStageIntLLRInputS2xD(347)(2) <= CNStageIntLLROutputS2xD(124)(5);
  VNStageIntLLRInputS2xD(16)(1) <= CNStageIntLLROutputS2xD(125)(0);
  VNStageIntLLRInputS2xD(74)(2) <= CNStageIntLLROutputS2xD(125)(1);
  VNStageIntLLRInputS2xD(164)(2) <= CNStageIntLLROutputS2xD(125)(2);
  VNStageIntLLRInputS2xD(237)(2) <= CNStageIntLLROutputS2xD(125)(3);
  VNStageIntLLRInputS2xD(282)(2) <= CNStageIntLLROutputS2xD(125)(4);
  VNStageIntLLRInputS2xD(341)(2) <= CNStageIntLLROutputS2xD(125)(5);
  VNStageIntLLRInputS2xD(15)(2) <= CNStageIntLLROutputS2xD(126)(0);
  VNStageIntLLRInputS2xD(99)(2) <= CNStageIntLLROutputS2xD(126)(1);
  VNStageIntLLRInputS2xD(172)(2) <= CNStageIntLLROutputS2xD(126)(2);
  VNStageIntLLRInputS2xD(217)(2) <= CNStageIntLLROutputS2xD(126)(3);
  VNStageIntLLRInputS2xD(276)(2) <= CNStageIntLLROutputS2xD(126)(4);
  VNStageIntLLRInputS2xD(320)(1) <= CNStageIntLLROutputS2xD(126)(5);
  VNStageIntLLRInputS2xD(14)(2) <= CNStageIntLLROutputS2xD(127)(0);
  VNStageIntLLRInputS2xD(107)(1) <= CNStageIntLLROutputS2xD(127)(1);
  VNStageIntLLRInputS2xD(152)(2) <= CNStageIntLLROutputS2xD(127)(2);
  VNStageIntLLRInputS2xD(211)(2) <= CNStageIntLLROutputS2xD(127)(3);
  VNStageIntLLRInputS2xD(256)(2) <= CNStageIntLLROutputS2xD(127)(4);
  VNStageIntLLRInputS2xD(340)(2) <= CNStageIntLLROutputS2xD(127)(5);
  VNStageIntLLRInputS2xD(13)(1) <= CNStageIntLLROutputS2xD(128)(0);
  VNStageIntLLRInputS2xD(87)(2) <= CNStageIntLLROutputS2xD(128)(1);
  VNStageIntLLRInputS2xD(146)(2) <= CNStageIntLLROutputS2xD(128)(2);
  VNStageIntLLRInputS2xD(192)(2) <= CNStageIntLLROutputS2xD(128)(3);
  VNStageIntLLRInputS2xD(275)(2) <= CNStageIntLLROutputS2xD(128)(4);
  VNStageIntLLRInputS2xD(345)(2) <= CNStageIntLLROutputS2xD(128)(5);
  VNStageIntLLRInputS2xD(12)(2) <= CNStageIntLLROutputS2xD(129)(0);
  VNStageIntLLRInputS2xD(81)(2) <= CNStageIntLLROutputS2xD(129)(1);
  VNStageIntLLRInputS2xD(128)(2) <= CNStageIntLLROutputS2xD(129)(2);
  VNStageIntLLRInputS2xD(210)(2) <= CNStageIntLLROutputS2xD(129)(3);
  VNStageIntLLRInputS2xD(280)(2) <= CNStageIntLLROutputS2xD(129)(4);
  VNStageIntLLRInputS2xD(364)(2) <= CNStageIntLLROutputS2xD(129)(5);
  VNStageIntLLRInputS2xD(11)(2) <= CNStageIntLLROutputS2xD(130)(0);
  VNStageIntLLRInputS2xD(64)(2) <= CNStageIntLLROutputS2xD(130)(1);
  VNStageIntLLRInputS2xD(145)(2) <= CNStageIntLLROutputS2xD(130)(2);
  VNStageIntLLRInputS2xD(215)(2) <= CNStageIntLLROutputS2xD(130)(3);
  VNStageIntLLRInputS2xD(299)(1) <= CNStageIntLLROutputS2xD(130)(4);
  VNStageIntLLRInputS2xD(355)(2) <= CNStageIntLLROutputS2xD(130)(5);
  VNStageIntLLRInputS2xD(10)(2) <= CNStageIntLLROutputS2xD(131)(0);
  VNStageIntLLRInputS2xD(80)(2) <= CNStageIntLLROutputS2xD(131)(1);
  VNStageIntLLRInputS2xD(150)(2) <= CNStageIntLLROutputS2xD(131)(2);
  VNStageIntLLRInputS2xD(234)(2) <= CNStageIntLLROutputS2xD(131)(3);
  VNStageIntLLRInputS2xD(290)(2) <= CNStageIntLLROutputS2xD(131)(4);
  VNStageIntLLRInputS2xD(329)(2) <= CNStageIntLLROutputS2xD(131)(5);
  VNStageIntLLRInputS2xD(9)(2) <= CNStageIntLLROutputS2xD(132)(0);
  VNStageIntLLRInputS2xD(85)(1) <= CNStageIntLLROutputS2xD(132)(1);
  VNStageIntLLRInputS2xD(169)(2) <= CNStageIntLLROutputS2xD(132)(2);
  VNStageIntLLRInputS2xD(225)(2) <= CNStageIntLLROutputS2xD(132)(3);
  VNStageIntLLRInputS2xD(264)(2) <= CNStageIntLLROutputS2xD(132)(4);
  VNStageIntLLRInputS2xD(330)(2) <= CNStageIntLLROutputS2xD(132)(5);
  VNStageIntLLRInputS2xD(8)(1) <= CNStageIntLLROutputS2xD(133)(0);
  VNStageIntLLRInputS2xD(104)(2) <= CNStageIntLLROutputS2xD(133)(1);
  VNStageIntLLRInputS2xD(160)(2) <= CNStageIntLLROutputS2xD(133)(2);
  VNStageIntLLRInputS2xD(199)(2) <= CNStageIntLLROutputS2xD(133)(3);
  VNStageIntLLRInputS2xD(265)(1) <= CNStageIntLLROutputS2xD(133)(4);
  VNStageIntLLRInputS2xD(354)(2) <= CNStageIntLLROutputS2xD(133)(5);
  VNStageIntLLRInputS2xD(7)(2) <= CNStageIntLLROutputS2xD(134)(0);
  VNStageIntLLRInputS2xD(95)(2) <= CNStageIntLLROutputS2xD(134)(1);
  VNStageIntLLRInputS2xD(134)(2) <= CNStageIntLLROutputS2xD(134)(2);
  VNStageIntLLRInputS2xD(200)(2) <= CNStageIntLLROutputS2xD(134)(3);
  VNStageIntLLRInputS2xD(289)(2) <= CNStageIntLLROutputS2xD(134)(4);
  VNStageIntLLRInputS2xD(375)(2) <= CNStageIntLLROutputS2xD(134)(5);
  VNStageIntLLRInputS2xD(6)(2) <= CNStageIntLLROutputS2xD(135)(0);
  VNStageIntLLRInputS2xD(69)(2) <= CNStageIntLLROutputS2xD(135)(1);
  VNStageIntLLRInputS2xD(135)(2) <= CNStageIntLLROutputS2xD(135)(2);
  VNStageIntLLRInputS2xD(224)(2) <= CNStageIntLLROutputS2xD(135)(3);
  VNStageIntLLRInputS2xD(310)(2) <= CNStageIntLLROutputS2xD(135)(4);
  VNStageIntLLRInputS2xD(371)(1) <= CNStageIntLLROutputS2xD(135)(5);
  VNStageIntLLRInputS2xD(5)(2) <= CNStageIntLLROutputS2xD(136)(0);
  VNStageIntLLRInputS2xD(70)(2) <= CNStageIntLLROutputS2xD(136)(1);
  VNStageIntLLRInputS2xD(159)(2) <= CNStageIntLLROutputS2xD(136)(2);
  VNStageIntLLRInputS2xD(245)(2) <= CNStageIntLLROutputS2xD(136)(3);
  VNStageIntLLRInputS2xD(306)(2) <= CNStageIntLLROutputS2xD(136)(4);
  VNStageIntLLRInputS2xD(323)(1) <= CNStageIntLLROutputS2xD(136)(5);
  VNStageIntLLRInputS2xD(3)(1) <= CNStageIntLLROutputS2xD(137)(0);
  VNStageIntLLRInputS2xD(115)(2) <= CNStageIntLLROutputS2xD(137)(1);
  VNStageIntLLRInputS2xD(176)(2) <= CNStageIntLLROutputS2xD(137)(2);
  VNStageIntLLRInputS2xD(193)(2) <= CNStageIntLLROutputS2xD(137)(3);
  VNStageIntLLRInputS2xD(284)(2) <= CNStageIntLLROutputS2xD(137)(4);
  VNStageIntLLRInputS2xD(325)(2) <= CNStageIntLLROutputS2xD(137)(5);
  VNStageIntLLRInputS2xD(2)(2) <= CNStageIntLLROutputS2xD(138)(0);
  VNStageIntLLRInputS2xD(111)(2) <= CNStageIntLLROutputS2xD(138)(1);
  VNStageIntLLRInputS2xD(191)(2) <= CNStageIntLLROutputS2xD(138)(2);
  VNStageIntLLRInputS2xD(219)(2) <= CNStageIntLLROutputS2xD(138)(3);
  VNStageIntLLRInputS2xD(260)(2) <= CNStageIntLLROutputS2xD(138)(4);
  VNStageIntLLRInputS2xD(357)(2) <= CNStageIntLLROutputS2xD(138)(5);
  VNStageIntLLRInputS2xD(1)(1) <= CNStageIntLLROutputS2xD(139)(0);
  VNStageIntLLRInputS2xD(126)(1) <= CNStageIntLLROutputS2xD(139)(1);
  VNStageIntLLRInputS2xD(154)(1) <= CNStageIntLLROutputS2xD(139)(2);
  VNStageIntLLRInputS2xD(195)(1) <= CNStageIntLLROutputS2xD(139)(3);
  VNStageIntLLRInputS2xD(292)(2) <= CNStageIntLLROutputS2xD(139)(4);
  VNStageIntLLRInputS2xD(373)(1) <= CNStageIntLLROutputS2xD(139)(5);
  VNStageIntLLRInputS2xD(63)(2) <= CNStageIntLLROutputS2xD(140)(0);
  VNStageIntLLRInputS2xD(89)(2) <= CNStageIntLLROutputS2xD(140)(1);
  VNStageIntLLRInputS2xD(130)(2) <= CNStageIntLLROutputS2xD(140)(2);
  VNStageIntLLRInputS2xD(227)(2) <= CNStageIntLLROutputS2xD(140)(3);
  VNStageIntLLRInputS2xD(308)(0) <= CNStageIntLLROutputS2xD(140)(4);
  VNStageIntLLRInputS2xD(343)(2) <= CNStageIntLLROutputS2xD(140)(5);
  VNStageIntLLRInputS2xD(62)(1) <= CNStageIntLLROutputS2xD(141)(0);
  VNStageIntLLRInputS2xD(65)(2) <= CNStageIntLLROutputS2xD(141)(1);
  VNStageIntLLRInputS2xD(162)(2) <= CNStageIntLLROutputS2xD(141)(2);
  VNStageIntLLRInputS2xD(243)(2) <= CNStageIntLLROutputS2xD(141)(3);
  VNStageIntLLRInputS2xD(278)(2) <= CNStageIntLLROutputS2xD(141)(4);
  VNStageIntLLRInputS2xD(352)(2) <= CNStageIntLLROutputS2xD(141)(5);
  VNStageIntLLRInputS2xD(61)(1) <= CNStageIntLLROutputS2xD(142)(0);
  VNStageIntLLRInputS2xD(97)(2) <= CNStageIntLLROutputS2xD(142)(1);
  VNStageIntLLRInputS2xD(178)(2) <= CNStageIntLLROutputS2xD(142)(2);
  VNStageIntLLRInputS2xD(213)(2) <= CNStageIntLLROutputS2xD(142)(3);
  VNStageIntLLRInputS2xD(287)(2) <= CNStageIntLLROutputS2xD(142)(4);
  VNStageIntLLRInputS2xD(365)(2) <= CNStageIntLLROutputS2xD(142)(5);
  VNStageIntLLRInputS2xD(60)(1) <= CNStageIntLLROutputS2xD(143)(0);
  VNStageIntLLRInputS2xD(113)(2) <= CNStageIntLLROutputS2xD(143)(1);
  VNStageIntLLRInputS2xD(148)(2) <= CNStageIntLLROutputS2xD(143)(2);
  VNStageIntLLRInputS2xD(222)(1) <= CNStageIntLLROutputS2xD(143)(3);
  VNStageIntLLRInputS2xD(300)(2) <= CNStageIntLLROutputS2xD(143)(4);
  VNStageIntLLRInputS2xD(344)(2) <= CNStageIntLLROutputS2xD(143)(5);
  VNStageIntLLRInputS2xD(59)(0) <= CNStageIntLLROutputS2xD(144)(0);
  VNStageIntLLRInputS2xD(83)(2) <= CNStageIntLLROutputS2xD(144)(1);
  VNStageIntLLRInputS2xD(157)(2) <= CNStageIntLLROutputS2xD(144)(2);
  VNStageIntLLRInputS2xD(235)(1) <= CNStageIntLLROutputS2xD(144)(3);
  VNStageIntLLRInputS2xD(279)(2) <= CNStageIntLLROutputS2xD(144)(4);
  VNStageIntLLRInputS2xD(372)(1) <= CNStageIntLLROutputS2xD(144)(5);
  VNStageIntLLRInputS2xD(58)(1) <= CNStageIntLLROutputS2xD(145)(0);
  VNStageIntLLRInputS2xD(92)(2) <= CNStageIntLLROutputS2xD(145)(1);
  VNStageIntLLRInputS2xD(170)(2) <= CNStageIntLLROutputS2xD(145)(2);
  VNStageIntLLRInputS2xD(214)(2) <= CNStageIntLLROutputS2xD(145)(3);
  VNStageIntLLRInputS2xD(307)(2) <= CNStageIntLLROutputS2xD(145)(4);
  VNStageIntLLRInputS2xD(374)(2) <= CNStageIntLLROutputS2xD(145)(5);
  VNStageIntLLRInputS2xD(57)(1) <= CNStageIntLLROutputS2xD(146)(0);
  VNStageIntLLRInputS2xD(105)(1) <= CNStageIntLLROutputS2xD(146)(1);
  VNStageIntLLRInputS2xD(149)(2) <= CNStageIntLLROutputS2xD(146)(2);
  VNStageIntLLRInputS2xD(242)(2) <= CNStageIntLLROutputS2xD(146)(3);
  VNStageIntLLRInputS2xD(309)(2) <= CNStageIntLLROutputS2xD(146)(4);
  VNStageIntLLRInputS2xD(356)(2) <= CNStageIntLLROutputS2xD(146)(5);
  VNStageIntLLRInputS2xD(56)(2) <= CNStageIntLLROutputS2xD(147)(0);
  VNStageIntLLRInputS2xD(84)(2) <= CNStageIntLLROutputS2xD(147)(1);
  VNStageIntLLRInputS2xD(177)(2) <= CNStageIntLLROutputS2xD(147)(2);
  VNStageIntLLRInputS2xD(244)(0) <= CNStageIntLLROutputS2xD(147)(3);
  VNStageIntLLRInputS2xD(291)(2) <= CNStageIntLLROutputS2xD(147)(4);
  VNStageIntLLRInputS2xD(363)(1) <= CNStageIntLLROutputS2xD(147)(5);
  VNStageIntLLRInputS2xD(55)(2) <= CNStageIntLLROutputS2xD(148)(0);
  VNStageIntLLRInputS2xD(112)(2) <= CNStageIntLLROutputS2xD(148)(1);
  VNStageIntLLRInputS2xD(179)(2) <= CNStageIntLLROutputS2xD(148)(2);
  VNStageIntLLRInputS2xD(226)(1) <= CNStageIntLLROutputS2xD(148)(3);
  VNStageIntLLRInputS2xD(298)(2) <= CNStageIntLLROutputS2xD(148)(4);
  VNStageIntLLRInputS2xD(327)(2) <= CNStageIntLLROutputS2xD(148)(5);
  VNStageIntLLRInputS2xD(54)(2) <= CNStageIntLLROutputS2xD(149)(0);
  VNStageIntLLRInputS2xD(114)(2) <= CNStageIntLLROutputS2xD(149)(1);
  VNStageIntLLRInputS2xD(161)(2) <= CNStageIntLLROutputS2xD(149)(2);
  VNStageIntLLRInputS2xD(233)(2) <= CNStageIntLLROutputS2xD(149)(3);
  VNStageIntLLRInputS2xD(262)(2) <= CNStageIntLLROutputS2xD(149)(4);
  VNStageIntLLRInputS2xD(378)(1) <= CNStageIntLLROutputS2xD(149)(5);
  VNStageIntLLRInputS2xD(53)(1) <= CNStageIntLLROutputS2xD(150)(0);
  VNStageIntLLRInputS2xD(96)(2) <= CNStageIntLLROutputS2xD(150)(1);
  VNStageIntLLRInputS2xD(168)(1) <= CNStageIntLLROutputS2xD(150)(2);
  VNStageIntLLRInputS2xD(197)(2) <= CNStageIntLLROutputS2xD(150)(3);
  VNStageIntLLRInputS2xD(313)(0) <= CNStageIntLLROutputS2xD(150)(4);
  VNStageIntLLRInputS2xD(321)(2) <= CNStageIntLLROutputS2xD(150)(5);
  VNStageIntLLRInputS2xD(52)(1) <= CNStageIntLLROutputS2xD(151)(0);
  VNStageIntLLRInputS2xD(103)(2) <= CNStageIntLLROutputS2xD(151)(1);
  VNStageIntLLRInputS2xD(132)(1) <= CNStageIntLLROutputS2xD(151)(2);
  VNStageIntLLRInputS2xD(248)(2) <= CNStageIntLLROutputS2xD(151)(3);
  VNStageIntLLRInputS2xD(319)(2) <= CNStageIntLLROutputS2xD(151)(4);
  VNStageIntLLRInputS2xD(379)(1) <= CNStageIntLLROutputS2xD(151)(5);
  VNStageIntLLRInputS2xD(50)(2) <= CNStageIntLLROutputS2xD(152)(0);
  VNStageIntLLRInputS2xD(118)(2) <= CNStageIntLLROutputS2xD(152)(1);
  VNStageIntLLRInputS2xD(189)(1) <= CNStageIntLLROutputS2xD(152)(2);
  VNStageIntLLRInputS2xD(249)(0) <= CNStageIntLLROutputS2xD(152)(3);
  VNStageIntLLRInputS2xD(261)(2) <= CNStageIntLLROutputS2xD(152)(4);
  VNStageIntLLRInputS2xD(348)(2) <= CNStageIntLLROutputS2xD(152)(5);
  VNStageIntLLRInputS2xD(49)(2) <= CNStageIntLLROutputS2xD(153)(0);
  VNStageIntLLRInputS2xD(124)(1) <= CNStageIntLLROutputS2xD(153)(1);
  VNStageIntLLRInputS2xD(184)(2) <= CNStageIntLLROutputS2xD(153)(2);
  VNStageIntLLRInputS2xD(196)(2) <= CNStageIntLLROutputS2xD(153)(3);
  VNStageIntLLRInputS2xD(283)(2) <= CNStageIntLLROutputS2xD(153)(4);
  VNStageIntLLRInputS2xD(366)(2) <= CNStageIntLLROutputS2xD(153)(5);
  VNStageIntLLRInputS2xD(48)(1) <= CNStageIntLLROutputS2xD(154)(0);
  VNStageIntLLRInputS2xD(119)(2) <= CNStageIntLLROutputS2xD(154)(1);
  VNStageIntLLRInputS2xD(131)(1) <= CNStageIntLLROutputS2xD(154)(2);
  VNStageIntLLRInputS2xD(218)(2) <= CNStageIntLLROutputS2xD(154)(3);
  VNStageIntLLRInputS2xD(301)(2) <= CNStageIntLLROutputS2xD(154)(4);
  VNStageIntLLRInputS2xD(351)(1) <= CNStageIntLLROutputS2xD(154)(5);
  VNStageIntLLRInputS2xD(47)(1) <= CNStageIntLLROutputS2xD(155)(0);
  VNStageIntLLRInputS2xD(66)(2) <= CNStageIntLLROutputS2xD(155)(1);
  VNStageIntLLRInputS2xD(153)(2) <= CNStageIntLLROutputS2xD(155)(2);
  VNStageIntLLRInputS2xD(236)(2) <= CNStageIntLLROutputS2xD(155)(3);
  VNStageIntLLRInputS2xD(286)(2) <= CNStageIntLLROutputS2xD(155)(4);
  VNStageIntLLRInputS2xD(338)(2) <= CNStageIntLLROutputS2xD(155)(5);
  VNStageIntLLRInputS2xD(46)(2) <= CNStageIntLLROutputS2xD(156)(0);
  VNStageIntLLRInputS2xD(88)(2) <= CNStageIntLLROutputS2xD(156)(1);
  VNStageIntLLRInputS2xD(171)(1) <= CNStageIntLLROutputS2xD(156)(2);
  VNStageIntLLRInputS2xD(221)(2) <= CNStageIntLLROutputS2xD(156)(3);
  VNStageIntLLRInputS2xD(273)(2) <= CNStageIntLLROutputS2xD(156)(4);
  VNStageIntLLRInputS2xD(369)(1) <= CNStageIntLLROutputS2xD(156)(5);
  VNStageIntLLRInputS2xD(45)(2) <= CNStageIntLLROutputS2xD(157)(0);
  VNStageIntLLRInputS2xD(106)(1) <= CNStageIntLLROutputS2xD(157)(1);
  VNStageIntLLRInputS2xD(156)(2) <= CNStageIntLLROutputS2xD(157)(2);
  VNStageIntLLRInputS2xD(208)(2) <= CNStageIntLLROutputS2xD(157)(3);
  VNStageIntLLRInputS2xD(304)(2) <= CNStageIntLLROutputS2xD(157)(4);
  VNStageIntLLRInputS2xD(381)(1) <= CNStageIntLLROutputS2xD(157)(5);
  VNStageIntLLRInputS2xD(44)(2) <= CNStageIntLLROutputS2xD(158)(0);
  VNStageIntLLRInputS2xD(91)(2) <= CNStageIntLLROutputS2xD(158)(1);
  VNStageIntLLRInputS2xD(143)(2) <= CNStageIntLLROutputS2xD(158)(2);
  VNStageIntLLRInputS2xD(239)(2) <= CNStageIntLLROutputS2xD(158)(3);
  VNStageIntLLRInputS2xD(316)(1) <= CNStageIntLLROutputS2xD(158)(4);
  VNStageIntLLRInputS2xD(332)(2) <= CNStageIntLLROutputS2xD(158)(5);
  VNStageIntLLRInputS2xD(43)(1) <= CNStageIntLLROutputS2xD(159)(0);
  VNStageIntLLRInputS2xD(78)(2) <= CNStageIntLLROutputS2xD(159)(1);
  VNStageIntLLRInputS2xD(174)(2) <= CNStageIntLLROutputS2xD(159)(2);
  VNStageIntLLRInputS2xD(251)(1) <= CNStageIntLLROutputS2xD(159)(3);
  VNStageIntLLRInputS2xD(267)(2) <= CNStageIntLLROutputS2xD(159)(4);
  VNStageIntLLRInputS2xD(376)(2) <= CNStageIntLLROutputS2xD(159)(5);
  VNStageIntLLRInputS2xD(42)(2) <= CNStageIntLLROutputS2xD(160)(0);
  VNStageIntLLRInputS2xD(109)(2) <= CNStageIntLLROutputS2xD(160)(1);
  VNStageIntLLRInputS2xD(186)(1) <= CNStageIntLLROutputS2xD(160)(2);
  VNStageIntLLRInputS2xD(202)(2) <= CNStageIntLLROutputS2xD(160)(3);
  VNStageIntLLRInputS2xD(311)(2) <= CNStageIntLLROutputS2xD(160)(4);
  VNStageIntLLRInputS2xD(353)(2) <= CNStageIntLLROutputS2xD(160)(5);
  VNStageIntLLRInputS2xD(41)(2) <= CNStageIntLLROutputS2xD(161)(0);
  VNStageIntLLRInputS2xD(121)(1) <= CNStageIntLLROutputS2xD(161)(1);
  VNStageIntLLRInputS2xD(137)(2) <= CNStageIntLLROutputS2xD(161)(2);
  VNStageIntLLRInputS2xD(246)(2) <= CNStageIntLLROutputS2xD(161)(3);
  VNStageIntLLRInputS2xD(288)(2) <= CNStageIntLLROutputS2xD(161)(4);
  VNStageIntLLRInputS2xD(342)(2) <= CNStageIntLLROutputS2xD(161)(5);
  VNStageIntLLRInputS2xD(40)(2) <= CNStageIntLLROutputS2xD(162)(0);
  VNStageIntLLRInputS2xD(72)(2) <= CNStageIntLLROutputS2xD(162)(1);
  VNStageIntLLRInputS2xD(181)(2) <= CNStageIntLLROutputS2xD(162)(2);
  VNStageIntLLRInputS2xD(223)(2) <= CNStageIntLLROutputS2xD(162)(3);
  VNStageIntLLRInputS2xD(277)(2) <= CNStageIntLLROutputS2xD(162)(4);
  VNStageIntLLRInputS2xD(346)(2) <= CNStageIntLLROutputS2xD(162)(5);
  VNStageIntLLRInputS2xD(39)(2) <= CNStageIntLLROutputS2xD(163)(0);
  VNStageIntLLRInputS2xD(116)(1) <= CNStageIntLLROutputS2xD(163)(1);
  VNStageIntLLRInputS2xD(158)(2) <= CNStageIntLLROutputS2xD(163)(2);
  VNStageIntLLRInputS2xD(212)(2) <= CNStageIntLLROutputS2xD(163)(3);
  VNStageIntLLRInputS2xD(281)(2) <= CNStageIntLLROutputS2xD(163)(4);
  VNStageIntLLRInputS2xD(339)(2) <= CNStageIntLLROutputS2xD(163)(5);
  VNStageIntLLRInputS2xD(38)(2) <= CNStageIntLLROutputS2xD(164)(0);
  VNStageIntLLRInputS2xD(93)(2) <= CNStageIntLLROutputS2xD(164)(1);
  VNStageIntLLRInputS2xD(147)(2) <= CNStageIntLLROutputS2xD(164)(2);
  VNStageIntLLRInputS2xD(216)(2) <= CNStageIntLLROutputS2xD(164)(3);
  VNStageIntLLRInputS2xD(274)(1) <= CNStageIntLLROutputS2xD(164)(4);
  VNStageIntLLRInputS2xD(350)(2) <= CNStageIntLLROutputS2xD(164)(5);
  VNStageIntLLRInputS2xD(37)(2) <= CNStageIntLLROutputS2xD(165)(0);
  VNStageIntLLRInputS2xD(82)(2) <= CNStageIntLLROutputS2xD(165)(1);
  VNStageIntLLRInputS2xD(151)(2) <= CNStageIntLLROutputS2xD(165)(2);
  VNStageIntLLRInputS2xD(209)(2) <= CNStageIntLLROutputS2xD(165)(3);
  VNStageIntLLRInputS2xD(285)(2) <= CNStageIntLLROutputS2xD(165)(4);
  VNStageIntLLRInputS2xD(322)(2) <= CNStageIntLLROutputS2xD(165)(5);
  VNStageIntLLRInputS2xD(36)(2) <= CNStageIntLLROutputS2xD(166)(0);
  VNStageIntLLRInputS2xD(86)(1) <= CNStageIntLLROutputS2xD(166)(1);
  VNStageIntLLRInputS2xD(144)(2) <= CNStageIntLLROutputS2xD(166)(2);
  VNStageIntLLRInputS2xD(220)(2) <= CNStageIntLLROutputS2xD(166)(3);
  VNStageIntLLRInputS2xD(257)(2) <= CNStageIntLLROutputS2xD(166)(4);
  VNStageIntLLRInputS2xD(377)(1) <= CNStageIntLLROutputS2xD(166)(5);
  VNStageIntLLRInputS2xD(35)(2) <= CNStageIntLLROutputS2xD(167)(0);
  VNStageIntLLRInputS2xD(79)(2) <= CNStageIntLLROutputS2xD(167)(1);
  VNStageIntLLRInputS2xD(155)(2) <= CNStageIntLLROutputS2xD(167)(2);
  VNStageIntLLRInputS2xD(255)(2) <= CNStageIntLLROutputS2xD(167)(3);
  VNStageIntLLRInputS2xD(312)(2) <= CNStageIntLLROutputS2xD(167)(4);
  VNStageIntLLRInputS2xD(331)(2) <= CNStageIntLLROutputS2xD(167)(5);
  VNStageIntLLRInputS2xD(34)(2) <= CNStageIntLLROutputS2xD(168)(0);
  VNStageIntLLRInputS2xD(90)(2) <= CNStageIntLLROutputS2xD(168)(1);
  VNStageIntLLRInputS2xD(190)(0) <= CNStageIntLLROutputS2xD(168)(2);
  VNStageIntLLRInputS2xD(247)(2) <= CNStageIntLLROutputS2xD(168)(3);
  VNStageIntLLRInputS2xD(266)(1) <= CNStageIntLLROutputS2xD(168)(4);
  VNStageIntLLRInputS2xD(328)(2) <= CNStageIntLLROutputS2xD(168)(5);
  VNStageIntLLRInputS2xD(33)(2) <= CNStageIntLLROutputS2xD(169)(0);
  VNStageIntLLRInputS2xD(125)(1) <= CNStageIntLLROutputS2xD(169)(1);
  VNStageIntLLRInputS2xD(182)(2) <= CNStageIntLLROutputS2xD(169)(2);
  VNStageIntLLRInputS2xD(201)(2) <= CNStageIntLLROutputS2xD(169)(3);
  VNStageIntLLRInputS2xD(263)(2) <= CNStageIntLLROutputS2xD(169)(4);
  VNStageIntLLRInputS2xD(362)(2) <= CNStageIntLLROutputS2xD(169)(5);
  VNStageIntLLRInputS2xD(0)(2) <= CNStageIntLLROutputS2xD(170)(0);
  VNStageIntLLRInputS2xD(75)(2) <= CNStageIntLLROutputS2xD(170)(1);
  VNStageIntLLRInputS2xD(140)(2) <= CNStageIntLLROutputS2xD(170)(2);
  VNStageIntLLRInputS2xD(205)(0) <= CNStageIntLLROutputS2xD(170)(3);
  VNStageIntLLRInputS2xD(270)(2) <= CNStageIntLLROutputS2xD(170)(4);
  VNStageIntLLRInputS2xD(335)(2) <= CNStageIntLLROutputS2xD(170)(5);
  VNStageIntLLRInputS2xD(62)(2) <= CNStageIntLLROutputS2xD(171)(0);
  VNStageIntLLRInputS2xD(109)(3) <= CNStageIntLLROutputS2xD(171)(1);
  VNStageIntLLRInputS2xD(161)(3) <= CNStageIntLLROutputS2xD(171)(2);
  VNStageIntLLRInputS2xD(194)(3) <= CNStageIntLLROutputS2xD(171)(3);
  VNStageIntLLRInputS2xD(271)(2) <= CNStageIntLLROutputS2xD(171)(4);
  VNStageIntLLRInputS2xD(350)(3) <= CNStageIntLLROutputS2xD(171)(5);
  VNStageIntLLRInputS2xD(61)(2) <= CNStageIntLLROutputS2xD(172)(0);
  VNStageIntLLRInputS2xD(96)(3) <= CNStageIntLLROutputS2xD(172)(1);
  VNStageIntLLRInputS2xD(129)(3) <= CNStageIntLLROutputS2xD(172)(2);
  VNStageIntLLRInputS2xD(206)(2) <= CNStageIntLLROutputS2xD(172)(3);
  VNStageIntLLRInputS2xD(285)(3) <= CNStageIntLLROutputS2xD(172)(4);
  VNStageIntLLRInputS2xD(331)(3) <= CNStageIntLLROutputS2xD(172)(5);
  VNStageIntLLRInputS2xD(60)(2) <= CNStageIntLLROutputS2xD(173)(0);
  VNStageIntLLRInputS2xD(127)(3) <= CNStageIntLLROutputS2xD(173)(1);
  VNStageIntLLRInputS2xD(141)(1) <= CNStageIntLLROutputS2xD(173)(2);
  VNStageIntLLRInputS2xD(220)(3) <= CNStageIntLLROutputS2xD(173)(3);
  VNStageIntLLRInputS2xD(266)(2) <= CNStageIntLLROutputS2xD(173)(4);
  VNStageIntLLRInputS2xD(371)(2) <= CNStageIntLLROutputS2xD(173)(5);
  VNStageIntLLRInputS2xD(59)(1) <= CNStageIntLLROutputS2xD(174)(0);
  VNStageIntLLRInputS2xD(76)(3) <= CNStageIntLLROutputS2xD(174)(1);
  VNStageIntLLRInputS2xD(155)(3) <= CNStageIntLLROutputS2xD(174)(2);
  VNStageIntLLRInputS2xD(201)(3) <= CNStageIntLLROutputS2xD(174)(3);
  VNStageIntLLRInputS2xD(306)(3) <= CNStageIntLLROutputS2xD(174)(4);
  VNStageIntLLRInputS2xD(360)(3) <= CNStageIntLLROutputS2xD(174)(5);
  VNStageIntLLRInputS2xD(58)(2) <= CNStageIntLLROutputS2xD(175)(0);
  VNStageIntLLRInputS2xD(90)(3) <= CNStageIntLLROutputS2xD(175)(1);
  VNStageIntLLRInputS2xD(136)(3) <= CNStageIntLLROutputS2xD(175)(2);
  VNStageIntLLRInputS2xD(241)(2) <= CNStageIntLLROutputS2xD(175)(3);
  VNStageIntLLRInputS2xD(295)(3) <= CNStageIntLLROutputS2xD(175)(4);
  VNStageIntLLRInputS2xD(364)(3) <= CNStageIntLLROutputS2xD(175)(5);
  VNStageIntLLRInputS2xD(57)(2) <= CNStageIntLLROutputS2xD(176)(0);
  VNStageIntLLRInputS2xD(71)(2) <= CNStageIntLLROutputS2xD(176)(1);
  VNStageIntLLRInputS2xD(176)(3) <= CNStageIntLLROutputS2xD(176)(2);
  VNStageIntLLRInputS2xD(230)(2) <= CNStageIntLLROutputS2xD(176)(3);
  VNStageIntLLRInputS2xD(299)(2) <= CNStageIntLLROutputS2xD(176)(4);
  VNStageIntLLRInputS2xD(357)(3) <= CNStageIntLLROutputS2xD(176)(5);
  VNStageIntLLRInputS2xD(56)(3) <= CNStageIntLLROutputS2xD(177)(0);
  VNStageIntLLRInputS2xD(111)(3) <= CNStageIntLLROutputS2xD(177)(1);
  VNStageIntLLRInputS2xD(165)(3) <= CNStageIntLLROutputS2xD(177)(2);
  VNStageIntLLRInputS2xD(234)(3) <= CNStageIntLLROutputS2xD(177)(3);
  VNStageIntLLRInputS2xD(292)(3) <= CNStageIntLLROutputS2xD(177)(4);
  VNStageIntLLRInputS2xD(368)(1) <= CNStageIntLLROutputS2xD(177)(5);
  VNStageIntLLRInputS2xD(55)(3) <= CNStageIntLLROutputS2xD(178)(0);
  VNStageIntLLRInputS2xD(100)(3) <= CNStageIntLLROutputS2xD(178)(1);
  VNStageIntLLRInputS2xD(169)(3) <= CNStageIntLLROutputS2xD(178)(2);
  VNStageIntLLRInputS2xD(227)(3) <= CNStageIntLLROutputS2xD(178)(3);
  VNStageIntLLRInputS2xD(303)(3) <= CNStageIntLLROutputS2xD(178)(4);
  VNStageIntLLRInputS2xD(340)(3) <= CNStageIntLLROutputS2xD(178)(5);
  VNStageIntLLRInputS2xD(54)(3) <= CNStageIntLLROutputS2xD(179)(0);
  VNStageIntLLRInputS2xD(104)(3) <= CNStageIntLLROutputS2xD(179)(1);
  VNStageIntLLRInputS2xD(162)(3) <= CNStageIntLLROutputS2xD(179)(2);
  VNStageIntLLRInputS2xD(238)(3) <= CNStageIntLLROutputS2xD(179)(3);
  VNStageIntLLRInputS2xD(275)(3) <= CNStageIntLLROutputS2xD(179)(4);
  VNStageIntLLRInputS2xD(332)(3) <= CNStageIntLLROutputS2xD(179)(5);
  VNStageIntLLRInputS2xD(53)(2) <= CNStageIntLLROutputS2xD(180)(0);
  VNStageIntLLRInputS2xD(97)(3) <= CNStageIntLLROutputS2xD(180)(1);
  VNStageIntLLRInputS2xD(173)(3) <= CNStageIntLLROutputS2xD(180)(2);
  VNStageIntLLRInputS2xD(210)(3) <= CNStageIntLLROutputS2xD(180)(3);
  VNStageIntLLRInputS2xD(267)(3) <= CNStageIntLLROutputS2xD(180)(4);
  VNStageIntLLRInputS2xD(349)(2) <= CNStageIntLLROutputS2xD(180)(5);
  VNStageIntLLRInputS2xD(52)(2) <= CNStageIntLLROutputS2xD(181)(0);
  VNStageIntLLRInputS2xD(108)(3) <= CNStageIntLLROutputS2xD(181)(1);
  VNStageIntLLRInputS2xD(145)(3) <= CNStageIntLLROutputS2xD(181)(2);
  VNStageIntLLRInputS2xD(202)(3) <= CNStageIntLLROutputS2xD(181)(3);
  VNStageIntLLRInputS2xD(284)(3) <= CNStageIntLLROutputS2xD(181)(4);
  VNStageIntLLRInputS2xD(346)(3) <= CNStageIntLLROutputS2xD(181)(5);
  VNStageIntLLRInputS2xD(51)(2) <= CNStageIntLLROutputS2xD(182)(0);
  VNStageIntLLRInputS2xD(80)(3) <= CNStageIntLLROutputS2xD(182)(1);
  VNStageIntLLRInputS2xD(137)(3) <= CNStageIntLLROutputS2xD(182)(2);
  VNStageIntLLRInputS2xD(219)(3) <= CNStageIntLLROutputS2xD(182)(3);
  VNStageIntLLRInputS2xD(281)(3) <= CNStageIntLLROutputS2xD(182)(4);
  VNStageIntLLRInputS2xD(380)(2) <= CNStageIntLLROutputS2xD(182)(5);
  VNStageIntLLRInputS2xD(50)(3) <= CNStageIntLLROutputS2xD(183)(0);
  VNStageIntLLRInputS2xD(72)(3) <= CNStageIntLLROutputS2xD(183)(1);
  VNStageIntLLRInputS2xD(154)(2) <= CNStageIntLLROutputS2xD(183)(2);
  VNStageIntLLRInputS2xD(216)(3) <= CNStageIntLLROutputS2xD(183)(3);
  VNStageIntLLRInputS2xD(315)(2) <= CNStageIntLLROutputS2xD(183)(4);
  VNStageIntLLRInputS2xD(337)(3) <= CNStageIntLLROutputS2xD(183)(5);
  VNStageIntLLRInputS2xD(49)(3) <= CNStageIntLLROutputS2xD(184)(0);
  VNStageIntLLRInputS2xD(89)(3) <= CNStageIntLLROutputS2xD(184)(1);
  VNStageIntLLRInputS2xD(151)(3) <= CNStageIntLLROutputS2xD(184)(2);
  VNStageIntLLRInputS2xD(250)(2) <= CNStageIntLLROutputS2xD(184)(3);
  VNStageIntLLRInputS2xD(272)(3) <= CNStageIntLLROutputS2xD(184)(4);
  VNStageIntLLRInputS2xD(323)(2) <= CNStageIntLLROutputS2xD(184)(5);
  VNStageIntLLRInputS2xD(46)(3) <= CNStageIntLLROutputS2xD(185)(0);
  VNStageIntLLRInputS2xD(77)(1) <= CNStageIntLLROutputS2xD(185)(1);
  VNStageIntLLRInputS2xD(191)(3) <= CNStageIntLLROutputS2xD(185)(2);
  VNStageIntLLRInputS2xD(246)(3) <= CNStageIntLLROutputS2xD(185)(3);
  VNStageIntLLRInputS2xD(277)(3) <= CNStageIntLLROutputS2xD(185)(4);
  VNStageIntLLRInputS2xD(325)(3) <= CNStageIntLLROutputS2xD(185)(5);
  VNStageIntLLRInputS2xD(45)(3) <= CNStageIntLLROutputS2xD(186)(0);
  VNStageIntLLRInputS2xD(126)(2) <= CNStageIntLLROutputS2xD(186)(1);
  VNStageIntLLRInputS2xD(181)(3) <= CNStageIntLLROutputS2xD(186)(2);
  VNStageIntLLRInputS2xD(212)(3) <= CNStageIntLLROutputS2xD(186)(3);
  VNStageIntLLRInputS2xD(260)(3) <= CNStageIntLLROutputS2xD(186)(4);
  VNStageIntLLRInputS2xD(355)(3) <= CNStageIntLLROutputS2xD(186)(5);
  VNStageIntLLRInputS2xD(44)(3) <= CNStageIntLLROutputS2xD(187)(0);
  VNStageIntLLRInputS2xD(116)(2) <= CNStageIntLLROutputS2xD(187)(1);
  VNStageIntLLRInputS2xD(147)(3) <= CNStageIntLLROutputS2xD(187)(2);
  VNStageIntLLRInputS2xD(195)(2) <= CNStageIntLLROutputS2xD(187)(3);
  VNStageIntLLRInputS2xD(290)(3) <= CNStageIntLLROutputS2xD(187)(4);
  VNStageIntLLRInputS2xD(378)(2) <= CNStageIntLLROutputS2xD(187)(5);
  VNStageIntLLRInputS2xD(43)(2) <= CNStageIntLLROutputS2xD(188)(0);
  VNStageIntLLRInputS2xD(82)(3) <= CNStageIntLLROutputS2xD(188)(1);
  VNStageIntLLRInputS2xD(130)(3) <= CNStageIntLLROutputS2xD(188)(2);
  VNStageIntLLRInputS2xD(225)(3) <= CNStageIntLLROutputS2xD(188)(3);
  VNStageIntLLRInputS2xD(313)(1) <= CNStageIntLLROutputS2xD(188)(4);
  VNStageIntLLRInputS2xD(351)(2) <= CNStageIntLLROutputS2xD(188)(5);
  VNStageIntLLRInputS2xD(42)(3) <= CNStageIntLLROutputS2xD(189)(0);
  VNStageIntLLRInputS2xD(65)(3) <= CNStageIntLLROutputS2xD(189)(1);
  VNStageIntLLRInputS2xD(160)(3) <= CNStageIntLLROutputS2xD(189)(2);
  VNStageIntLLRInputS2xD(248)(3) <= CNStageIntLLROutputS2xD(189)(3);
  VNStageIntLLRInputS2xD(286)(3) <= CNStageIntLLROutputS2xD(189)(4);
  VNStageIntLLRInputS2xD(335)(3) <= CNStageIntLLROutputS2xD(189)(5);
  VNStageIntLLRInputS2xD(41)(3) <= CNStageIntLLROutputS2xD(190)(0);
  VNStageIntLLRInputS2xD(95)(3) <= CNStageIntLLROutputS2xD(190)(1);
  VNStageIntLLRInputS2xD(183)(2) <= CNStageIntLLROutputS2xD(190)(2);
  VNStageIntLLRInputS2xD(221)(3) <= CNStageIntLLROutputS2xD(190)(3);
  VNStageIntLLRInputS2xD(270)(3) <= CNStageIntLLROutputS2xD(190)(4);
  VNStageIntLLRInputS2xD(338)(3) <= CNStageIntLLROutputS2xD(190)(5);
  VNStageIntLLRInputS2xD(39)(3) <= CNStageIntLLROutputS2xD(191)(0);
  VNStageIntLLRInputS2xD(91)(3) <= CNStageIntLLROutputS2xD(191)(1);
  VNStageIntLLRInputS2xD(140)(3) <= CNStageIntLLROutputS2xD(191)(2);
  VNStageIntLLRInputS2xD(208)(3) <= CNStageIntLLROutputS2xD(191)(3);
  VNStageIntLLRInputS2xD(314)(0) <= CNStageIntLLROutputS2xD(191)(4);
  VNStageIntLLRInputS2xD(354)(3) <= CNStageIntLLROutputS2xD(191)(5);
  VNStageIntLLRInputS2xD(38)(3) <= CNStageIntLLROutputS2xD(192)(0);
  VNStageIntLLRInputS2xD(75)(3) <= CNStageIntLLROutputS2xD(192)(1);
  VNStageIntLLRInputS2xD(143)(3) <= CNStageIntLLROutputS2xD(192)(2);
  VNStageIntLLRInputS2xD(249)(1) <= CNStageIntLLROutputS2xD(192)(3);
  VNStageIntLLRInputS2xD(289)(3) <= CNStageIntLLROutputS2xD(192)(4);
  VNStageIntLLRInputS2xD(352)(3) <= CNStageIntLLROutputS2xD(192)(5);
  VNStageIntLLRInputS2xD(37)(3) <= CNStageIntLLROutputS2xD(193)(0);
  VNStageIntLLRInputS2xD(78)(3) <= CNStageIntLLROutputS2xD(193)(1);
  VNStageIntLLRInputS2xD(184)(3) <= CNStageIntLLROutputS2xD(193)(2);
  VNStageIntLLRInputS2xD(224)(3) <= CNStageIntLLROutputS2xD(193)(3);
  VNStageIntLLRInputS2xD(287)(3) <= CNStageIntLLROutputS2xD(193)(4);
  VNStageIntLLRInputS2xD(377)(2) <= CNStageIntLLROutputS2xD(193)(5);
  VNStageIntLLRInputS2xD(35)(3) <= CNStageIntLLROutputS2xD(194)(0);
  VNStageIntLLRInputS2xD(94)(2) <= CNStageIntLLROutputS2xD(194)(1);
  VNStageIntLLRInputS2xD(157)(3) <= CNStageIntLLROutputS2xD(194)(2);
  VNStageIntLLRInputS2xD(247)(3) <= CNStageIntLLROutputS2xD(194)(3);
  VNStageIntLLRInputS2xD(257)(3) <= CNStageIntLLROutputS2xD(194)(4);
  VNStageIntLLRInputS2xD(365)(3) <= CNStageIntLLROutputS2xD(194)(5);
  VNStageIntLLRInputS2xD(34)(3) <= CNStageIntLLROutputS2xD(195)(0);
  VNStageIntLLRInputS2xD(92)(3) <= CNStageIntLLROutputS2xD(195)(1);
  VNStageIntLLRInputS2xD(182)(3) <= CNStageIntLLROutputS2xD(195)(2);
  VNStageIntLLRInputS2xD(255)(3) <= CNStageIntLLROutputS2xD(195)(3);
  VNStageIntLLRInputS2xD(300)(3) <= CNStageIntLLROutputS2xD(195)(4);
  VNStageIntLLRInputS2xD(359)(3) <= CNStageIntLLROutputS2xD(195)(5);
  VNStageIntLLRInputS2xD(33)(3) <= CNStageIntLLROutputS2xD(196)(0);
  VNStageIntLLRInputS2xD(117)(3) <= CNStageIntLLROutputS2xD(196)(1);
  VNStageIntLLRInputS2xD(190)(1) <= CNStageIntLLROutputS2xD(196)(2);
  VNStageIntLLRInputS2xD(235)(2) <= CNStageIntLLROutputS2xD(196)(3);
  VNStageIntLLRInputS2xD(294)(3) <= CNStageIntLLROutputS2xD(196)(4);
  VNStageIntLLRInputS2xD(320)(2) <= CNStageIntLLROutputS2xD(196)(5);
  VNStageIntLLRInputS2xD(31)(2) <= CNStageIntLLROutputS2xD(197)(0);
  VNStageIntLLRInputS2xD(105)(2) <= CNStageIntLLROutputS2xD(197)(1);
  VNStageIntLLRInputS2xD(164)(3) <= CNStageIntLLROutputS2xD(197)(2);
  VNStageIntLLRInputS2xD(192)(3) <= CNStageIntLLROutputS2xD(197)(3);
  VNStageIntLLRInputS2xD(293)(3) <= CNStageIntLLROutputS2xD(197)(4);
  VNStageIntLLRInputS2xD(363)(2) <= CNStageIntLLROutputS2xD(197)(5);
  VNStageIntLLRInputS2xD(30)(3) <= CNStageIntLLROutputS2xD(198)(0);
  VNStageIntLLRInputS2xD(99)(3) <= CNStageIntLLROutputS2xD(198)(1);
  VNStageIntLLRInputS2xD(128)(3) <= CNStageIntLLROutputS2xD(198)(2);
  VNStageIntLLRInputS2xD(228)(3) <= CNStageIntLLROutputS2xD(198)(3);
  VNStageIntLLRInputS2xD(298)(3) <= CNStageIntLLROutputS2xD(198)(4);
  VNStageIntLLRInputS2xD(382)(2) <= CNStageIntLLROutputS2xD(198)(5);
  VNStageIntLLRInputS2xD(28)(3) <= CNStageIntLLROutputS2xD(199)(0);
  VNStageIntLLRInputS2xD(98)(2) <= CNStageIntLLROutputS2xD(199)(1);
  VNStageIntLLRInputS2xD(168)(2) <= CNStageIntLLROutputS2xD(199)(2);
  VNStageIntLLRInputS2xD(252)(2) <= CNStageIntLLROutputS2xD(199)(3);
  VNStageIntLLRInputS2xD(308)(1) <= CNStageIntLLROutputS2xD(199)(4);
  VNStageIntLLRInputS2xD(347)(3) <= CNStageIntLLROutputS2xD(199)(5);
  VNStageIntLLRInputS2xD(27)(3) <= CNStageIntLLROutputS2xD(200)(0);
  VNStageIntLLRInputS2xD(103)(3) <= CNStageIntLLROutputS2xD(200)(1);
  VNStageIntLLRInputS2xD(187)(2) <= CNStageIntLLROutputS2xD(200)(2);
  VNStageIntLLRInputS2xD(243)(3) <= CNStageIntLLROutputS2xD(200)(3);
  VNStageIntLLRInputS2xD(282)(3) <= CNStageIntLLROutputS2xD(200)(4);
  VNStageIntLLRInputS2xD(348)(3) <= CNStageIntLLROutputS2xD(200)(5);
  VNStageIntLLRInputS2xD(26)(3) <= CNStageIntLLROutputS2xD(201)(0);
  VNStageIntLLRInputS2xD(122)(2) <= CNStageIntLLROutputS2xD(201)(1);
  VNStageIntLLRInputS2xD(178)(3) <= CNStageIntLLROutputS2xD(201)(2);
  VNStageIntLLRInputS2xD(217)(3) <= CNStageIntLLROutputS2xD(201)(3);
  VNStageIntLLRInputS2xD(283)(3) <= CNStageIntLLROutputS2xD(201)(4);
  VNStageIntLLRInputS2xD(372)(2) <= CNStageIntLLROutputS2xD(201)(5);
  VNStageIntLLRInputS2xD(25)(3) <= CNStageIntLLROutputS2xD(202)(0);
  VNStageIntLLRInputS2xD(113)(3) <= CNStageIntLLROutputS2xD(202)(1);
  VNStageIntLLRInputS2xD(152)(3) <= CNStageIntLLROutputS2xD(202)(2);
  VNStageIntLLRInputS2xD(218)(3) <= CNStageIntLLROutputS2xD(202)(3);
  VNStageIntLLRInputS2xD(307)(3) <= CNStageIntLLROutputS2xD(202)(4);
  VNStageIntLLRInputS2xD(330)(3) <= CNStageIntLLROutputS2xD(202)(5);
  VNStageIntLLRInputS2xD(24)(3) <= CNStageIntLLROutputS2xD(203)(0);
  VNStageIntLLRInputS2xD(87)(3) <= CNStageIntLLROutputS2xD(203)(1);
  VNStageIntLLRInputS2xD(153)(3) <= CNStageIntLLROutputS2xD(203)(2);
  VNStageIntLLRInputS2xD(242)(3) <= CNStageIntLLROutputS2xD(203)(3);
  VNStageIntLLRInputS2xD(265)(2) <= CNStageIntLLROutputS2xD(203)(4);
  VNStageIntLLRInputS2xD(326)(2) <= CNStageIntLLROutputS2xD(203)(5);
  VNStageIntLLRInputS2xD(23)(3) <= CNStageIntLLROutputS2xD(204)(0);
  VNStageIntLLRInputS2xD(88)(3) <= CNStageIntLLROutputS2xD(204)(1);
  VNStageIntLLRInputS2xD(177)(3) <= CNStageIntLLROutputS2xD(204)(2);
  VNStageIntLLRInputS2xD(200)(3) <= CNStageIntLLROutputS2xD(204)(3);
  VNStageIntLLRInputS2xD(261)(3) <= CNStageIntLLROutputS2xD(204)(4);
  VNStageIntLLRInputS2xD(341)(3) <= CNStageIntLLROutputS2xD(204)(5);
  VNStageIntLLRInputS2xD(22)(3) <= CNStageIntLLROutputS2xD(205)(0);
  VNStageIntLLRInputS2xD(112)(3) <= CNStageIntLLROutputS2xD(205)(1);
  VNStageIntLLRInputS2xD(135)(3) <= CNStageIntLLROutputS2xD(205)(2);
  VNStageIntLLRInputS2xD(196)(3) <= CNStageIntLLROutputS2xD(205)(3);
  VNStageIntLLRInputS2xD(276)(3) <= CNStageIntLLROutputS2xD(205)(4);
  VNStageIntLLRInputS2xD(367)(3) <= CNStageIntLLROutputS2xD(205)(5);
  VNStageIntLLRInputS2xD(21)(3) <= CNStageIntLLROutputS2xD(206)(0);
  VNStageIntLLRInputS2xD(70)(3) <= CNStageIntLLROutputS2xD(206)(1);
  VNStageIntLLRInputS2xD(131)(2) <= CNStageIntLLROutputS2xD(206)(2);
  VNStageIntLLRInputS2xD(211)(3) <= CNStageIntLLROutputS2xD(206)(3);
  VNStageIntLLRInputS2xD(302)(3) <= CNStageIntLLROutputS2xD(206)(4);
  VNStageIntLLRInputS2xD(343)(3) <= CNStageIntLLROutputS2xD(206)(5);
  VNStageIntLLRInputS2xD(18)(3) <= CNStageIntLLROutputS2xD(207)(0);
  VNStageIntLLRInputS2xD(107)(2) <= CNStageIntLLROutputS2xD(207)(1);
  VNStageIntLLRInputS2xD(148)(3) <= CNStageIntLLROutputS2xD(207)(2);
  VNStageIntLLRInputS2xD(245)(3) <= CNStageIntLLROutputS2xD(207)(3);
  VNStageIntLLRInputS2xD(263)(3) <= CNStageIntLLROutputS2xD(207)(4);
  VNStageIntLLRInputS2xD(361)(3) <= CNStageIntLLROutputS2xD(207)(5);
  VNStageIntLLRInputS2xD(17)(3) <= CNStageIntLLROutputS2xD(208)(0);
  VNStageIntLLRInputS2xD(83)(3) <= CNStageIntLLROutputS2xD(208)(1);
  VNStageIntLLRInputS2xD(180)(1) <= CNStageIntLLROutputS2xD(208)(2);
  VNStageIntLLRInputS2xD(198)(3) <= CNStageIntLLROutputS2xD(208)(3);
  VNStageIntLLRInputS2xD(296)(3) <= CNStageIntLLROutputS2xD(208)(4);
  VNStageIntLLRInputS2xD(370)(2) <= CNStageIntLLROutputS2xD(208)(5);
  VNStageIntLLRInputS2xD(16)(2) <= CNStageIntLLROutputS2xD(209)(0);
  VNStageIntLLRInputS2xD(115)(3) <= CNStageIntLLROutputS2xD(209)(1);
  VNStageIntLLRInputS2xD(133)(1) <= CNStageIntLLROutputS2xD(209)(2);
  VNStageIntLLRInputS2xD(231)(2) <= CNStageIntLLROutputS2xD(209)(3);
  VNStageIntLLRInputS2xD(305)(3) <= CNStageIntLLROutputS2xD(209)(4);
  VNStageIntLLRInputS2xD(383)(3) <= CNStageIntLLROutputS2xD(209)(5);
  VNStageIntLLRInputS2xD(15)(3) <= CNStageIntLLROutputS2xD(210)(0);
  VNStageIntLLRInputS2xD(68)(2) <= CNStageIntLLROutputS2xD(210)(1);
  VNStageIntLLRInputS2xD(166)(3) <= CNStageIntLLROutputS2xD(210)(2);
  VNStageIntLLRInputS2xD(240)(3) <= CNStageIntLLROutputS2xD(210)(3);
  VNStageIntLLRInputS2xD(318)(1) <= CNStageIntLLROutputS2xD(210)(4);
  VNStageIntLLRInputS2xD(362)(3) <= CNStageIntLLROutputS2xD(210)(5);
  VNStageIntLLRInputS2xD(14)(3) <= CNStageIntLLROutputS2xD(211)(0);
  VNStageIntLLRInputS2xD(101)(3) <= CNStageIntLLROutputS2xD(211)(1);
  VNStageIntLLRInputS2xD(175)(3) <= CNStageIntLLROutputS2xD(211)(2);
  VNStageIntLLRInputS2xD(253)(2) <= CNStageIntLLROutputS2xD(211)(3);
  VNStageIntLLRInputS2xD(297)(3) <= CNStageIntLLROutputS2xD(211)(4);
  VNStageIntLLRInputS2xD(327)(3) <= CNStageIntLLROutputS2xD(211)(5);
  VNStageIntLLRInputS2xD(13)(2) <= CNStageIntLLROutputS2xD(212)(0);
  VNStageIntLLRInputS2xD(110)(3) <= CNStageIntLLROutputS2xD(212)(1);
  VNStageIntLLRInputS2xD(188)(1) <= CNStageIntLLROutputS2xD(212)(2);
  VNStageIntLLRInputS2xD(232)(2) <= CNStageIntLLROutputS2xD(212)(3);
  VNStageIntLLRInputS2xD(262)(3) <= CNStageIntLLROutputS2xD(212)(4);
  VNStageIntLLRInputS2xD(329)(3) <= CNStageIntLLROutputS2xD(212)(5);
  VNStageIntLLRInputS2xD(12)(3) <= CNStageIntLLROutputS2xD(213)(0);
  VNStageIntLLRInputS2xD(123)(2) <= CNStageIntLLROutputS2xD(213)(1);
  VNStageIntLLRInputS2xD(167)(3) <= CNStageIntLLROutputS2xD(213)(2);
  VNStageIntLLRInputS2xD(197)(3) <= CNStageIntLLROutputS2xD(213)(3);
  VNStageIntLLRInputS2xD(264)(3) <= CNStageIntLLROutputS2xD(213)(4);
  VNStageIntLLRInputS2xD(374)(3) <= CNStageIntLLROutputS2xD(213)(5);
  VNStageIntLLRInputS2xD(11)(3) <= CNStageIntLLROutputS2xD(214)(0);
  VNStageIntLLRInputS2xD(102)(3) <= CNStageIntLLROutputS2xD(214)(1);
  VNStageIntLLRInputS2xD(132)(2) <= CNStageIntLLROutputS2xD(214)(2);
  VNStageIntLLRInputS2xD(199)(3) <= CNStageIntLLROutputS2xD(214)(3);
  VNStageIntLLRInputS2xD(309)(3) <= CNStageIntLLROutputS2xD(214)(4);
  VNStageIntLLRInputS2xD(381)(2) <= CNStageIntLLROutputS2xD(214)(5);
  VNStageIntLLRInputS2xD(9)(3) <= CNStageIntLLROutputS2xD(215)(0);
  VNStageIntLLRInputS2xD(69)(3) <= CNStageIntLLROutputS2xD(215)(1);
  VNStageIntLLRInputS2xD(179)(3) <= CNStageIntLLROutputS2xD(215)(2);
  VNStageIntLLRInputS2xD(251)(2) <= CNStageIntLLROutputS2xD(215)(3);
  VNStageIntLLRInputS2xD(280)(3) <= CNStageIntLLROutputS2xD(215)(4);
  VNStageIntLLRInputS2xD(333)(2) <= CNStageIntLLROutputS2xD(215)(5);
  VNStageIntLLRInputS2xD(8)(2) <= CNStageIntLLROutputS2xD(216)(0);
  VNStageIntLLRInputS2xD(114)(3) <= CNStageIntLLROutputS2xD(216)(1);
  VNStageIntLLRInputS2xD(186)(2) <= CNStageIntLLROutputS2xD(216)(2);
  VNStageIntLLRInputS2xD(215)(3) <= CNStageIntLLROutputS2xD(216)(3);
  VNStageIntLLRInputS2xD(268)(3) <= CNStageIntLLROutputS2xD(216)(4);
  VNStageIntLLRInputS2xD(339)(3) <= CNStageIntLLROutputS2xD(216)(5);
  VNStageIntLLRInputS2xD(7)(3) <= CNStageIntLLROutputS2xD(217)(0);
  VNStageIntLLRInputS2xD(121)(2) <= CNStageIntLLROutputS2xD(217)(1);
  VNStageIntLLRInputS2xD(150)(3) <= CNStageIntLLROutputS2xD(217)(2);
  VNStageIntLLRInputS2xD(203)(3) <= CNStageIntLLROutputS2xD(217)(3);
  VNStageIntLLRInputS2xD(274)(2) <= CNStageIntLLROutputS2xD(217)(4);
  VNStageIntLLRInputS2xD(334)(2) <= CNStageIntLLROutputS2xD(217)(5);
  VNStageIntLLRInputS2xD(6)(3) <= CNStageIntLLROutputS2xD(218)(0);
  VNStageIntLLRInputS2xD(85)(2) <= CNStageIntLLROutputS2xD(218)(1);
  VNStageIntLLRInputS2xD(138)(3) <= CNStageIntLLROutputS2xD(218)(2);
  VNStageIntLLRInputS2xD(209)(3) <= CNStageIntLLROutputS2xD(218)(3);
  VNStageIntLLRInputS2xD(269)(2) <= CNStageIntLLROutputS2xD(218)(4);
  VNStageIntLLRInputS2xD(344)(3) <= CNStageIntLLROutputS2xD(218)(5);
  VNStageIntLLRInputS2xD(5)(3) <= CNStageIntLLROutputS2xD(219)(0);
  VNStageIntLLRInputS2xD(73)(3) <= CNStageIntLLROutputS2xD(219)(1);
  VNStageIntLLRInputS2xD(144)(3) <= CNStageIntLLROutputS2xD(219)(2);
  VNStageIntLLRInputS2xD(204)(3) <= CNStageIntLLROutputS2xD(219)(3);
  VNStageIntLLRInputS2xD(279)(3) <= CNStageIntLLROutputS2xD(219)(4);
  VNStageIntLLRInputS2xD(366)(3) <= CNStageIntLLROutputS2xD(219)(5);
  VNStageIntLLRInputS2xD(4)(2) <= CNStageIntLLROutputS2xD(220)(0);
  VNStageIntLLRInputS2xD(79)(3) <= CNStageIntLLROutputS2xD(220)(1);
  VNStageIntLLRInputS2xD(139)(3) <= CNStageIntLLROutputS2xD(220)(2);
  VNStageIntLLRInputS2xD(214)(3) <= CNStageIntLLROutputS2xD(220)(3);
  VNStageIntLLRInputS2xD(301)(3) <= CNStageIntLLROutputS2xD(220)(4);
  VNStageIntLLRInputS2xD(321)(3) <= CNStageIntLLROutputS2xD(220)(5);
  VNStageIntLLRInputS2xD(3)(2) <= CNStageIntLLROutputS2xD(221)(0);
  VNStageIntLLRInputS2xD(74)(3) <= CNStageIntLLROutputS2xD(221)(1);
  VNStageIntLLRInputS2xD(149)(3) <= CNStageIntLLROutputS2xD(221)(2);
  VNStageIntLLRInputS2xD(236)(3) <= CNStageIntLLROutputS2xD(221)(3);
  VNStageIntLLRInputS2xD(319)(3) <= CNStageIntLLROutputS2xD(221)(4);
  VNStageIntLLRInputS2xD(369)(2) <= CNStageIntLLROutputS2xD(221)(5);
  VNStageIntLLRInputS2xD(2)(3) <= CNStageIntLLROutputS2xD(222)(0);
  VNStageIntLLRInputS2xD(84)(3) <= CNStageIntLLROutputS2xD(222)(1);
  VNStageIntLLRInputS2xD(171)(2) <= CNStageIntLLROutputS2xD(222)(2);
  VNStageIntLLRInputS2xD(254)(1) <= CNStageIntLLROutputS2xD(222)(3);
  VNStageIntLLRInputS2xD(304)(3) <= CNStageIntLLROutputS2xD(222)(4);
  VNStageIntLLRInputS2xD(356)(3) <= CNStageIntLLROutputS2xD(222)(5);
  VNStageIntLLRInputS2xD(1)(2) <= CNStageIntLLROutputS2xD(223)(0);
  VNStageIntLLRInputS2xD(106)(2) <= CNStageIntLLROutputS2xD(223)(1);
  VNStageIntLLRInputS2xD(189)(2) <= CNStageIntLLROutputS2xD(223)(2);
  VNStageIntLLRInputS2xD(239)(3) <= CNStageIntLLROutputS2xD(223)(3);
  VNStageIntLLRInputS2xD(291)(3) <= CNStageIntLLROutputS2xD(223)(4);
  VNStageIntLLRInputS2xD(324)(3) <= CNStageIntLLROutputS2xD(223)(5);
  VNStageIntLLRInputS2xD(0)(3) <= CNStageIntLLROutputS2xD(224)(0);
  VNStageIntLLRInputS2xD(93)(3) <= CNStageIntLLROutputS2xD(224)(1);
  VNStageIntLLRInputS2xD(158)(3) <= CNStageIntLLROutputS2xD(224)(2);
  VNStageIntLLRInputS2xD(223)(3) <= CNStageIntLLROutputS2xD(224)(3);
  VNStageIntLLRInputS2xD(288)(3) <= CNStageIntLLROutputS2xD(224)(4);
  VNStageIntLLRInputS2xD(353)(3) <= CNStageIntLLROutputS2xD(224)(5);
  VNStageIntLLRInputS2xD(18)(4) <= CNStageIntLLROutputS2xD(225)(0);
  VNStageIntLLRInputS2xD(110)(4) <= CNStageIntLLROutputS2xD(225)(1);
  VNStageIntLLRInputS2xD(167)(4) <= CNStageIntLLROutputS2xD(225)(2);
  VNStageIntLLRInputS2xD(249)(2) <= CNStageIntLLROutputS2xD(225)(3);
  VNStageIntLLRInputS2xD(311)(3) <= CNStageIntLLROutputS2xD(225)(4);
  VNStageIntLLRInputS2xD(347)(4) <= CNStageIntLLROutputS2xD(225)(5);
  VNStageIntLLRInputS2xD(17)(4) <= CNStageIntLLROutputS2xD(226)(0);
  VNStageIntLLRInputS2xD(102)(4) <= CNStageIntLLROutputS2xD(226)(1);
  VNStageIntLLRInputS2xD(184)(4) <= CNStageIntLLROutputS2xD(226)(2);
  VNStageIntLLRInputS2xD(246)(4) <= CNStageIntLLROutputS2xD(226)(3);
  VNStageIntLLRInputS2xD(282)(4) <= CNStageIntLLROutputS2xD(226)(4);
  VNStageIntLLRInputS2xD(367)(4) <= CNStageIntLLROutputS2xD(226)(5);
  VNStageIntLLRInputS2xD(16)(3) <= CNStageIntLLROutputS2xD(227)(0);
  VNStageIntLLRInputS2xD(119)(3) <= CNStageIntLLROutputS2xD(227)(1);
  VNStageIntLLRInputS2xD(181)(4) <= CNStageIntLLROutputS2xD(227)(2);
  VNStageIntLLRInputS2xD(217)(4) <= CNStageIntLLROutputS2xD(227)(3);
  VNStageIntLLRInputS2xD(302)(4) <= CNStageIntLLROutputS2xD(227)(4);
  VNStageIntLLRInputS2xD(353)(4) <= CNStageIntLLROutputS2xD(227)(5);
  VNStageIntLLRInputS2xD(15)(4) <= CNStageIntLLROutputS2xD(228)(0);
  VNStageIntLLRInputS2xD(116)(3) <= CNStageIntLLROutputS2xD(228)(1);
  VNStageIntLLRInputS2xD(152)(4) <= CNStageIntLLROutputS2xD(228)(2);
  VNStageIntLLRInputS2xD(237)(3) <= CNStageIntLLROutputS2xD(228)(3);
  VNStageIntLLRInputS2xD(288)(4) <= CNStageIntLLROutputS2xD(228)(4);
  VNStageIntLLRInputS2xD(343)(4) <= CNStageIntLLROutputS2xD(228)(5);
  VNStageIntLLRInputS2xD(14)(4) <= CNStageIntLLROutputS2xD(229)(0);
  VNStageIntLLRInputS2xD(87)(4) <= CNStageIntLLROutputS2xD(229)(1);
  VNStageIntLLRInputS2xD(172)(3) <= CNStageIntLLROutputS2xD(229)(2);
  VNStageIntLLRInputS2xD(223)(4) <= CNStageIntLLROutputS2xD(229)(3);
  VNStageIntLLRInputS2xD(278)(3) <= CNStageIntLLROutputS2xD(229)(4);
  VNStageIntLLRInputS2xD(372)(3) <= CNStageIntLLROutputS2xD(229)(5);
  VNStageIntLLRInputS2xD(13)(3) <= CNStageIntLLROutputS2xD(230)(0);
  VNStageIntLLRInputS2xD(107)(3) <= CNStageIntLLROutputS2xD(230)(1);
  VNStageIntLLRInputS2xD(158)(4) <= CNStageIntLLROutputS2xD(230)(2);
  VNStageIntLLRInputS2xD(213)(3) <= CNStageIntLLROutputS2xD(230)(3);
  VNStageIntLLRInputS2xD(307)(4) <= CNStageIntLLROutputS2xD(230)(4);
  VNStageIntLLRInputS2xD(355)(4) <= CNStageIntLLROutputS2xD(230)(5);
  VNStageIntLLRInputS2xD(12)(4) <= CNStageIntLLROutputS2xD(231)(0);
  VNStageIntLLRInputS2xD(93)(4) <= CNStageIntLLROutputS2xD(231)(1);
  VNStageIntLLRInputS2xD(148)(4) <= CNStageIntLLROutputS2xD(231)(2);
  VNStageIntLLRInputS2xD(242)(4) <= CNStageIntLLROutputS2xD(231)(3);
  VNStageIntLLRInputS2xD(290)(4) <= CNStageIntLLROutputS2xD(231)(4);
  VNStageIntLLRInputS2xD(322)(3) <= CNStageIntLLROutputS2xD(231)(5);
  VNStageIntLLRInputS2xD(11)(4) <= CNStageIntLLROutputS2xD(232)(0);
  VNStageIntLLRInputS2xD(83)(4) <= CNStageIntLLROutputS2xD(232)(1);
  VNStageIntLLRInputS2xD(177)(4) <= CNStageIntLLROutputS2xD(232)(2);
  VNStageIntLLRInputS2xD(225)(4) <= CNStageIntLLROutputS2xD(232)(3);
  VNStageIntLLRInputS2xD(257)(4) <= CNStageIntLLROutputS2xD(232)(4);
  VNStageIntLLRInputS2xD(345)(3) <= CNStageIntLLROutputS2xD(232)(5);
  VNStageIntLLRInputS2xD(10)(3) <= CNStageIntLLROutputS2xD(233)(0);
  VNStageIntLLRInputS2xD(112)(4) <= CNStageIntLLROutputS2xD(233)(1);
  VNStageIntLLRInputS2xD(160)(4) <= CNStageIntLLROutputS2xD(233)(2);
  VNStageIntLLRInputS2xD(255)(4) <= CNStageIntLLROutputS2xD(233)(3);
  VNStageIntLLRInputS2xD(280)(4) <= CNStageIntLLROutputS2xD(233)(4);
  VNStageIntLLRInputS2xD(381)(3) <= CNStageIntLLROutputS2xD(233)(5);
  VNStageIntLLRInputS2xD(9)(4) <= CNStageIntLLROutputS2xD(234)(0);
  VNStageIntLLRInputS2xD(95)(4) <= CNStageIntLLROutputS2xD(234)(1);
  VNStageIntLLRInputS2xD(190)(2) <= CNStageIntLLROutputS2xD(234)(2);
  VNStageIntLLRInputS2xD(215)(4) <= CNStageIntLLROutputS2xD(234)(3);
  VNStageIntLLRInputS2xD(316)(2) <= CNStageIntLLROutputS2xD(234)(4);
  VNStageIntLLRInputS2xD(365)(4) <= CNStageIntLLROutputS2xD(234)(5);
  VNStageIntLLRInputS2xD(7)(4) <= CNStageIntLLROutputS2xD(235)(0);
  VNStageIntLLRInputS2xD(85)(3) <= CNStageIntLLROutputS2xD(235)(1);
  VNStageIntLLRInputS2xD(186)(3) <= CNStageIntLLROutputS2xD(235)(2);
  VNStageIntLLRInputS2xD(235)(3) <= CNStageIntLLROutputS2xD(235)(3);
  VNStageIntLLRInputS2xD(303)(4) <= CNStageIntLLROutputS2xD(235)(4);
  VNStageIntLLRInputS2xD(346)(4) <= CNStageIntLLROutputS2xD(235)(5);
  VNStageIntLLRInputS2xD(6)(4) <= CNStageIntLLROutputS2xD(236)(0);
  VNStageIntLLRInputS2xD(121)(3) <= CNStageIntLLROutputS2xD(236)(1);
  VNStageIntLLRInputS2xD(170)(3) <= CNStageIntLLROutputS2xD(236)(2);
  VNStageIntLLRInputS2xD(238)(4) <= CNStageIntLLROutputS2xD(236)(3);
  VNStageIntLLRInputS2xD(281)(4) <= CNStageIntLLROutputS2xD(236)(4);
  VNStageIntLLRInputS2xD(321)(4) <= CNStageIntLLROutputS2xD(236)(5);
  VNStageIntLLRInputS2xD(5)(4) <= CNStageIntLLROutputS2xD(237)(0);
  VNStageIntLLRInputS2xD(105)(3) <= CNStageIntLLROutputS2xD(237)(1);
  VNStageIntLLRInputS2xD(173)(4) <= CNStageIntLLROutputS2xD(237)(2);
  VNStageIntLLRInputS2xD(216)(4) <= CNStageIntLLROutputS2xD(237)(3);
  VNStageIntLLRInputS2xD(319)(4) <= CNStageIntLLROutputS2xD(237)(4);
  VNStageIntLLRInputS2xD(382)(3) <= CNStageIntLLROutputS2xD(237)(5);
  VNStageIntLLRInputS2xD(4)(3) <= CNStageIntLLROutputS2xD(238)(0);
  VNStageIntLLRInputS2xD(108)(4) <= CNStageIntLLROutputS2xD(238)(1);
  VNStageIntLLRInputS2xD(151)(4) <= CNStageIntLLROutputS2xD(238)(2);
  VNStageIntLLRInputS2xD(254)(2) <= CNStageIntLLROutputS2xD(238)(3);
  VNStageIntLLRInputS2xD(317)(1) <= CNStageIntLLROutputS2xD(238)(4);
  VNStageIntLLRInputS2xD(344)(4) <= CNStageIntLLROutputS2xD(238)(5);
  VNStageIntLLRInputS2xD(3)(3) <= CNStageIntLLROutputS2xD(239)(0);
  VNStageIntLLRInputS2xD(86)(2) <= CNStageIntLLROutputS2xD(239)(1);
  VNStageIntLLRInputS2xD(189)(3) <= CNStageIntLLROutputS2xD(239)(2);
  VNStageIntLLRInputS2xD(252)(3) <= CNStageIntLLROutputS2xD(239)(3);
  VNStageIntLLRInputS2xD(279)(4) <= CNStageIntLLROutputS2xD(239)(4);
  VNStageIntLLRInputS2xD(352)(4) <= CNStageIntLLROutputS2xD(239)(5);
  VNStageIntLLRInputS2xD(2)(4) <= CNStageIntLLROutputS2xD(240)(0);
  VNStageIntLLRInputS2xD(124)(2) <= CNStageIntLLROutputS2xD(240)(1);
  VNStageIntLLRInputS2xD(187)(3) <= CNStageIntLLROutputS2xD(240)(2);
  VNStageIntLLRInputS2xD(214)(4) <= CNStageIntLLROutputS2xD(240)(3);
  VNStageIntLLRInputS2xD(287)(4) <= CNStageIntLLROutputS2xD(240)(4);
  VNStageIntLLRInputS2xD(332)(4) <= CNStageIntLLROutputS2xD(240)(5);
  VNStageIntLLRInputS2xD(1)(3) <= CNStageIntLLROutputS2xD(241)(0);
  VNStageIntLLRInputS2xD(122)(3) <= CNStageIntLLROutputS2xD(241)(1);
  VNStageIntLLRInputS2xD(149)(4) <= CNStageIntLLROutputS2xD(241)(2);
  VNStageIntLLRInputS2xD(222)(2) <= CNStageIntLLROutputS2xD(241)(3);
  VNStageIntLLRInputS2xD(267)(4) <= CNStageIntLLROutputS2xD(241)(4);
  VNStageIntLLRInputS2xD(326)(3) <= CNStageIntLLROutputS2xD(241)(5);
  VNStageIntLLRInputS2xD(62)(3) <= CNStageIntLLROutputS2xD(242)(0);
  VNStageIntLLRInputS2xD(92)(4) <= CNStageIntLLROutputS2xD(242)(1);
  VNStageIntLLRInputS2xD(137)(4) <= CNStageIntLLROutputS2xD(242)(2);
  VNStageIntLLRInputS2xD(196)(4) <= CNStageIntLLROutputS2xD(242)(3);
  VNStageIntLLRInputS2xD(256)(3) <= CNStageIntLLROutputS2xD(242)(4);
  VNStageIntLLRInputS2xD(325)(4) <= CNStageIntLLROutputS2xD(242)(5);
  VNStageIntLLRInputS2xD(61)(3) <= CNStageIntLLROutputS2xD(243)(0);
  VNStageIntLLRInputS2xD(72)(4) <= CNStageIntLLROutputS2xD(243)(1);
  VNStageIntLLRInputS2xD(131)(3) <= CNStageIntLLROutputS2xD(243)(2);
  VNStageIntLLRInputS2xD(192)(4) <= CNStageIntLLROutputS2xD(243)(3);
  VNStageIntLLRInputS2xD(260)(4) <= CNStageIntLLROutputS2xD(243)(4);
  VNStageIntLLRInputS2xD(330)(4) <= CNStageIntLLROutputS2xD(243)(5);
  VNStageIntLLRInputS2xD(60)(3) <= CNStageIntLLROutputS2xD(244)(0);
  VNStageIntLLRInputS2xD(66)(3) <= CNStageIntLLROutputS2xD(244)(1);
  VNStageIntLLRInputS2xD(128)(4) <= CNStageIntLLROutputS2xD(244)(2);
  VNStageIntLLRInputS2xD(195)(3) <= CNStageIntLLROutputS2xD(244)(3);
  VNStageIntLLRInputS2xD(265)(3) <= CNStageIntLLROutputS2xD(244)(4);
  VNStageIntLLRInputS2xD(349)(3) <= CNStageIntLLROutputS2xD(244)(5);
  VNStageIntLLRInputS2xD(59)(2) <= CNStageIntLLROutputS2xD(245)(0);
  VNStageIntLLRInputS2xD(64)(3) <= CNStageIntLLROutputS2xD(245)(1);
  VNStageIntLLRInputS2xD(130)(4) <= CNStageIntLLROutputS2xD(245)(2);
  VNStageIntLLRInputS2xD(200)(4) <= CNStageIntLLROutputS2xD(245)(3);
  VNStageIntLLRInputS2xD(284)(4) <= CNStageIntLLROutputS2xD(245)(4);
  VNStageIntLLRInputS2xD(340)(4) <= CNStageIntLLROutputS2xD(245)(5);
  VNStageIntLLRInputS2xD(57)(3) <= CNStageIntLLROutputS2xD(246)(0);
  VNStageIntLLRInputS2xD(70)(4) <= CNStageIntLLROutputS2xD(246)(1);
  VNStageIntLLRInputS2xD(154)(3) <= CNStageIntLLROutputS2xD(246)(2);
  VNStageIntLLRInputS2xD(210)(4) <= CNStageIntLLROutputS2xD(246)(3);
  VNStageIntLLRInputS2xD(312)(3) <= CNStageIntLLROutputS2xD(246)(4);
  VNStageIntLLRInputS2xD(378)(3) <= CNStageIntLLROutputS2xD(246)(5);
  VNStageIntLLRInputS2xD(56)(4) <= CNStageIntLLROutputS2xD(247)(0);
  VNStageIntLLRInputS2xD(89)(4) <= CNStageIntLLROutputS2xD(247)(1);
  VNStageIntLLRInputS2xD(145)(4) <= CNStageIntLLROutputS2xD(247)(2);
  VNStageIntLLRInputS2xD(247)(4) <= CNStageIntLLROutputS2xD(247)(3);
  VNStageIntLLRInputS2xD(313)(2) <= CNStageIntLLROutputS2xD(247)(4);
  VNStageIntLLRInputS2xD(339)(4) <= CNStageIntLLROutputS2xD(247)(5);
  VNStageIntLLRInputS2xD(55)(4) <= CNStageIntLLROutputS2xD(248)(0);
  VNStageIntLLRInputS2xD(80)(4) <= CNStageIntLLROutputS2xD(248)(1);
  VNStageIntLLRInputS2xD(182)(4) <= CNStageIntLLROutputS2xD(248)(2);
  VNStageIntLLRInputS2xD(248)(4) <= CNStageIntLLROutputS2xD(248)(3);
  VNStageIntLLRInputS2xD(274)(3) <= CNStageIntLLROutputS2xD(248)(4);
  VNStageIntLLRInputS2xD(360)(4) <= CNStageIntLLROutputS2xD(248)(5);
  VNStageIntLLRInputS2xD(53)(3) <= CNStageIntLLROutputS2xD(249)(0);
  VNStageIntLLRInputS2xD(118)(3) <= CNStageIntLLROutputS2xD(249)(1);
  VNStageIntLLRInputS2xD(144)(4) <= CNStageIntLLROutputS2xD(249)(2);
  VNStageIntLLRInputS2xD(230)(3) <= CNStageIntLLROutputS2xD(249)(3);
  VNStageIntLLRInputS2xD(291)(4) <= CNStageIntLLROutputS2xD(249)(4);
  VNStageIntLLRInputS2xD(371)(3) <= CNStageIntLLROutputS2xD(249)(5);
  VNStageIntLLRInputS2xD(51)(3) <= CNStageIntLLROutputS2xD(250)(0);
  VNStageIntLLRInputS2xD(100)(4) <= CNStageIntLLROutputS2xD(250)(1);
  VNStageIntLLRInputS2xD(161)(4) <= CNStageIntLLROutputS2xD(250)(2);
  VNStageIntLLRInputS2xD(241)(3) <= CNStageIntLLROutputS2xD(250)(3);
  VNStageIntLLRInputS2xD(269)(3) <= CNStageIntLLROutputS2xD(250)(4);
  VNStageIntLLRInputS2xD(373)(2) <= CNStageIntLLROutputS2xD(250)(5);
  VNStageIntLLRInputS2xD(50)(4) <= CNStageIntLLROutputS2xD(251)(0);
  VNStageIntLLRInputS2xD(96)(4) <= CNStageIntLLROutputS2xD(251)(1);
  VNStageIntLLRInputS2xD(176)(4) <= CNStageIntLLROutputS2xD(251)(2);
  VNStageIntLLRInputS2xD(204)(4) <= CNStageIntLLROutputS2xD(251)(3);
  VNStageIntLLRInputS2xD(308)(2) <= CNStageIntLLROutputS2xD(251)(4);
  VNStageIntLLRInputS2xD(342)(3) <= CNStageIntLLROutputS2xD(251)(5);
  VNStageIntLLRInputS2xD(49)(4) <= CNStageIntLLROutputS2xD(252)(0);
  VNStageIntLLRInputS2xD(111)(4) <= CNStageIntLLROutputS2xD(252)(1);
  VNStageIntLLRInputS2xD(139)(4) <= CNStageIntLLROutputS2xD(252)(2);
  VNStageIntLLRInputS2xD(243)(4) <= CNStageIntLLROutputS2xD(252)(3);
  VNStageIntLLRInputS2xD(277)(4) <= CNStageIntLLROutputS2xD(252)(4);
  VNStageIntLLRInputS2xD(358)(3) <= CNStageIntLLROutputS2xD(252)(5);
  VNStageIntLLRInputS2xD(47)(2) <= CNStageIntLLROutputS2xD(253)(0);
  VNStageIntLLRInputS2xD(113)(4) <= CNStageIntLLROutputS2xD(253)(1);
  VNStageIntLLRInputS2xD(147)(4) <= CNStageIntLLROutputS2xD(253)(2);
  VNStageIntLLRInputS2xD(228)(4) <= CNStageIntLLROutputS2xD(253)(3);
  VNStageIntLLRInputS2xD(263)(4) <= CNStageIntLLROutputS2xD(253)(4);
  VNStageIntLLRInputS2xD(337)(4) <= CNStageIntLLROutputS2xD(253)(5);
  VNStageIntLLRInputS2xD(46)(4) <= CNStageIntLLROutputS2xD(254)(0);
  VNStageIntLLRInputS2xD(82)(4) <= CNStageIntLLROutputS2xD(254)(1);
  VNStageIntLLRInputS2xD(163)(3) <= CNStageIntLLROutputS2xD(254)(2);
  VNStageIntLLRInputS2xD(198)(4) <= CNStageIntLLROutputS2xD(254)(3);
  VNStageIntLLRInputS2xD(272)(4) <= CNStageIntLLROutputS2xD(254)(4);
  VNStageIntLLRInputS2xD(350)(4) <= CNStageIntLLROutputS2xD(254)(5);
  VNStageIntLLRInputS2xD(45)(4) <= CNStageIntLLROutputS2xD(255)(0);
  VNStageIntLLRInputS2xD(98)(3) <= CNStageIntLLROutputS2xD(255)(1);
  VNStageIntLLRInputS2xD(133)(2) <= CNStageIntLLROutputS2xD(255)(2);
  VNStageIntLLRInputS2xD(207)(3) <= CNStageIntLLROutputS2xD(255)(3);
  VNStageIntLLRInputS2xD(285)(4) <= CNStageIntLLROutputS2xD(255)(4);
  VNStageIntLLRInputS2xD(329)(4) <= CNStageIntLLROutputS2xD(255)(5);
  VNStageIntLLRInputS2xD(44)(4) <= CNStageIntLLROutputS2xD(256)(0);
  VNStageIntLLRInputS2xD(68)(3) <= CNStageIntLLROutputS2xD(256)(1);
  VNStageIntLLRInputS2xD(142)(3) <= CNStageIntLLROutputS2xD(256)(2);
  VNStageIntLLRInputS2xD(220)(4) <= CNStageIntLLROutputS2xD(256)(3);
  VNStageIntLLRInputS2xD(264)(4) <= CNStageIntLLROutputS2xD(256)(4);
  VNStageIntLLRInputS2xD(357)(4) <= CNStageIntLLROutputS2xD(256)(5);
  VNStageIntLLRInputS2xD(43)(3) <= CNStageIntLLROutputS2xD(257)(0);
  VNStageIntLLRInputS2xD(77)(2) <= CNStageIntLLROutputS2xD(257)(1);
  VNStageIntLLRInputS2xD(155)(4) <= CNStageIntLLROutputS2xD(257)(2);
  VNStageIntLLRInputS2xD(199)(4) <= CNStageIntLLROutputS2xD(257)(3);
  VNStageIntLLRInputS2xD(292)(4) <= CNStageIntLLROutputS2xD(257)(4);
  VNStageIntLLRInputS2xD(359)(4) <= CNStageIntLLROutputS2xD(257)(5);
  VNStageIntLLRInputS2xD(42)(4) <= CNStageIntLLROutputS2xD(258)(0);
  VNStageIntLLRInputS2xD(90)(4) <= CNStageIntLLROutputS2xD(258)(1);
  VNStageIntLLRInputS2xD(134)(3) <= CNStageIntLLROutputS2xD(258)(2);
  VNStageIntLLRInputS2xD(227)(4) <= CNStageIntLLROutputS2xD(258)(3);
  VNStageIntLLRInputS2xD(294)(4) <= CNStageIntLLROutputS2xD(258)(4);
  VNStageIntLLRInputS2xD(341)(4) <= CNStageIntLLROutputS2xD(258)(5);
  VNStageIntLLRInputS2xD(41)(4) <= CNStageIntLLROutputS2xD(259)(0);
  VNStageIntLLRInputS2xD(69)(4) <= CNStageIntLLROutputS2xD(259)(1);
  VNStageIntLLRInputS2xD(162)(4) <= CNStageIntLLROutputS2xD(259)(2);
  VNStageIntLLRInputS2xD(229)(3) <= CNStageIntLLROutputS2xD(259)(3);
  VNStageIntLLRInputS2xD(276)(4) <= CNStageIntLLROutputS2xD(259)(4);
  VNStageIntLLRInputS2xD(348)(4) <= CNStageIntLLROutputS2xD(259)(5);
  VNStageIntLLRInputS2xD(40)(3) <= CNStageIntLLROutputS2xD(260)(0);
  VNStageIntLLRInputS2xD(97)(4) <= CNStageIntLLROutputS2xD(260)(1);
  VNStageIntLLRInputS2xD(164)(4) <= CNStageIntLLROutputS2xD(260)(2);
  VNStageIntLLRInputS2xD(211)(4) <= CNStageIntLLROutputS2xD(260)(3);
  VNStageIntLLRInputS2xD(283)(4) <= CNStageIntLLROutputS2xD(260)(4);
  VNStageIntLLRInputS2xD(375)(3) <= CNStageIntLLROutputS2xD(260)(5);
  VNStageIntLLRInputS2xD(39)(4) <= CNStageIntLLROutputS2xD(261)(0);
  VNStageIntLLRInputS2xD(99)(4) <= CNStageIntLLROutputS2xD(261)(1);
  VNStageIntLLRInputS2xD(146)(3) <= CNStageIntLLROutputS2xD(261)(2);
  VNStageIntLLRInputS2xD(218)(4) <= CNStageIntLLROutputS2xD(261)(3);
  VNStageIntLLRInputS2xD(310)(3) <= CNStageIntLLROutputS2xD(261)(4);
  VNStageIntLLRInputS2xD(363)(3) <= CNStageIntLLROutputS2xD(261)(5);
  VNStageIntLLRInputS2xD(38)(4) <= CNStageIntLLROutputS2xD(262)(0);
  VNStageIntLLRInputS2xD(81)(3) <= CNStageIntLLROutputS2xD(262)(1);
  VNStageIntLLRInputS2xD(153)(4) <= CNStageIntLLROutputS2xD(262)(2);
  VNStageIntLLRInputS2xD(245)(4) <= CNStageIntLLROutputS2xD(262)(3);
  VNStageIntLLRInputS2xD(298)(4) <= CNStageIntLLROutputS2xD(262)(4);
  VNStageIntLLRInputS2xD(369)(3) <= CNStageIntLLROutputS2xD(262)(5);
  VNStageIntLLRInputS2xD(37)(4) <= CNStageIntLLROutputS2xD(263)(0);
  VNStageIntLLRInputS2xD(88)(4) <= CNStageIntLLROutputS2xD(263)(1);
  VNStageIntLLRInputS2xD(180)(2) <= CNStageIntLLROutputS2xD(263)(2);
  VNStageIntLLRInputS2xD(233)(3) <= CNStageIntLLROutputS2xD(263)(3);
  VNStageIntLLRInputS2xD(304)(4) <= CNStageIntLLROutputS2xD(263)(4);
  VNStageIntLLRInputS2xD(364)(4) <= CNStageIntLLROutputS2xD(263)(5);
  VNStageIntLLRInputS2xD(36)(3) <= CNStageIntLLROutputS2xD(264)(0);
  VNStageIntLLRInputS2xD(115)(4) <= CNStageIntLLROutputS2xD(264)(1);
  VNStageIntLLRInputS2xD(168)(3) <= CNStageIntLLROutputS2xD(264)(2);
  VNStageIntLLRInputS2xD(239)(4) <= CNStageIntLLROutputS2xD(264)(3);
  VNStageIntLLRInputS2xD(299)(3) <= CNStageIntLLROutputS2xD(264)(4);
  VNStageIntLLRInputS2xD(374)(4) <= CNStageIntLLROutputS2xD(264)(5);
  VNStageIntLLRInputS2xD(35)(4) <= CNStageIntLLROutputS2xD(265)(0);
  VNStageIntLLRInputS2xD(103)(4) <= CNStageIntLLROutputS2xD(265)(1);
  VNStageIntLLRInputS2xD(174)(3) <= CNStageIntLLROutputS2xD(265)(2);
  VNStageIntLLRInputS2xD(234)(4) <= CNStageIntLLROutputS2xD(265)(3);
  VNStageIntLLRInputS2xD(309)(4) <= CNStageIntLLROutputS2xD(265)(4);
  VNStageIntLLRInputS2xD(333)(3) <= CNStageIntLLROutputS2xD(265)(5);
  VNStageIntLLRInputS2xD(34)(4) <= CNStageIntLLROutputS2xD(266)(0);
  VNStageIntLLRInputS2xD(109)(4) <= CNStageIntLLROutputS2xD(266)(1);
  VNStageIntLLRInputS2xD(169)(4) <= CNStageIntLLROutputS2xD(266)(2);
  VNStageIntLLRInputS2xD(244)(1) <= CNStageIntLLROutputS2xD(266)(3);
  VNStageIntLLRInputS2xD(268)(4) <= CNStageIntLLROutputS2xD(266)(4);
  VNStageIntLLRInputS2xD(351)(3) <= CNStageIntLLROutputS2xD(266)(5);
  VNStageIntLLRInputS2xD(33)(4) <= CNStageIntLLROutputS2xD(267)(0);
  VNStageIntLLRInputS2xD(104)(4) <= CNStageIntLLROutputS2xD(267)(1);
  VNStageIntLLRInputS2xD(179)(4) <= CNStageIntLLROutputS2xD(267)(2);
  VNStageIntLLRInputS2xD(203)(4) <= CNStageIntLLROutputS2xD(267)(3);
  VNStageIntLLRInputS2xD(286)(4) <= CNStageIntLLROutputS2xD(267)(4);
  VNStageIntLLRInputS2xD(336)(3) <= CNStageIntLLROutputS2xD(267)(5);
  VNStageIntLLRInputS2xD(32)(3) <= CNStageIntLLROutputS2xD(268)(0);
  VNStageIntLLRInputS2xD(114)(4) <= CNStageIntLLROutputS2xD(268)(1);
  VNStageIntLLRInputS2xD(138)(4) <= CNStageIntLLROutputS2xD(268)(2);
  VNStageIntLLRInputS2xD(221)(4) <= CNStageIntLLROutputS2xD(268)(3);
  VNStageIntLLRInputS2xD(271)(3) <= CNStageIntLLROutputS2xD(268)(4);
  VNStageIntLLRInputS2xD(323)(3) <= CNStageIntLLROutputS2xD(268)(5);
  VNStageIntLLRInputS2xD(30)(4) <= CNStageIntLLROutputS2xD(269)(0);
  VNStageIntLLRInputS2xD(91)(4) <= CNStageIntLLROutputS2xD(269)(1);
  VNStageIntLLRInputS2xD(141)(2) <= CNStageIntLLROutputS2xD(269)(2);
  VNStageIntLLRInputS2xD(193)(3) <= CNStageIntLLROutputS2xD(269)(3);
  VNStageIntLLRInputS2xD(289)(4) <= CNStageIntLLROutputS2xD(269)(4);
  VNStageIntLLRInputS2xD(366)(4) <= CNStageIntLLROutputS2xD(269)(5);
  VNStageIntLLRInputS2xD(29)(3) <= CNStageIntLLROutputS2xD(270)(0);
  VNStageIntLLRInputS2xD(76)(4) <= CNStageIntLLROutputS2xD(270)(1);
  VNStageIntLLRInputS2xD(191)(4) <= CNStageIntLLROutputS2xD(270)(2);
  VNStageIntLLRInputS2xD(224)(4) <= CNStageIntLLROutputS2xD(270)(3);
  VNStageIntLLRInputS2xD(301)(4) <= CNStageIntLLROutputS2xD(270)(4);
  VNStageIntLLRInputS2xD(380)(3) <= CNStageIntLLROutputS2xD(270)(5);
  VNStageIntLLRInputS2xD(28)(4) <= CNStageIntLLROutputS2xD(271)(0);
  VNStageIntLLRInputS2xD(126)(3) <= CNStageIntLLROutputS2xD(271)(1);
  VNStageIntLLRInputS2xD(159)(3) <= CNStageIntLLROutputS2xD(271)(2);
  VNStageIntLLRInputS2xD(236)(4) <= CNStageIntLLROutputS2xD(271)(3);
  VNStageIntLLRInputS2xD(315)(3) <= CNStageIntLLROutputS2xD(271)(4);
  VNStageIntLLRInputS2xD(361)(4) <= CNStageIntLLROutputS2xD(271)(5);
  VNStageIntLLRInputS2xD(26)(4) <= CNStageIntLLROutputS2xD(272)(0);
  VNStageIntLLRInputS2xD(106)(3) <= CNStageIntLLROutputS2xD(272)(1);
  VNStageIntLLRInputS2xD(185)(1) <= CNStageIntLLROutputS2xD(272)(2);
  VNStageIntLLRInputS2xD(231)(3) <= CNStageIntLLROutputS2xD(272)(3);
  VNStageIntLLRInputS2xD(273)(3) <= CNStageIntLLROutputS2xD(272)(4);
  VNStageIntLLRInputS2xD(327)(4) <= CNStageIntLLROutputS2xD(272)(5);
  VNStageIntLLRInputS2xD(24)(4) <= CNStageIntLLROutputS2xD(273)(0);
  VNStageIntLLRInputS2xD(101)(4) <= CNStageIntLLROutputS2xD(273)(1);
  VNStageIntLLRInputS2xD(143)(4) <= CNStageIntLLROutputS2xD(273)(2);
  VNStageIntLLRInputS2xD(197)(4) <= CNStageIntLLROutputS2xD(273)(3);
  VNStageIntLLRInputS2xD(266)(3) <= CNStageIntLLROutputS2xD(273)(4);
  VNStageIntLLRInputS2xD(324)(4) <= CNStageIntLLROutputS2xD(273)(5);
  VNStageIntLLRInputS2xD(23)(4) <= CNStageIntLLROutputS2xD(274)(0);
  VNStageIntLLRInputS2xD(78)(4) <= CNStageIntLLROutputS2xD(274)(1);
  VNStageIntLLRInputS2xD(132)(3) <= CNStageIntLLROutputS2xD(274)(2);
  VNStageIntLLRInputS2xD(201)(4) <= CNStageIntLLROutputS2xD(274)(3);
  VNStageIntLLRInputS2xD(259)(2) <= CNStageIntLLROutputS2xD(274)(4);
  VNStageIntLLRInputS2xD(335)(4) <= CNStageIntLLROutputS2xD(274)(5);
  VNStageIntLLRInputS2xD(22)(4) <= CNStageIntLLROutputS2xD(275)(0);
  VNStageIntLLRInputS2xD(67)(1) <= CNStageIntLLROutputS2xD(275)(1);
  VNStageIntLLRInputS2xD(136)(4) <= CNStageIntLLROutputS2xD(275)(2);
  VNStageIntLLRInputS2xD(194)(4) <= CNStageIntLLROutputS2xD(275)(3);
  VNStageIntLLRInputS2xD(270)(4) <= CNStageIntLLROutputS2xD(275)(4);
  VNStageIntLLRInputS2xD(370)(3) <= CNStageIntLLROutputS2xD(275)(5);
  VNStageIntLLRInputS2xD(21)(4) <= CNStageIntLLROutputS2xD(276)(0);
  VNStageIntLLRInputS2xD(71)(3) <= CNStageIntLLROutputS2xD(276)(1);
  VNStageIntLLRInputS2xD(129)(4) <= CNStageIntLLROutputS2xD(276)(2);
  VNStageIntLLRInputS2xD(205)(1) <= CNStageIntLLROutputS2xD(276)(3);
  VNStageIntLLRInputS2xD(305)(4) <= CNStageIntLLROutputS2xD(276)(4);
  VNStageIntLLRInputS2xD(362)(4) <= CNStageIntLLROutputS2xD(276)(5);
  VNStageIntLLRInputS2xD(20)(2) <= CNStageIntLLROutputS2xD(277)(0);
  VNStageIntLLRInputS2xD(127)(4) <= CNStageIntLLROutputS2xD(277)(1);
  VNStageIntLLRInputS2xD(140)(4) <= CNStageIntLLROutputS2xD(277)(2);
  VNStageIntLLRInputS2xD(240)(4) <= CNStageIntLLROutputS2xD(277)(3);
  VNStageIntLLRInputS2xD(297)(4) <= CNStageIntLLROutputS2xD(277)(4);
  VNStageIntLLRInputS2xD(379)(2) <= CNStageIntLLROutputS2xD(277)(5);
  VNStageIntLLRInputS2xD(19)(3) <= CNStageIntLLROutputS2xD(278)(0);
  VNStageIntLLRInputS2xD(75)(4) <= CNStageIntLLROutputS2xD(278)(1);
  VNStageIntLLRInputS2xD(175)(4) <= CNStageIntLLROutputS2xD(278)(2);
  VNStageIntLLRInputS2xD(232)(3) <= CNStageIntLLROutputS2xD(278)(3);
  VNStageIntLLRInputS2xD(314)(1) <= CNStageIntLLROutputS2xD(278)(4);
  VNStageIntLLRInputS2xD(376)(3) <= CNStageIntLLROutputS2xD(278)(5);
  VNStageIntLLRInputS2xD(0)(4) <= CNStageIntLLROutputS2xD(279)(0);
  VNStageIntLLRInputS2xD(123)(3) <= CNStageIntLLROutputS2xD(279)(1);
  VNStageIntLLRInputS2xD(188)(2) <= CNStageIntLLROutputS2xD(279)(2);
  VNStageIntLLRInputS2xD(253)(3) <= CNStageIntLLROutputS2xD(279)(3);
  VNStageIntLLRInputS2xD(318)(2) <= CNStageIntLLROutputS2xD(279)(4);
  VNStageIntLLRInputS2xD(383)(4) <= CNStageIntLLROutputS2xD(279)(5);
  VNStageIntLLRInputS2xD(35)(5) <= CNStageIntLLROutputS2xD(280)(0);
  VNStageIntLLRInputS2xD(91)(5) <= CNStageIntLLROutputS2xD(280)(1);
  VNStageIntLLRInputS2xD(191)(5) <= CNStageIntLLROutputS2xD(280)(2);
  VNStageIntLLRInputS2xD(248)(5) <= CNStageIntLLROutputS2xD(280)(3);
  VNStageIntLLRInputS2xD(267)(5) <= CNStageIntLLROutputS2xD(280)(4);
  VNStageIntLLRInputS2xD(329)(5) <= CNStageIntLLROutputS2xD(280)(5);
  VNStageIntLLRInputS2xD(34)(5) <= CNStageIntLLROutputS2xD(281)(0);
  VNStageIntLLRInputS2xD(126)(4) <= CNStageIntLLROutputS2xD(281)(1);
  VNStageIntLLRInputS2xD(183)(3) <= CNStageIntLLROutputS2xD(281)(2);
  VNStageIntLLRInputS2xD(202)(4) <= CNStageIntLLROutputS2xD(281)(3);
  VNStageIntLLRInputS2xD(264)(5) <= CNStageIntLLROutputS2xD(281)(4);
  VNStageIntLLRInputS2xD(363)(4) <= CNStageIntLLROutputS2xD(281)(5);
  VNStageIntLLRInputS2xD(33)(5) <= CNStageIntLLROutputS2xD(282)(0);
  VNStageIntLLRInputS2xD(118)(4) <= CNStageIntLLROutputS2xD(282)(1);
  VNStageIntLLRInputS2xD(137)(5) <= CNStageIntLLROutputS2xD(282)(2);
  VNStageIntLLRInputS2xD(199)(5) <= CNStageIntLLROutputS2xD(282)(3);
  VNStageIntLLRInputS2xD(298)(5) <= CNStageIntLLROutputS2xD(282)(4);
  VNStageIntLLRInputS2xD(383)(5) <= CNStageIntLLROutputS2xD(282)(5);
  VNStageIntLLRInputS2xD(31)(3) <= CNStageIntLLROutputS2xD(283)(0);
  VNStageIntLLRInputS2xD(69)(5) <= CNStageIntLLROutputS2xD(283)(1);
  VNStageIntLLRInputS2xD(168)(4) <= CNStageIntLLROutputS2xD(283)(2);
  VNStageIntLLRInputS2xD(253)(4) <= CNStageIntLLROutputS2xD(283)(3);
  VNStageIntLLRInputS2xD(304)(5) <= CNStageIntLLROutputS2xD(283)(4);
  VNStageIntLLRInputS2xD(359)(5) <= CNStageIntLLROutputS2xD(283)(5);
  VNStageIntLLRInputS2xD(30)(5) <= CNStageIntLLROutputS2xD(284)(0);
  VNStageIntLLRInputS2xD(103)(5) <= CNStageIntLLROutputS2xD(284)(1);
  VNStageIntLLRInputS2xD(188)(3) <= CNStageIntLLROutputS2xD(284)(2);
  VNStageIntLLRInputS2xD(239)(5) <= CNStageIntLLROutputS2xD(284)(3);
  VNStageIntLLRInputS2xD(294)(5) <= CNStageIntLLROutputS2xD(284)(4);
  VNStageIntLLRInputS2xD(325)(5) <= CNStageIntLLROutputS2xD(284)(5);
  VNStageIntLLRInputS2xD(27)(4) <= CNStageIntLLROutputS2xD(285)(0);
  VNStageIntLLRInputS2xD(99)(5) <= CNStageIntLLROutputS2xD(285)(1);
  VNStageIntLLRInputS2xD(130)(5) <= CNStageIntLLROutputS2xD(285)(2);
  VNStageIntLLRInputS2xD(241)(4) <= CNStageIntLLROutputS2xD(285)(3);
  VNStageIntLLRInputS2xD(273)(4) <= CNStageIntLLROutputS2xD(285)(4);
  VNStageIntLLRInputS2xD(361)(5) <= CNStageIntLLROutputS2xD(285)(5);
  VNStageIntLLRInputS2xD(26)(5) <= CNStageIntLLROutputS2xD(286)(0);
  VNStageIntLLRInputS2xD(65)(4) <= CNStageIntLLROutputS2xD(286)(1);
  VNStageIntLLRInputS2xD(176)(5) <= CNStageIntLLROutputS2xD(286)(2);
  VNStageIntLLRInputS2xD(208)(4) <= CNStageIntLLROutputS2xD(286)(3);
  VNStageIntLLRInputS2xD(296)(4) <= CNStageIntLLROutputS2xD(286)(4);
  VNStageIntLLRInputS2xD(334)(3) <= CNStageIntLLROutputS2xD(286)(5);
  VNStageIntLLRInputS2xD(25)(4) <= CNStageIntLLROutputS2xD(287)(0);
  VNStageIntLLRInputS2xD(111)(5) <= CNStageIntLLROutputS2xD(287)(1);
  VNStageIntLLRInputS2xD(143)(5) <= CNStageIntLLROutputS2xD(287)(2);
  VNStageIntLLRInputS2xD(231)(4) <= CNStageIntLLROutputS2xD(287)(3);
  VNStageIntLLRInputS2xD(269)(4) <= CNStageIntLLROutputS2xD(287)(4);
  VNStageIntLLRInputS2xD(381)(4) <= CNStageIntLLROutputS2xD(287)(5);
  VNStageIntLLRInputS2xD(24)(5) <= CNStageIntLLROutputS2xD(288)(0);
  VNStageIntLLRInputS2xD(78)(5) <= CNStageIntLLROutputS2xD(288)(1);
  VNStageIntLLRInputS2xD(166)(4) <= CNStageIntLLROutputS2xD(288)(2);
  VNStageIntLLRInputS2xD(204)(5) <= CNStageIntLLROutputS2xD(288)(3);
  VNStageIntLLRInputS2xD(316)(3) <= CNStageIntLLROutputS2xD(288)(4);
  VNStageIntLLRInputS2xD(321)(5) <= CNStageIntLLROutputS2xD(288)(5);
  VNStageIntLLRInputS2xD(23)(5) <= CNStageIntLLROutputS2xD(289)(0);
  VNStageIntLLRInputS2xD(101)(5) <= CNStageIntLLROutputS2xD(289)(1);
  VNStageIntLLRInputS2xD(139)(5) <= CNStageIntLLROutputS2xD(289)(2);
  VNStageIntLLRInputS2xD(251)(3) <= CNStageIntLLROutputS2xD(289)(3);
  VNStageIntLLRInputS2xD(319)(5) <= CNStageIntLLROutputS2xD(289)(4);
  VNStageIntLLRInputS2xD(362)(5) <= CNStageIntLLROutputS2xD(289)(5);
  VNStageIntLLRInputS2xD(22)(5) <= CNStageIntLLROutputS2xD(290)(0);
  VNStageIntLLRInputS2xD(74)(4) <= CNStageIntLLROutputS2xD(290)(1);
  VNStageIntLLRInputS2xD(186)(4) <= CNStageIntLLROutputS2xD(290)(2);
  VNStageIntLLRInputS2xD(254)(3) <= CNStageIntLLROutputS2xD(290)(3);
  VNStageIntLLRInputS2xD(297)(5) <= CNStageIntLLROutputS2xD(290)(4);
  VNStageIntLLRInputS2xD(337)(5) <= CNStageIntLLROutputS2xD(290)(5);
  VNStageIntLLRInputS2xD(21)(5) <= CNStageIntLLROutputS2xD(291)(0);
  VNStageIntLLRInputS2xD(121)(4) <= CNStageIntLLROutputS2xD(291)(1);
  VNStageIntLLRInputS2xD(189)(4) <= CNStageIntLLROutputS2xD(291)(2);
  VNStageIntLLRInputS2xD(232)(4) <= CNStageIntLLROutputS2xD(291)(3);
  VNStageIntLLRInputS2xD(272)(5) <= CNStageIntLLROutputS2xD(291)(4);
  VNStageIntLLRInputS2xD(335)(5) <= CNStageIntLLROutputS2xD(291)(5);
  VNStageIntLLRInputS2xD(20)(3) <= CNStageIntLLROutputS2xD(292)(0);
  VNStageIntLLRInputS2xD(124)(3) <= CNStageIntLLROutputS2xD(292)(1);
  VNStageIntLLRInputS2xD(167)(5) <= CNStageIntLLROutputS2xD(292)(2);
  VNStageIntLLRInputS2xD(207)(4) <= CNStageIntLLROutputS2xD(292)(3);
  VNStageIntLLRInputS2xD(270)(5) <= CNStageIntLLROutputS2xD(292)(4);
  VNStageIntLLRInputS2xD(360)(5) <= CNStageIntLLROutputS2xD(292)(5);
  VNStageIntLLRInputS2xD(18)(5) <= CNStageIntLLROutputS2xD(293)(0);
  VNStageIntLLRInputS2xD(77)(3) <= CNStageIntLLROutputS2xD(293)(1);
  VNStageIntLLRInputS2xD(140)(5) <= CNStageIntLLROutputS2xD(293)(2);
  VNStageIntLLRInputS2xD(230)(4) <= CNStageIntLLROutputS2xD(293)(3);
  VNStageIntLLRInputS2xD(303)(5) <= CNStageIntLLROutputS2xD(293)(4);
  VNStageIntLLRInputS2xD(348)(5) <= CNStageIntLLROutputS2xD(293)(5);
  VNStageIntLLRInputS2xD(17)(5) <= CNStageIntLLROutputS2xD(294)(0);
  VNStageIntLLRInputS2xD(75)(5) <= CNStageIntLLROutputS2xD(294)(1);
  VNStageIntLLRInputS2xD(165)(4) <= CNStageIntLLROutputS2xD(294)(2);
  VNStageIntLLRInputS2xD(238)(5) <= CNStageIntLLROutputS2xD(294)(3);
  VNStageIntLLRInputS2xD(283)(5) <= CNStageIntLLROutputS2xD(294)(4);
  VNStageIntLLRInputS2xD(342)(4) <= CNStageIntLLROutputS2xD(294)(5);
  VNStageIntLLRInputS2xD(16)(4) <= CNStageIntLLROutputS2xD(295)(0);
  VNStageIntLLRInputS2xD(100)(5) <= CNStageIntLLROutputS2xD(295)(1);
  VNStageIntLLRInputS2xD(173)(5) <= CNStageIntLLROutputS2xD(295)(2);
  VNStageIntLLRInputS2xD(218)(5) <= CNStageIntLLROutputS2xD(295)(3);
  VNStageIntLLRInputS2xD(277)(5) <= CNStageIntLLROutputS2xD(295)(4);
  VNStageIntLLRInputS2xD(320)(3) <= CNStageIntLLROutputS2xD(295)(5);
  VNStageIntLLRInputS2xD(15)(5) <= CNStageIntLLROutputS2xD(296)(0);
  VNStageIntLLRInputS2xD(108)(5) <= CNStageIntLLROutputS2xD(296)(1);
  VNStageIntLLRInputS2xD(153)(5) <= CNStageIntLLROutputS2xD(296)(2);
  VNStageIntLLRInputS2xD(212)(4) <= CNStageIntLLROutputS2xD(296)(3);
  VNStageIntLLRInputS2xD(256)(4) <= CNStageIntLLROutputS2xD(296)(4);
  VNStageIntLLRInputS2xD(341)(5) <= CNStageIntLLROutputS2xD(296)(5);
  VNStageIntLLRInputS2xD(14)(5) <= CNStageIntLLROutputS2xD(297)(0);
  VNStageIntLLRInputS2xD(88)(5) <= CNStageIntLLROutputS2xD(297)(1);
  VNStageIntLLRInputS2xD(147)(5) <= CNStageIntLLROutputS2xD(297)(2);
  VNStageIntLLRInputS2xD(192)(5) <= CNStageIntLLROutputS2xD(297)(3);
  VNStageIntLLRInputS2xD(276)(5) <= CNStageIntLLROutputS2xD(297)(4);
  VNStageIntLLRInputS2xD(346)(5) <= CNStageIntLLROutputS2xD(297)(5);
  VNStageIntLLRInputS2xD(13)(4) <= CNStageIntLLROutputS2xD(298)(0);
  VNStageIntLLRInputS2xD(82)(5) <= CNStageIntLLROutputS2xD(298)(1);
  VNStageIntLLRInputS2xD(128)(5) <= CNStageIntLLROutputS2xD(298)(2);
  VNStageIntLLRInputS2xD(211)(5) <= CNStageIntLLROutputS2xD(298)(3);
  VNStageIntLLRInputS2xD(281)(5) <= CNStageIntLLROutputS2xD(298)(4);
  VNStageIntLLRInputS2xD(365)(5) <= CNStageIntLLROutputS2xD(298)(5);
  VNStageIntLLRInputS2xD(12)(5) <= CNStageIntLLROutputS2xD(299)(0);
  VNStageIntLLRInputS2xD(64)(4) <= CNStageIntLLROutputS2xD(299)(1);
  VNStageIntLLRInputS2xD(146)(4) <= CNStageIntLLROutputS2xD(299)(2);
  VNStageIntLLRInputS2xD(216)(5) <= CNStageIntLLROutputS2xD(299)(3);
  VNStageIntLLRInputS2xD(300)(4) <= CNStageIntLLROutputS2xD(299)(4);
  VNStageIntLLRInputS2xD(356)(4) <= CNStageIntLLROutputS2xD(299)(5);
  VNStageIntLLRInputS2xD(9)(5) <= CNStageIntLLROutputS2xD(300)(0);
  VNStageIntLLRInputS2xD(105)(4) <= CNStageIntLLROutputS2xD(300)(1);
  VNStageIntLLRInputS2xD(161)(5) <= CNStageIntLLROutputS2xD(300)(2);
  VNStageIntLLRInputS2xD(200)(5) <= CNStageIntLLROutputS2xD(300)(3);
  VNStageIntLLRInputS2xD(266)(4) <= CNStageIntLLROutputS2xD(300)(4);
  VNStageIntLLRInputS2xD(355)(5) <= CNStageIntLLROutputS2xD(300)(5);
  VNStageIntLLRInputS2xD(7)(5) <= CNStageIntLLROutputS2xD(301)(0);
  VNStageIntLLRInputS2xD(70)(5) <= CNStageIntLLROutputS2xD(301)(1);
  VNStageIntLLRInputS2xD(136)(5) <= CNStageIntLLROutputS2xD(301)(2);
  VNStageIntLLRInputS2xD(225)(5) <= CNStageIntLLROutputS2xD(301)(3);
  VNStageIntLLRInputS2xD(311)(4) <= CNStageIntLLROutputS2xD(301)(4);
  VNStageIntLLRInputS2xD(372)(4) <= CNStageIntLLROutputS2xD(301)(5);
  VNStageIntLLRInputS2xD(6)(5) <= CNStageIntLLROutputS2xD(302)(0);
  VNStageIntLLRInputS2xD(71)(4) <= CNStageIntLLROutputS2xD(302)(1);
  VNStageIntLLRInputS2xD(160)(5) <= CNStageIntLLROutputS2xD(302)(2);
  VNStageIntLLRInputS2xD(246)(5) <= CNStageIntLLROutputS2xD(302)(3);
  VNStageIntLLRInputS2xD(307)(5) <= CNStageIntLLROutputS2xD(302)(4);
  VNStageIntLLRInputS2xD(324)(5) <= CNStageIntLLROutputS2xD(302)(5);
  VNStageIntLLRInputS2xD(5)(5) <= CNStageIntLLROutputS2xD(303)(0);
  VNStageIntLLRInputS2xD(95)(5) <= CNStageIntLLROutputS2xD(303)(1);
  VNStageIntLLRInputS2xD(181)(5) <= CNStageIntLLROutputS2xD(303)(2);
  VNStageIntLLRInputS2xD(242)(5) <= CNStageIntLLROutputS2xD(303)(3);
  VNStageIntLLRInputS2xD(259)(3) <= CNStageIntLLROutputS2xD(303)(4);
  VNStageIntLLRInputS2xD(350)(5) <= CNStageIntLLROutputS2xD(303)(5);
  VNStageIntLLRInputS2xD(4)(4) <= CNStageIntLLROutputS2xD(304)(0);
  VNStageIntLLRInputS2xD(116)(4) <= CNStageIntLLROutputS2xD(304)(1);
  VNStageIntLLRInputS2xD(177)(5) <= CNStageIntLLROutputS2xD(304)(2);
  VNStageIntLLRInputS2xD(194)(5) <= CNStageIntLLROutputS2xD(304)(3);
  VNStageIntLLRInputS2xD(285)(5) <= CNStageIntLLROutputS2xD(304)(4);
  VNStageIntLLRInputS2xD(326)(4) <= CNStageIntLLROutputS2xD(304)(5);
  VNStageIntLLRInputS2xD(3)(4) <= CNStageIntLLROutputS2xD(305)(0);
  VNStageIntLLRInputS2xD(112)(5) <= CNStageIntLLROutputS2xD(305)(1);
  VNStageIntLLRInputS2xD(129)(5) <= CNStageIntLLROutputS2xD(305)(2);
  VNStageIntLLRInputS2xD(220)(5) <= CNStageIntLLROutputS2xD(305)(3);
  VNStageIntLLRInputS2xD(261)(4) <= CNStageIntLLROutputS2xD(305)(4);
  VNStageIntLLRInputS2xD(358)(4) <= CNStageIntLLROutputS2xD(305)(5);
  VNStageIntLLRInputS2xD(2)(5) <= CNStageIntLLROutputS2xD(306)(0);
  VNStageIntLLRInputS2xD(127)(5) <= CNStageIntLLROutputS2xD(306)(1);
  VNStageIntLLRInputS2xD(155)(5) <= CNStageIntLLROutputS2xD(306)(2);
  VNStageIntLLRInputS2xD(196)(5) <= CNStageIntLLROutputS2xD(306)(3);
  VNStageIntLLRInputS2xD(293)(4) <= CNStageIntLLROutputS2xD(306)(4);
  VNStageIntLLRInputS2xD(374)(5) <= CNStageIntLLROutputS2xD(306)(5);
  VNStageIntLLRInputS2xD(1)(4) <= CNStageIntLLROutputS2xD(307)(0);
  VNStageIntLLRInputS2xD(90)(5) <= CNStageIntLLROutputS2xD(307)(1);
  VNStageIntLLRInputS2xD(131)(4) <= CNStageIntLLROutputS2xD(307)(2);
  VNStageIntLLRInputS2xD(228)(5) <= CNStageIntLLROutputS2xD(307)(3);
  VNStageIntLLRInputS2xD(309)(5) <= CNStageIntLLROutputS2xD(307)(4);
  VNStageIntLLRInputS2xD(344)(5) <= CNStageIntLLROutputS2xD(307)(5);
  VNStageIntLLRInputS2xD(62)(4) <= CNStageIntLLROutputS2xD(308)(0);
  VNStageIntLLRInputS2xD(98)(4) <= CNStageIntLLROutputS2xD(308)(1);
  VNStageIntLLRInputS2xD(179)(5) <= CNStageIntLLROutputS2xD(308)(2);
  VNStageIntLLRInputS2xD(214)(5) <= CNStageIntLLROutputS2xD(308)(3);
  VNStageIntLLRInputS2xD(288)(5) <= CNStageIntLLROutputS2xD(308)(4);
  VNStageIntLLRInputS2xD(366)(5) <= CNStageIntLLROutputS2xD(308)(5);
  VNStageIntLLRInputS2xD(61)(4) <= CNStageIntLLROutputS2xD(309)(0);
  VNStageIntLLRInputS2xD(114)(5) <= CNStageIntLLROutputS2xD(309)(1);
  VNStageIntLLRInputS2xD(149)(5) <= CNStageIntLLROutputS2xD(309)(2);
  VNStageIntLLRInputS2xD(223)(5) <= CNStageIntLLROutputS2xD(309)(3);
  VNStageIntLLRInputS2xD(301)(5) <= CNStageIntLLROutputS2xD(309)(4);
  VNStageIntLLRInputS2xD(345)(4) <= CNStageIntLLROutputS2xD(309)(5);
  VNStageIntLLRInputS2xD(60)(4) <= CNStageIntLLROutputS2xD(310)(0);
  VNStageIntLLRInputS2xD(84)(4) <= CNStageIntLLROutputS2xD(310)(1);
  VNStageIntLLRInputS2xD(158)(5) <= CNStageIntLLROutputS2xD(310)(2);
  VNStageIntLLRInputS2xD(236)(5) <= CNStageIntLLROutputS2xD(310)(3);
  VNStageIntLLRInputS2xD(280)(5) <= CNStageIntLLROutputS2xD(310)(4);
  VNStageIntLLRInputS2xD(373)(3) <= CNStageIntLLROutputS2xD(310)(5);
  VNStageIntLLRInputS2xD(59)(3) <= CNStageIntLLROutputS2xD(311)(0);
  VNStageIntLLRInputS2xD(93)(5) <= CNStageIntLLROutputS2xD(311)(1);
  VNStageIntLLRInputS2xD(171)(3) <= CNStageIntLLROutputS2xD(311)(2);
  VNStageIntLLRInputS2xD(215)(5) <= CNStageIntLLROutputS2xD(311)(3);
  VNStageIntLLRInputS2xD(308)(3) <= CNStageIntLLROutputS2xD(311)(4);
  VNStageIntLLRInputS2xD(375)(4) <= CNStageIntLLROutputS2xD(311)(5);
  VNStageIntLLRInputS2xD(58)(3) <= CNStageIntLLROutputS2xD(312)(0);
  VNStageIntLLRInputS2xD(106)(4) <= CNStageIntLLROutputS2xD(312)(1);
  VNStageIntLLRInputS2xD(150)(4) <= CNStageIntLLROutputS2xD(312)(2);
  VNStageIntLLRInputS2xD(243)(5) <= CNStageIntLLROutputS2xD(312)(3);
  VNStageIntLLRInputS2xD(310)(4) <= CNStageIntLLROutputS2xD(312)(4);
  VNStageIntLLRInputS2xD(357)(5) <= CNStageIntLLROutputS2xD(312)(5);
  VNStageIntLLRInputS2xD(57)(4) <= CNStageIntLLROutputS2xD(313)(0);
  VNStageIntLLRInputS2xD(85)(4) <= CNStageIntLLROutputS2xD(313)(1);
  VNStageIntLLRInputS2xD(178)(4) <= CNStageIntLLROutputS2xD(313)(2);
  VNStageIntLLRInputS2xD(245)(5) <= CNStageIntLLROutputS2xD(313)(3);
  VNStageIntLLRInputS2xD(292)(5) <= CNStageIntLLROutputS2xD(313)(4);
  VNStageIntLLRInputS2xD(364)(5) <= CNStageIntLLROutputS2xD(313)(5);
  VNStageIntLLRInputS2xD(56)(5) <= CNStageIntLLROutputS2xD(314)(0);
  VNStageIntLLRInputS2xD(113)(5) <= CNStageIntLLROutputS2xD(314)(1);
  VNStageIntLLRInputS2xD(180)(3) <= CNStageIntLLROutputS2xD(314)(2);
  VNStageIntLLRInputS2xD(227)(5) <= CNStageIntLLROutputS2xD(314)(3);
  VNStageIntLLRInputS2xD(299)(4) <= CNStageIntLLROutputS2xD(314)(4);
  VNStageIntLLRInputS2xD(328)(3) <= CNStageIntLLROutputS2xD(314)(5);
  VNStageIntLLRInputS2xD(55)(5) <= CNStageIntLLROutputS2xD(315)(0);
  VNStageIntLLRInputS2xD(115)(5) <= CNStageIntLLROutputS2xD(315)(1);
  VNStageIntLLRInputS2xD(162)(5) <= CNStageIntLLROutputS2xD(315)(2);
  VNStageIntLLRInputS2xD(234)(5) <= CNStageIntLLROutputS2xD(315)(3);
  VNStageIntLLRInputS2xD(263)(5) <= CNStageIntLLROutputS2xD(315)(4);
  VNStageIntLLRInputS2xD(379)(3) <= CNStageIntLLROutputS2xD(315)(5);
  VNStageIntLLRInputS2xD(54)(4) <= CNStageIntLLROutputS2xD(316)(0);
  VNStageIntLLRInputS2xD(97)(5) <= CNStageIntLLROutputS2xD(316)(1);
  VNStageIntLLRInputS2xD(169)(5) <= CNStageIntLLROutputS2xD(316)(2);
  VNStageIntLLRInputS2xD(198)(5) <= CNStageIntLLROutputS2xD(316)(3);
  VNStageIntLLRInputS2xD(314)(2) <= CNStageIntLLROutputS2xD(316)(4);
  VNStageIntLLRInputS2xD(322)(4) <= CNStageIntLLROutputS2xD(316)(5);
  VNStageIntLLRInputS2xD(53)(4) <= CNStageIntLLROutputS2xD(317)(0);
  VNStageIntLLRInputS2xD(104)(5) <= CNStageIntLLROutputS2xD(317)(1);
  VNStageIntLLRInputS2xD(133)(3) <= CNStageIntLLROutputS2xD(317)(2);
  VNStageIntLLRInputS2xD(249)(3) <= CNStageIntLLROutputS2xD(317)(3);
  VNStageIntLLRInputS2xD(257)(5) <= CNStageIntLLROutputS2xD(317)(4);
  VNStageIntLLRInputS2xD(380)(4) <= CNStageIntLLROutputS2xD(317)(5);
  VNStageIntLLRInputS2xD(52)(3) <= CNStageIntLLROutputS2xD(318)(0);
  VNStageIntLLRInputS2xD(68)(4) <= CNStageIntLLROutputS2xD(318)(1);
  VNStageIntLLRInputS2xD(184)(5) <= CNStageIntLLROutputS2xD(318)(2);
  VNStageIntLLRInputS2xD(255)(5) <= CNStageIntLLROutputS2xD(318)(3);
  VNStageIntLLRInputS2xD(315)(4) <= CNStageIntLLROutputS2xD(318)(4);
  VNStageIntLLRInputS2xD(327)(5) <= CNStageIntLLROutputS2xD(318)(5);
  VNStageIntLLRInputS2xD(51)(4) <= CNStageIntLLROutputS2xD(319)(0);
  VNStageIntLLRInputS2xD(119)(4) <= CNStageIntLLROutputS2xD(319)(1);
  VNStageIntLLRInputS2xD(190)(3) <= CNStageIntLLROutputS2xD(319)(2);
  VNStageIntLLRInputS2xD(250)(3) <= CNStageIntLLROutputS2xD(319)(3);
  VNStageIntLLRInputS2xD(262)(4) <= CNStageIntLLROutputS2xD(319)(4);
  VNStageIntLLRInputS2xD(349)(4) <= CNStageIntLLROutputS2xD(319)(5);
  VNStageIntLLRInputS2xD(50)(5) <= CNStageIntLLROutputS2xD(320)(0);
  VNStageIntLLRInputS2xD(125)(2) <= CNStageIntLLROutputS2xD(320)(1);
  VNStageIntLLRInputS2xD(185)(2) <= CNStageIntLLROutputS2xD(320)(2);
  VNStageIntLLRInputS2xD(197)(5) <= CNStageIntLLROutputS2xD(320)(3);
  VNStageIntLLRInputS2xD(284)(5) <= CNStageIntLLROutputS2xD(320)(4);
  VNStageIntLLRInputS2xD(367)(5) <= CNStageIntLLROutputS2xD(320)(5);
  VNStageIntLLRInputS2xD(49)(5) <= CNStageIntLLROutputS2xD(321)(0);
  VNStageIntLLRInputS2xD(120)(2) <= CNStageIntLLROutputS2xD(321)(1);
  VNStageIntLLRInputS2xD(132)(4) <= CNStageIntLLROutputS2xD(321)(2);
  VNStageIntLLRInputS2xD(219)(4) <= CNStageIntLLROutputS2xD(321)(3);
  VNStageIntLLRInputS2xD(302)(5) <= CNStageIntLLROutputS2xD(321)(4);
  VNStageIntLLRInputS2xD(352)(5) <= CNStageIntLLROutputS2xD(321)(5);
  VNStageIntLLRInputS2xD(48)(2) <= CNStageIntLLROutputS2xD(322)(0);
  VNStageIntLLRInputS2xD(67)(2) <= CNStageIntLLROutputS2xD(322)(1);
  VNStageIntLLRInputS2xD(154)(4) <= CNStageIntLLROutputS2xD(322)(2);
  VNStageIntLLRInputS2xD(237)(4) <= CNStageIntLLROutputS2xD(322)(3);
  VNStageIntLLRInputS2xD(287)(5) <= CNStageIntLLROutputS2xD(322)(4);
  VNStageIntLLRInputS2xD(339)(5) <= CNStageIntLLROutputS2xD(322)(5);
  VNStageIntLLRInputS2xD(46)(5) <= CNStageIntLLROutputS2xD(323)(0);
  VNStageIntLLRInputS2xD(107)(4) <= CNStageIntLLROutputS2xD(323)(1);
  VNStageIntLLRInputS2xD(157)(4) <= CNStageIntLLROutputS2xD(323)(2);
  VNStageIntLLRInputS2xD(209)(4) <= CNStageIntLLROutputS2xD(323)(3);
  VNStageIntLLRInputS2xD(305)(5) <= CNStageIntLLROutputS2xD(323)(4);
  VNStageIntLLRInputS2xD(382)(4) <= CNStageIntLLROutputS2xD(323)(5);
  VNStageIntLLRInputS2xD(45)(5) <= CNStageIntLLROutputS2xD(324)(0);
  VNStageIntLLRInputS2xD(92)(5) <= CNStageIntLLROutputS2xD(324)(1);
  VNStageIntLLRInputS2xD(144)(5) <= CNStageIntLLROutputS2xD(324)(2);
  VNStageIntLLRInputS2xD(240)(5) <= CNStageIntLLROutputS2xD(324)(3);
  VNStageIntLLRInputS2xD(317)(2) <= CNStageIntLLROutputS2xD(324)(4);
  VNStageIntLLRInputS2xD(333)(4) <= CNStageIntLLROutputS2xD(324)(5);
  VNStageIntLLRInputS2xD(44)(5) <= CNStageIntLLROutputS2xD(325)(0);
  VNStageIntLLRInputS2xD(79)(4) <= CNStageIntLLROutputS2xD(325)(1);
  VNStageIntLLRInputS2xD(175)(5) <= CNStageIntLLROutputS2xD(325)(2);
  VNStageIntLLRInputS2xD(252)(4) <= CNStageIntLLROutputS2xD(325)(3);
  VNStageIntLLRInputS2xD(268)(5) <= CNStageIntLLROutputS2xD(325)(4);
  VNStageIntLLRInputS2xD(377)(3) <= CNStageIntLLROutputS2xD(325)(5);
  VNStageIntLLRInputS2xD(43)(4) <= CNStageIntLLROutputS2xD(326)(0);
  VNStageIntLLRInputS2xD(110)(5) <= CNStageIntLLROutputS2xD(326)(1);
  VNStageIntLLRInputS2xD(187)(4) <= CNStageIntLLROutputS2xD(326)(2);
  VNStageIntLLRInputS2xD(203)(5) <= CNStageIntLLROutputS2xD(326)(3);
  VNStageIntLLRInputS2xD(312)(4) <= CNStageIntLLROutputS2xD(326)(4);
  VNStageIntLLRInputS2xD(354)(4) <= CNStageIntLLROutputS2xD(326)(5);
  VNStageIntLLRInputS2xD(42)(5) <= CNStageIntLLROutputS2xD(327)(0);
  VNStageIntLLRInputS2xD(122)(4) <= CNStageIntLLROutputS2xD(327)(1);
  VNStageIntLLRInputS2xD(138)(5) <= CNStageIntLLROutputS2xD(327)(2);
  VNStageIntLLRInputS2xD(247)(5) <= CNStageIntLLROutputS2xD(327)(3);
  VNStageIntLLRInputS2xD(289)(5) <= CNStageIntLLROutputS2xD(327)(4);
  VNStageIntLLRInputS2xD(343)(5) <= CNStageIntLLROutputS2xD(327)(5);
  VNStageIntLLRInputS2xD(41)(5) <= CNStageIntLLROutputS2xD(328)(0);
  VNStageIntLLRInputS2xD(73)(4) <= CNStageIntLLROutputS2xD(328)(1);
  VNStageIntLLRInputS2xD(182)(5) <= CNStageIntLLROutputS2xD(328)(2);
  VNStageIntLLRInputS2xD(224)(5) <= CNStageIntLLROutputS2xD(328)(3);
  VNStageIntLLRInputS2xD(278)(4) <= CNStageIntLLROutputS2xD(328)(4);
  VNStageIntLLRInputS2xD(347)(5) <= CNStageIntLLROutputS2xD(328)(5);
  VNStageIntLLRInputS2xD(39)(5) <= CNStageIntLLROutputS2xD(329)(0);
  VNStageIntLLRInputS2xD(94)(3) <= CNStageIntLLROutputS2xD(329)(1);
  VNStageIntLLRInputS2xD(148)(5) <= CNStageIntLLROutputS2xD(329)(2);
  VNStageIntLLRInputS2xD(217)(5) <= CNStageIntLLROutputS2xD(329)(3);
  VNStageIntLLRInputS2xD(275)(4) <= CNStageIntLLROutputS2xD(329)(4);
  VNStageIntLLRInputS2xD(351)(4) <= CNStageIntLLROutputS2xD(329)(5);
  VNStageIntLLRInputS2xD(38)(5) <= CNStageIntLLROutputS2xD(330)(0);
  VNStageIntLLRInputS2xD(83)(5) <= CNStageIntLLROutputS2xD(330)(1);
  VNStageIntLLRInputS2xD(152)(5) <= CNStageIntLLROutputS2xD(330)(2);
  VNStageIntLLRInputS2xD(210)(5) <= CNStageIntLLROutputS2xD(330)(3);
  VNStageIntLLRInputS2xD(286)(5) <= CNStageIntLLROutputS2xD(330)(4);
  VNStageIntLLRInputS2xD(323)(4) <= CNStageIntLLROutputS2xD(330)(5);
  VNStageIntLLRInputS2xD(37)(5) <= CNStageIntLLROutputS2xD(331)(0);
  VNStageIntLLRInputS2xD(87)(5) <= CNStageIntLLROutputS2xD(331)(1);
  VNStageIntLLRInputS2xD(145)(5) <= CNStageIntLLROutputS2xD(331)(2);
  VNStageIntLLRInputS2xD(221)(5) <= CNStageIntLLROutputS2xD(331)(3);
  VNStageIntLLRInputS2xD(258)(2) <= CNStageIntLLROutputS2xD(331)(4);
  VNStageIntLLRInputS2xD(378)(4) <= CNStageIntLLROutputS2xD(331)(5);
  VNStageIntLLRInputS2xD(0)(5) <= CNStageIntLLROutputS2xD(332)(0);
  VNStageIntLLRInputS2xD(76)(5) <= CNStageIntLLROutputS2xD(332)(1);
  VNStageIntLLRInputS2xD(141)(3) <= CNStageIntLLROutputS2xD(332)(2);
  VNStageIntLLRInputS2xD(206)(3) <= CNStageIntLLROutputS2xD(332)(3);
  VNStageIntLLRInputS2xD(271)(4) <= CNStageIntLLROutputS2xD(332)(4);
  VNStageIntLLRInputS2xD(336)(4) <= CNStageIntLLROutputS2xD(332)(5);
  VNStageIntLLRInputS2xD(28)(5) <= CNStageIntLLROutputS2xD(333)(0);
  VNStageIntLLRInputS2xD(106)(5) <= CNStageIntLLROutputS2xD(333)(1);
  VNStageIntLLRInputS2xD(144)(6) <= CNStageIntLLROutputS2xD(333)(2);
  VNStageIntLLRInputS2xD(193)(4) <= CNStageIntLLROutputS2xD(333)(3);
  VNStageIntLLRInputS2xD(261)(5) <= CNStageIntLLROutputS2xD(333)(4);
  VNStageIntLLRInputS2xD(367)(6) <= CNStageIntLLROutputS2xD(333)(5);
  VNStageIntLLRInputS2xD(26)(6) <= CNStageIntLLROutputS2xD(334)(0);
  VNStageIntLLRInputS2xD(126)(5) <= CNStageIntLLROutputS2xD(334)(1);
  VNStageIntLLRInputS2xD(131)(5) <= CNStageIntLLROutputS2xD(334)(2);
  VNStageIntLLRInputS2xD(237)(5) <= CNStageIntLLROutputS2xD(334)(3);
  VNStageIntLLRInputS2xD(277)(6) <= CNStageIntLLROutputS2xD(334)(4);
  VNStageIntLLRInputS2xD(340)(5) <= CNStageIntLLROutputS2xD(334)(5);
  VNStageIntLLRInputS2xD(24)(6) <= CNStageIntLLROutputS2xD(335)(0);
  VNStageIntLLRInputS2xD(107)(5) <= CNStageIntLLROutputS2xD(335)(1);
  VNStageIntLLRInputS2xD(147)(6) <= CNStageIntLLROutputS2xD(335)(2);
  VNStageIntLLRInputS2xD(210)(6) <= CNStageIntLLROutputS2xD(335)(3);
  VNStageIntLLRInputS2xD(300)(5) <= CNStageIntLLROutputS2xD(335)(4);
  VNStageIntLLRInputS2xD(373)(4) <= CNStageIntLLROutputS2xD(335)(5);
  VNStageIntLLRInputS2xD(23)(6) <= CNStageIntLLROutputS2xD(336)(0);
  VNStageIntLLRInputS2xD(82)(6) <= CNStageIntLLROutputS2xD(336)(1);
  VNStageIntLLRInputS2xD(145)(6) <= CNStageIntLLROutputS2xD(336)(2);
  VNStageIntLLRInputS2xD(235)(4) <= CNStageIntLLROutputS2xD(336)(3);
  VNStageIntLLRInputS2xD(308)(4) <= CNStageIntLLROutputS2xD(336)(4);
  VNStageIntLLRInputS2xD(353)(5) <= CNStageIntLLROutputS2xD(336)(5);
  VNStageIntLLRInputS2xD(22)(6) <= CNStageIntLLROutputS2xD(337)(0);
  VNStageIntLLRInputS2xD(80)(5) <= CNStageIntLLROutputS2xD(337)(1);
  VNStageIntLLRInputS2xD(170)(4) <= CNStageIntLLROutputS2xD(337)(2);
  VNStageIntLLRInputS2xD(243)(6) <= CNStageIntLLROutputS2xD(337)(3);
  VNStageIntLLRInputS2xD(288)(6) <= CNStageIntLLROutputS2xD(337)(4);
  VNStageIntLLRInputS2xD(347)(6) <= CNStageIntLLROutputS2xD(337)(5);
  VNStageIntLLRInputS2xD(21)(6) <= CNStageIntLLROutputS2xD(338)(0);
  VNStageIntLLRInputS2xD(105)(5) <= CNStageIntLLROutputS2xD(338)(1);
  VNStageIntLLRInputS2xD(178)(5) <= CNStageIntLLROutputS2xD(338)(2);
  VNStageIntLLRInputS2xD(223)(6) <= CNStageIntLLROutputS2xD(338)(3);
  VNStageIntLLRInputS2xD(282)(5) <= CNStageIntLLROutputS2xD(338)(4);
  VNStageIntLLRInputS2xD(320)(4) <= CNStageIntLLROutputS2xD(338)(5);
  VNStageIntLLRInputS2xD(20)(4) <= CNStageIntLLROutputS2xD(339)(0);
  VNStageIntLLRInputS2xD(113)(6) <= CNStageIntLLROutputS2xD(339)(1);
  VNStageIntLLRInputS2xD(158)(6) <= CNStageIntLLROutputS2xD(339)(2);
  VNStageIntLLRInputS2xD(217)(6) <= CNStageIntLLROutputS2xD(339)(3);
  VNStageIntLLRInputS2xD(256)(5) <= CNStageIntLLROutputS2xD(339)(4);
  VNStageIntLLRInputS2xD(346)(6) <= CNStageIntLLROutputS2xD(339)(5);
  VNStageIntLLRInputS2xD(19)(4) <= CNStageIntLLROutputS2xD(340)(0);
  VNStageIntLLRInputS2xD(93)(6) <= CNStageIntLLROutputS2xD(340)(1);
  VNStageIntLLRInputS2xD(152)(6) <= CNStageIntLLROutputS2xD(340)(2);
  VNStageIntLLRInputS2xD(192)(6) <= CNStageIntLLROutputS2xD(340)(3);
  VNStageIntLLRInputS2xD(281)(6) <= CNStageIntLLROutputS2xD(340)(4);
  VNStageIntLLRInputS2xD(351)(5) <= CNStageIntLLROutputS2xD(340)(5);
  VNStageIntLLRInputS2xD(18)(6) <= CNStageIntLLROutputS2xD(341)(0);
  VNStageIntLLRInputS2xD(87)(6) <= CNStageIntLLROutputS2xD(341)(1);
  VNStageIntLLRInputS2xD(128)(6) <= CNStageIntLLROutputS2xD(341)(2);
  VNStageIntLLRInputS2xD(216)(6) <= CNStageIntLLROutputS2xD(341)(3);
  VNStageIntLLRInputS2xD(286)(6) <= CNStageIntLLROutputS2xD(341)(4);
  VNStageIntLLRInputS2xD(370)(4) <= CNStageIntLLROutputS2xD(341)(5);
  VNStageIntLLRInputS2xD(17)(6) <= CNStageIntLLROutputS2xD(342)(0);
  VNStageIntLLRInputS2xD(64)(5) <= CNStageIntLLROutputS2xD(342)(1);
  VNStageIntLLRInputS2xD(151)(5) <= CNStageIntLLROutputS2xD(342)(2);
  VNStageIntLLRInputS2xD(221)(6) <= CNStageIntLLROutputS2xD(342)(3);
  VNStageIntLLRInputS2xD(305)(6) <= CNStageIntLLROutputS2xD(342)(4);
  VNStageIntLLRInputS2xD(361)(6) <= CNStageIntLLROutputS2xD(342)(5);
  VNStageIntLLRInputS2xD(16)(5) <= CNStageIntLLROutputS2xD(343)(0);
  VNStageIntLLRInputS2xD(86)(3) <= CNStageIntLLROutputS2xD(343)(1);
  VNStageIntLLRInputS2xD(156)(3) <= CNStageIntLLROutputS2xD(343)(2);
  VNStageIntLLRInputS2xD(240)(6) <= CNStageIntLLROutputS2xD(343)(3);
  VNStageIntLLRInputS2xD(296)(5) <= CNStageIntLLROutputS2xD(343)(4);
  VNStageIntLLRInputS2xD(335)(6) <= CNStageIntLLROutputS2xD(343)(5);
  VNStageIntLLRInputS2xD(15)(6) <= CNStageIntLLROutputS2xD(344)(0);
  VNStageIntLLRInputS2xD(91)(6) <= CNStageIntLLROutputS2xD(344)(1);
  VNStageIntLLRInputS2xD(175)(6) <= CNStageIntLLROutputS2xD(344)(2);
  VNStageIntLLRInputS2xD(231)(5) <= CNStageIntLLROutputS2xD(344)(3);
  VNStageIntLLRInputS2xD(270)(6) <= CNStageIntLLROutputS2xD(344)(4);
  VNStageIntLLRInputS2xD(336)(5) <= CNStageIntLLROutputS2xD(344)(5);
  VNStageIntLLRInputS2xD(14)(6) <= CNStageIntLLROutputS2xD(345)(0);
  VNStageIntLLRInputS2xD(110)(6) <= CNStageIntLLROutputS2xD(345)(1);
  VNStageIntLLRInputS2xD(166)(5) <= CNStageIntLLROutputS2xD(345)(2);
  VNStageIntLLRInputS2xD(205)(2) <= CNStageIntLLROutputS2xD(345)(3);
  VNStageIntLLRInputS2xD(271)(5) <= CNStageIntLLROutputS2xD(345)(4);
  VNStageIntLLRInputS2xD(360)(6) <= CNStageIntLLROutputS2xD(345)(5);
  VNStageIntLLRInputS2xD(13)(5) <= CNStageIntLLROutputS2xD(346)(0);
  VNStageIntLLRInputS2xD(101)(6) <= CNStageIntLLROutputS2xD(346)(1);
  VNStageIntLLRInputS2xD(140)(6) <= CNStageIntLLROutputS2xD(346)(2);
  VNStageIntLLRInputS2xD(206)(4) <= CNStageIntLLROutputS2xD(346)(3);
  VNStageIntLLRInputS2xD(295)(4) <= CNStageIntLLROutputS2xD(346)(4);
  VNStageIntLLRInputS2xD(381)(5) <= CNStageIntLLROutputS2xD(346)(5);
  VNStageIntLLRInputS2xD(12)(6) <= CNStageIntLLROutputS2xD(347)(0);
  VNStageIntLLRInputS2xD(75)(6) <= CNStageIntLLROutputS2xD(347)(1);
  VNStageIntLLRInputS2xD(141)(4) <= CNStageIntLLROutputS2xD(347)(2);
  VNStageIntLLRInputS2xD(230)(5) <= CNStageIntLLROutputS2xD(347)(3);
  VNStageIntLLRInputS2xD(316)(4) <= CNStageIntLLROutputS2xD(347)(4);
  VNStageIntLLRInputS2xD(377)(4) <= CNStageIntLLROutputS2xD(347)(5);
  VNStageIntLLRInputS2xD(11)(5) <= CNStageIntLLROutputS2xD(348)(0);
  VNStageIntLLRInputS2xD(76)(6) <= CNStageIntLLROutputS2xD(348)(1);
  VNStageIntLLRInputS2xD(165)(5) <= CNStageIntLLROutputS2xD(348)(2);
  VNStageIntLLRInputS2xD(251)(4) <= CNStageIntLLROutputS2xD(348)(3);
  VNStageIntLLRInputS2xD(312)(5) <= CNStageIntLLROutputS2xD(348)(4);
  VNStageIntLLRInputS2xD(329)(6) <= CNStageIntLLROutputS2xD(348)(5);
  VNStageIntLLRInputS2xD(10)(4) <= CNStageIntLLROutputS2xD(349)(0);
  VNStageIntLLRInputS2xD(100)(6) <= CNStageIntLLROutputS2xD(349)(1);
  VNStageIntLLRInputS2xD(186)(5) <= CNStageIntLLROutputS2xD(349)(2);
  VNStageIntLLRInputS2xD(247)(6) <= CNStageIntLLROutputS2xD(349)(3);
  VNStageIntLLRInputS2xD(264)(6) <= CNStageIntLLROutputS2xD(349)(4);
  VNStageIntLLRInputS2xD(355)(6) <= CNStageIntLLROutputS2xD(349)(5);
  VNStageIntLLRInputS2xD(9)(6) <= CNStageIntLLROutputS2xD(350)(0);
  VNStageIntLLRInputS2xD(121)(5) <= CNStageIntLLROutputS2xD(350)(1);
  VNStageIntLLRInputS2xD(182)(6) <= CNStageIntLLROutputS2xD(350)(2);
  VNStageIntLLRInputS2xD(199)(6) <= CNStageIntLLROutputS2xD(350)(3);
  VNStageIntLLRInputS2xD(290)(5) <= CNStageIntLLROutputS2xD(350)(4);
  VNStageIntLLRInputS2xD(331)(4) <= CNStageIntLLROutputS2xD(350)(5);
  VNStageIntLLRInputS2xD(7)(6) <= CNStageIntLLROutputS2xD(351)(0);
  VNStageIntLLRInputS2xD(69)(6) <= CNStageIntLLROutputS2xD(351)(1);
  VNStageIntLLRInputS2xD(160)(6) <= CNStageIntLLROutputS2xD(351)(2);
  VNStageIntLLRInputS2xD(201)(5) <= CNStageIntLLROutputS2xD(351)(3);
  VNStageIntLLRInputS2xD(298)(6) <= CNStageIntLLROutputS2xD(351)(4);
  VNStageIntLLRInputS2xD(379)(4) <= CNStageIntLLROutputS2xD(351)(5);
  VNStageIntLLRInputS2xD(6)(6) <= CNStageIntLLROutputS2xD(352)(0);
  VNStageIntLLRInputS2xD(95)(6) <= CNStageIntLLROutputS2xD(352)(1);
  VNStageIntLLRInputS2xD(136)(6) <= CNStageIntLLROutputS2xD(352)(2);
  VNStageIntLLRInputS2xD(233)(4) <= CNStageIntLLROutputS2xD(352)(3);
  VNStageIntLLRInputS2xD(314)(3) <= CNStageIntLLROutputS2xD(352)(4);
  VNStageIntLLRInputS2xD(349)(5) <= CNStageIntLLROutputS2xD(352)(5);
  VNStageIntLLRInputS2xD(5)(6) <= CNStageIntLLROutputS2xD(353)(0);
  VNStageIntLLRInputS2xD(71)(5) <= CNStageIntLLROutputS2xD(353)(1);
  VNStageIntLLRInputS2xD(168)(5) <= CNStageIntLLROutputS2xD(353)(2);
  VNStageIntLLRInputS2xD(249)(4) <= CNStageIntLLROutputS2xD(353)(3);
  VNStageIntLLRInputS2xD(284)(6) <= CNStageIntLLROutputS2xD(353)(4);
  VNStageIntLLRInputS2xD(358)(5) <= CNStageIntLLROutputS2xD(353)(5);
  VNStageIntLLRInputS2xD(4)(5) <= CNStageIntLLROutputS2xD(354)(0);
  VNStageIntLLRInputS2xD(103)(6) <= CNStageIntLLROutputS2xD(354)(1);
  VNStageIntLLRInputS2xD(184)(6) <= CNStageIntLLROutputS2xD(354)(2);
  VNStageIntLLRInputS2xD(219)(5) <= CNStageIntLLROutputS2xD(354)(3);
  VNStageIntLLRInputS2xD(293)(5) <= CNStageIntLLROutputS2xD(354)(4);
  VNStageIntLLRInputS2xD(371)(4) <= CNStageIntLLROutputS2xD(354)(5);
  VNStageIntLLRInputS2xD(2)(6) <= CNStageIntLLROutputS2xD(355)(0);
  VNStageIntLLRInputS2xD(89)(5) <= CNStageIntLLROutputS2xD(355)(1);
  VNStageIntLLRInputS2xD(163)(4) <= CNStageIntLLROutputS2xD(355)(2);
  VNStageIntLLRInputS2xD(241)(5) <= CNStageIntLLROutputS2xD(355)(3);
  VNStageIntLLRInputS2xD(285)(6) <= CNStageIntLLROutputS2xD(355)(4);
  VNStageIntLLRInputS2xD(378)(5) <= CNStageIntLLROutputS2xD(355)(5);
  VNStageIntLLRInputS2xD(1)(5) <= CNStageIntLLROutputS2xD(356)(0);
  VNStageIntLLRInputS2xD(98)(5) <= CNStageIntLLROutputS2xD(356)(1);
  VNStageIntLLRInputS2xD(176)(6) <= CNStageIntLLROutputS2xD(356)(2);
  VNStageIntLLRInputS2xD(220)(6) <= CNStageIntLLROutputS2xD(356)(3);
  VNStageIntLLRInputS2xD(313)(3) <= CNStageIntLLROutputS2xD(356)(4);
  VNStageIntLLRInputS2xD(380)(5) <= CNStageIntLLROutputS2xD(356)(5);
  VNStageIntLLRInputS2xD(63)(3) <= CNStageIntLLROutputS2xD(357)(0);
  VNStageIntLLRInputS2xD(111)(6) <= CNStageIntLLROutputS2xD(357)(1);
  VNStageIntLLRInputS2xD(155)(6) <= CNStageIntLLROutputS2xD(357)(2);
  VNStageIntLLRInputS2xD(248)(6) <= CNStageIntLLROutputS2xD(357)(3);
  VNStageIntLLRInputS2xD(315)(5) <= CNStageIntLLROutputS2xD(357)(4);
  VNStageIntLLRInputS2xD(362)(6) <= CNStageIntLLROutputS2xD(357)(5);
  VNStageIntLLRInputS2xD(62)(5) <= CNStageIntLLROutputS2xD(358)(0);
  VNStageIntLLRInputS2xD(90)(6) <= CNStageIntLLROutputS2xD(358)(1);
  VNStageIntLLRInputS2xD(183)(4) <= CNStageIntLLROutputS2xD(358)(2);
  VNStageIntLLRInputS2xD(250)(4) <= CNStageIntLLROutputS2xD(358)(3);
  VNStageIntLLRInputS2xD(297)(6) <= CNStageIntLLROutputS2xD(358)(4);
  VNStageIntLLRInputS2xD(369)(4) <= CNStageIntLLROutputS2xD(358)(5);
  VNStageIntLLRInputS2xD(61)(5) <= CNStageIntLLROutputS2xD(359)(0);
  VNStageIntLLRInputS2xD(118)(5) <= CNStageIntLLROutputS2xD(359)(1);
  VNStageIntLLRInputS2xD(185)(3) <= CNStageIntLLROutputS2xD(359)(2);
  VNStageIntLLRInputS2xD(232)(5) <= CNStageIntLLROutputS2xD(359)(3);
  VNStageIntLLRInputS2xD(304)(6) <= CNStageIntLLROutputS2xD(359)(4);
  VNStageIntLLRInputS2xD(333)(5) <= CNStageIntLLROutputS2xD(359)(5);
  VNStageIntLLRInputS2xD(60)(5) <= CNStageIntLLROutputS2xD(360)(0);
  VNStageIntLLRInputS2xD(120)(3) <= CNStageIntLLROutputS2xD(360)(1);
  VNStageIntLLRInputS2xD(167)(6) <= CNStageIntLLROutputS2xD(360)(2);
  VNStageIntLLRInputS2xD(239)(6) <= CNStageIntLLROutputS2xD(360)(3);
  VNStageIntLLRInputS2xD(268)(6) <= CNStageIntLLROutputS2xD(360)(4);
  VNStageIntLLRInputS2xD(321)(6) <= CNStageIntLLROutputS2xD(360)(5);
  VNStageIntLLRInputS2xD(59)(4) <= CNStageIntLLROutputS2xD(361)(0);
  VNStageIntLLRInputS2xD(102)(5) <= CNStageIntLLROutputS2xD(361)(1);
  VNStageIntLLRInputS2xD(174)(4) <= CNStageIntLLROutputS2xD(361)(2);
  VNStageIntLLRInputS2xD(203)(6) <= CNStageIntLLROutputS2xD(361)(3);
  VNStageIntLLRInputS2xD(319)(6) <= CNStageIntLLROutputS2xD(361)(4);
  VNStageIntLLRInputS2xD(327)(6) <= CNStageIntLLROutputS2xD(361)(5);
  VNStageIntLLRInputS2xD(58)(4) <= CNStageIntLLROutputS2xD(362)(0);
  VNStageIntLLRInputS2xD(109)(5) <= CNStageIntLLROutputS2xD(362)(1);
  VNStageIntLLRInputS2xD(138)(6) <= CNStageIntLLROutputS2xD(362)(2);
  VNStageIntLLRInputS2xD(254)(4) <= CNStageIntLLROutputS2xD(362)(3);
  VNStageIntLLRInputS2xD(262)(5) <= CNStageIntLLROutputS2xD(362)(4);
  VNStageIntLLRInputS2xD(322)(5) <= CNStageIntLLROutputS2xD(362)(5);
  VNStageIntLLRInputS2xD(57)(5) <= CNStageIntLLROutputS2xD(363)(0);
  VNStageIntLLRInputS2xD(73)(5) <= CNStageIntLLROutputS2xD(363)(1);
  VNStageIntLLRInputS2xD(189)(5) <= CNStageIntLLROutputS2xD(363)(2);
  VNStageIntLLRInputS2xD(197)(6) <= CNStageIntLLROutputS2xD(363)(3);
  VNStageIntLLRInputS2xD(257)(6) <= CNStageIntLLROutputS2xD(363)(4);
  VNStageIntLLRInputS2xD(332)(5) <= CNStageIntLLROutputS2xD(363)(5);
  VNStageIntLLRInputS2xD(56)(6) <= CNStageIntLLROutputS2xD(364)(0);
  VNStageIntLLRInputS2xD(124)(4) <= CNStageIntLLROutputS2xD(364)(1);
  VNStageIntLLRInputS2xD(132)(5) <= CNStageIntLLROutputS2xD(364)(2);
  VNStageIntLLRInputS2xD(255)(6) <= CNStageIntLLROutputS2xD(364)(3);
  VNStageIntLLRInputS2xD(267)(6) <= CNStageIntLLROutputS2xD(364)(4);
  VNStageIntLLRInputS2xD(354)(5) <= CNStageIntLLROutputS2xD(364)(5);
  VNStageIntLLRInputS2xD(55)(6) <= CNStageIntLLROutputS2xD(365)(0);
  VNStageIntLLRInputS2xD(67)(3) <= CNStageIntLLROutputS2xD(365)(1);
  VNStageIntLLRInputS2xD(190)(4) <= CNStageIntLLROutputS2xD(365)(2);
  VNStageIntLLRInputS2xD(202)(5) <= CNStageIntLLROutputS2xD(365)(3);
  VNStageIntLLRInputS2xD(289)(6) <= CNStageIntLLROutputS2xD(365)(4);
  VNStageIntLLRInputS2xD(372)(5) <= CNStageIntLLROutputS2xD(365)(5);
  VNStageIntLLRInputS2xD(54)(5) <= CNStageIntLLROutputS2xD(366)(0);
  VNStageIntLLRInputS2xD(125)(3) <= CNStageIntLLROutputS2xD(366)(1);
  VNStageIntLLRInputS2xD(137)(6) <= CNStageIntLLROutputS2xD(366)(2);
  VNStageIntLLRInputS2xD(224)(6) <= CNStageIntLLROutputS2xD(366)(3);
  VNStageIntLLRInputS2xD(307)(6) <= CNStageIntLLROutputS2xD(366)(4);
  VNStageIntLLRInputS2xD(357)(6) <= CNStageIntLLROutputS2xD(366)(5);
  VNStageIntLLRInputS2xD(53)(5) <= CNStageIntLLROutputS2xD(367)(0);
  VNStageIntLLRInputS2xD(72)(5) <= CNStageIntLLROutputS2xD(367)(1);
  VNStageIntLLRInputS2xD(159)(4) <= CNStageIntLLROutputS2xD(367)(2);
  VNStageIntLLRInputS2xD(242)(6) <= CNStageIntLLROutputS2xD(367)(3);
  VNStageIntLLRInputS2xD(292)(6) <= CNStageIntLLROutputS2xD(367)(4);
  VNStageIntLLRInputS2xD(344)(6) <= CNStageIntLLROutputS2xD(367)(5);
  VNStageIntLLRInputS2xD(52)(4) <= CNStageIntLLROutputS2xD(368)(0);
  VNStageIntLLRInputS2xD(94)(4) <= CNStageIntLLROutputS2xD(368)(1);
  VNStageIntLLRInputS2xD(177)(6) <= CNStageIntLLROutputS2xD(368)(2);
  VNStageIntLLRInputS2xD(227)(6) <= CNStageIntLLROutputS2xD(368)(3);
  VNStageIntLLRInputS2xD(279)(5) <= CNStageIntLLROutputS2xD(368)(4);
  VNStageIntLLRInputS2xD(375)(5) <= CNStageIntLLROutputS2xD(368)(5);
  VNStageIntLLRInputS2xD(51)(5) <= CNStageIntLLROutputS2xD(369)(0);
  VNStageIntLLRInputS2xD(112)(6) <= CNStageIntLLROutputS2xD(369)(1);
  VNStageIntLLRInputS2xD(162)(6) <= CNStageIntLLROutputS2xD(369)(2);
  VNStageIntLLRInputS2xD(214)(6) <= CNStageIntLLROutputS2xD(369)(3);
  VNStageIntLLRInputS2xD(310)(5) <= CNStageIntLLROutputS2xD(369)(4);
  VNStageIntLLRInputS2xD(324)(6) <= CNStageIntLLROutputS2xD(369)(5);
  VNStageIntLLRInputS2xD(50)(6) <= CNStageIntLLROutputS2xD(370)(0);
  VNStageIntLLRInputS2xD(97)(6) <= CNStageIntLLROutputS2xD(370)(1);
  VNStageIntLLRInputS2xD(149)(6) <= CNStageIntLLROutputS2xD(370)(2);
  VNStageIntLLRInputS2xD(245)(6) <= CNStageIntLLROutputS2xD(370)(3);
  VNStageIntLLRInputS2xD(259)(4) <= CNStageIntLLROutputS2xD(370)(4);
  VNStageIntLLRInputS2xD(338)(4) <= CNStageIntLLROutputS2xD(370)(5);
  VNStageIntLLRInputS2xD(49)(6) <= CNStageIntLLROutputS2xD(371)(0);
  VNStageIntLLRInputS2xD(84)(5) <= CNStageIntLLROutputS2xD(371)(1);
  VNStageIntLLRInputS2xD(180)(4) <= CNStageIntLLROutputS2xD(371)(2);
  VNStageIntLLRInputS2xD(194)(6) <= CNStageIntLLROutputS2xD(371)(3);
  VNStageIntLLRInputS2xD(273)(5) <= CNStageIntLLROutputS2xD(371)(4);
  VNStageIntLLRInputS2xD(382)(5) <= CNStageIntLLROutputS2xD(371)(5);
  VNStageIntLLRInputS2xD(48)(3) <= CNStageIntLLROutputS2xD(372)(0);
  VNStageIntLLRInputS2xD(115)(6) <= CNStageIntLLROutputS2xD(372)(1);
  VNStageIntLLRInputS2xD(129)(6) <= CNStageIntLLROutputS2xD(372)(2);
  VNStageIntLLRInputS2xD(208)(5) <= CNStageIntLLROutputS2xD(372)(3);
  VNStageIntLLRInputS2xD(317)(3) <= CNStageIntLLROutputS2xD(372)(4);
  VNStageIntLLRInputS2xD(359)(6) <= CNStageIntLLROutputS2xD(372)(5);
  VNStageIntLLRInputS2xD(47)(3) <= CNStageIntLLROutputS2xD(373)(0);
  VNStageIntLLRInputS2xD(127)(6) <= CNStageIntLLROutputS2xD(373)(1);
  VNStageIntLLRInputS2xD(143)(6) <= CNStageIntLLROutputS2xD(373)(2);
  VNStageIntLLRInputS2xD(252)(5) <= CNStageIntLLROutputS2xD(373)(3);
  VNStageIntLLRInputS2xD(294)(6) <= CNStageIntLLROutputS2xD(373)(4);
  VNStageIntLLRInputS2xD(348)(6) <= CNStageIntLLROutputS2xD(373)(5);
  VNStageIntLLRInputS2xD(46)(6) <= CNStageIntLLROutputS2xD(374)(0);
  VNStageIntLLRInputS2xD(78)(6) <= CNStageIntLLROutputS2xD(374)(1);
  VNStageIntLLRInputS2xD(187)(5) <= CNStageIntLLROutputS2xD(374)(2);
  VNStageIntLLRInputS2xD(229)(4) <= CNStageIntLLROutputS2xD(374)(3);
  VNStageIntLLRInputS2xD(283)(6) <= CNStageIntLLROutputS2xD(374)(4);
  VNStageIntLLRInputS2xD(352)(6) <= CNStageIntLLROutputS2xD(374)(5);
  VNStageIntLLRInputS2xD(45)(6) <= CNStageIntLLROutputS2xD(375)(0);
  VNStageIntLLRInputS2xD(122)(5) <= CNStageIntLLROutputS2xD(375)(1);
  VNStageIntLLRInputS2xD(164)(5) <= CNStageIntLLROutputS2xD(375)(2);
  VNStageIntLLRInputS2xD(218)(6) <= CNStageIntLLROutputS2xD(375)(3);
  VNStageIntLLRInputS2xD(287)(6) <= CNStageIntLLROutputS2xD(375)(4);
  VNStageIntLLRInputS2xD(345)(5) <= CNStageIntLLROutputS2xD(375)(5);
  VNStageIntLLRInputS2xD(44)(6) <= CNStageIntLLROutputS2xD(376)(0);
  VNStageIntLLRInputS2xD(99)(6) <= CNStageIntLLROutputS2xD(376)(1);
  VNStageIntLLRInputS2xD(153)(6) <= CNStageIntLLROutputS2xD(376)(2);
  VNStageIntLLRInputS2xD(222)(3) <= CNStageIntLLROutputS2xD(376)(3);
  VNStageIntLLRInputS2xD(280)(6) <= CNStageIntLLROutputS2xD(376)(4);
  VNStageIntLLRInputS2xD(356)(5) <= CNStageIntLLROutputS2xD(376)(5);
  VNStageIntLLRInputS2xD(43)(5) <= CNStageIntLLROutputS2xD(377)(0);
  VNStageIntLLRInputS2xD(88)(6) <= CNStageIntLLROutputS2xD(377)(1);
  VNStageIntLLRInputS2xD(157)(5) <= CNStageIntLLROutputS2xD(377)(2);
  VNStageIntLLRInputS2xD(215)(6) <= CNStageIntLLROutputS2xD(377)(3);
  VNStageIntLLRInputS2xD(291)(5) <= CNStageIntLLROutputS2xD(377)(4);
  VNStageIntLLRInputS2xD(328)(4) <= CNStageIntLLROutputS2xD(377)(5);
  VNStageIntLLRInputS2xD(42)(6) <= CNStageIntLLROutputS2xD(378)(0);
  VNStageIntLLRInputS2xD(92)(6) <= CNStageIntLLROutputS2xD(378)(1);
  VNStageIntLLRInputS2xD(150)(5) <= CNStageIntLLROutputS2xD(378)(2);
  VNStageIntLLRInputS2xD(226)(2) <= CNStageIntLLROutputS2xD(378)(3);
  VNStageIntLLRInputS2xD(263)(6) <= CNStageIntLLROutputS2xD(378)(4);
  VNStageIntLLRInputS2xD(383)(6) <= CNStageIntLLROutputS2xD(378)(5);
  VNStageIntLLRInputS2xD(41)(6) <= CNStageIntLLROutputS2xD(379)(0);
  VNStageIntLLRInputS2xD(85)(5) <= CNStageIntLLROutputS2xD(379)(1);
  VNStageIntLLRInputS2xD(161)(6) <= CNStageIntLLROutputS2xD(379)(2);
  VNStageIntLLRInputS2xD(198)(6) <= CNStageIntLLROutputS2xD(379)(3);
  VNStageIntLLRInputS2xD(318)(3) <= CNStageIntLLROutputS2xD(379)(4);
  VNStageIntLLRInputS2xD(337)(6) <= CNStageIntLLROutputS2xD(379)(5);
  VNStageIntLLRInputS2xD(40)(4) <= CNStageIntLLROutputS2xD(380)(0);
  VNStageIntLLRInputS2xD(96)(5) <= CNStageIntLLROutputS2xD(380)(1);
  VNStageIntLLRInputS2xD(133)(4) <= CNStageIntLLROutputS2xD(380)(2);
  VNStageIntLLRInputS2xD(253)(5) <= CNStageIntLLROutputS2xD(380)(3);
  VNStageIntLLRInputS2xD(272)(6) <= CNStageIntLLROutputS2xD(380)(4);
  VNStageIntLLRInputS2xD(334)(4) <= CNStageIntLLROutputS2xD(380)(5);
  VNStageIntLLRInputS2xD(39)(6) <= CNStageIntLLROutputS2xD(381)(0);
  VNStageIntLLRInputS2xD(68)(5) <= CNStageIntLLROutputS2xD(381)(1);
  VNStageIntLLRInputS2xD(188)(4) <= CNStageIntLLROutputS2xD(381)(2);
  VNStageIntLLRInputS2xD(207)(5) <= CNStageIntLLROutputS2xD(381)(3);
  VNStageIntLLRInputS2xD(269)(5) <= CNStageIntLLROutputS2xD(381)(4);
  VNStageIntLLRInputS2xD(368)(2) <= CNStageIntLLROutputS2xD(381)(5);
  VNStageIntLLRInputS2xD(38)(6) <= CNStageIntLLROutputS2xD(382)(0);
  VNStageIntLLRInputS2xD(123)(4) <= CNStageIntLLROutputS2xD(382)(1);
  VNStageIntLLRInputS2xD(142)(4) <= CNStageIntLLROutputS2xD(382)(2);
  VNStageIntLLRInputS2xD(204)(6) <= CNStageIntLLROutputS2xD(382)(3);
  VNStageIntLLRInputS2xD(303)(6) <= CNStageIntLLROutputS2xD(382)(4);
  VNStageIntLLRInputS2xD(325)(6) <= CNStageIntLLROutputS2xD(382)(5);
  VNStageIntLLRInputS2xD(37)(6) <= CNStageIntLLROutputS2xD(383)(0);
  VNStageIntLLRInputS2xD(77)(4) <= CNStageIntLLROutputS2xD(383)(1);
  VNStageIntLLRInputS2xD(139)(6) <= CNStageIntLLROutputS2xD(383)(2);
  VNStageIntLLRInputS2xD(238)(6) <= CNStageIntLLROutputS2xD(383)(3);
  VNStageIntLLRInputS2xD(260)(5) <= CNStageIntLLROutputS2xD(383)(4);
  VNStageIntLLRInputS2xD(374)(6) <= CNStageIntLLROutputS2xD(383)(5);

  -- Check Nodes (Iteration 3)
  CNStageIntLLRInputS3xD(53)(0) <= VNStageIntLLROutputS2xD(0)(0);
  CNStageIntLLRInputS3xD(110)(0) <= VNStageIntLLROutputS2xD(0)(1);
  CNStageIntLLRInputS3xD(170)(0) <= VNStageIntLLROutputS2xD(0)(2);
  CNStageIntLLRInputS3xD(224)(0) <= VNStageIntLLROutputS2xD(0)(3);
  CNStageIntLLRInputS3xD(279)(0) <= VNStageIntLLROutputS2xD(0)(4);
  CNStageIntLLRInputS3xD(332)(0) <= VNStageIntLLROutputS2xD(0)(5);
  CNStageIntLLRInputS3xD(51)(0) <= VNStageIntLLROutputS2xD(1)(0);
  CNStageIntLLRInputS3xD(139)(0) <= VNStageIntLLROutputS2xD(1)(1);
  CNStageIntLLRInputS3xD(223)(0) <= VNStageIntLLROutputS2xD(1)(2);
  CNStageIntLLRInputS3xD(241)(0) <= VNStageIntLLROutputS2xD(1)(3);
  CNStageIntLLRInputS3xD(307)(0) <= VNStageIntLLROutputS2xD(1)(4);
  CNStageIntLLRInputS3xD(356)(0) <= VNStageIntLLROutputS2xD(1)(5);
  CNStageIntLLRInputS3xD(50)(0) <= VNStageIntLLROutputS2xD(2)(0);
  CNStageIntLLRInputS3xD(92)(0) <= VNStageIntLLROutputS2xD(2)(1);
  CNStageIntLLRInputS3xD(138)(0) <= VNStageIntLLROutputS2xD(2)(2);
  CNStageIntLLRInputS3xD(222)(0) <= VNStageIntLLROutputS2xD(2)(3);
  CNStageIntLLRInputS3xD(240)(0) <= VNStageIntLLROutputS2xD(2)(4);
  CNStageIntLLRInputS3xD(306)(0) <= VNStageIntLLROutputS2xD(2)(5);
  CNStageIntLLRInputS3xD(355)(0) <= VNStageIntLLROutputS2xD(2)(6);
  CNStageIntLLRInputS3xD(91)(0) <= VNStageIntLLROutputS2xD(3)(0);
  CNStageIntLLRInputS3xD(137)(0) <= VNStageIntLLROutputS2xD(3)(1);
  CNStageIntLLRInputS3xD(221)(0) <= VNStageIntLLROutputS2xD(3)(2);
  CNStageIntLLRInputS3xD(239)(0) <= VNStageIntLLROutputS2xD(3)(3);
  CNStageIntLLRInputS3xD(305)(0) <= VNStageIntLLROutputS2xD(3)(4);
  CNStageIntLLRInputS3xD(49)(0) <= VNStageIntLLROutputS2xD(4)(0);
  CNStageIntLLRInputS3xD(90)(0) <= VNStageIntLLROutputS2xD(4)(1);
  CNStageIntLLRInputS3xD(220)(0) <= VNStageIntLLROutputS2xD(4)(2);
  CNStageIntLLRInputS3xD(238)(0) <= VNStageIntLLROutputS2xD(4)(3);
  CNStageIntLLRInputS3xD(304)(0) <= VNStageIntLLROutputS2xD(4)(4);
  CNStageIntLLRInputS3xD(354)(0) <= VNStageIntLLROutputS2xD(4)(5);
  CNStageIntLLRInputS3xD(48)(0) <= VNStageIntLLROutputS2xD(5)(0);
  CNStageIntLLRInputS3xD(89)(0) <= VNStageIntLLROutputS2xD(5)(1);
  CNStageIntLLRInputS3xD(136)(0) <= VNStageIntLLROutputS2xD(5)(2);
  CNStageIntLLRInputS3xD(219)(0) <= VNStageIntLLROutputS2xD(5)(3);
  CNStageIntLLRInputS3xD(237)(0) <= VNStageIntLLROutputS2xD(5)(4);
  CNStageIntLLRInputS3xD(303)(0) <= VNStageIntLLROutputS2xD(5)(5);
  CNStageIntLLRInputS3xD(353)(0) <= VNStageIntLLROutputS2xD(5)(6);
  CNStageIntLLRInputS3xD(47)(0) <= VNStageIntLLROutputS2xD(6)(0);
  CNStageIntLLRInputS3xD(88)(0) <= VNStageIntLLROutputS2xD(6)(1);
  CNStageIntLLRInputS3xD(135)(0) <= VNStageIntLLROutputS2xD(6)(2);
  CNStageIntLLRInputS3xD(218)(0) <= VNStageIntLLROutputS2xD(6)(3);
  CNStageIntLLRInputS3xD(236)(0) <= VNStageIntLLROutputS2xD(6)(4);
  CNStageIntLLRInputS3xD(302)(0) <= VNStageIntLLROutputS2xD(6)(5);
  CNStageIntLLRInputS3xD(352)(0) <= VNStageIntLLROutputS2xD(6)(6);
  CNStageIntLLRInputS3xD(46)(0) <= VNStageIntLLROutputS2xD(7)(0);
  CNStageIntLLRInputS3xD(87)(0) <= VNStageIntLLROutputS2xD(7)(1);
  CNStageIntLLRInputS3xD(134)(0) <= VNStageIntLLROutputS2xD(7)(2);
  CNStageIntLLRInputS3xD(217)(0) <= VNStageIntLLROutputS2xD(7)(3);
  CNStageIntLLRInputS3xD(235)(0) <= VNStageIntLLROutputS2xD(7)(4);
  CNStageIntLLRInputS3xD(301)(0) <= VNStageIntLLROutputS2xD(7)(5);
  CNStageIntLLRInputS3xD(351)(0) <= VNStageIntLLROutputS2xD(7)(6);
  CNStageIntLLRInputS3xD(45)(0) <= VNStageIntLLROutputS2xD(8)(0);
  CNStageIntLLRInputS3xD(133)(0) <= VNStageIntLLROutputS2xD(8)(1);
  CNStageIntLLRInputS3xD(216)(0) <= VNStageIntLLROutputS2xD(8)(2);
  CNStageIntLLRInputS3xD(44)(0) <= VNStageIntLLROutputS2xD(9)(0);
  CNStageIntLLRInputS3xD(86)(0) <= VNStageIntLLROutputS2xD(9)(1);
  CNStageIntLLRInputS3xD(132)(0) <= VNStageIntLLROutputS2xD(9)(2);
  CNStageIntLLRInputS3xD(215)(0) <= VNStageIntLLROutputS2xD(9)(3);
  CNStageIntLLRInputS3xD(234)(0) <= VNStageIntLLROutputS2xD(9)(4);
  CNStageIntLLRInputS3xD(300)(0) <= VNStageIntLLROutputS2xD(9)(5);
  CNStageIntLLRInputS3xD(350)(0) <= VNStageIntLLROutputS2xD(9)(6);
  CNStageIntLLRInputS3xD(43)(0) <= VNStageIntLLROutputS2xD(10)(0);
  CNStageIntLLRInputS3xD(85)(0) <= VNStageIntLLROutputS2xD(10)(1);
  CNStageIntLLRInputS3xD(131)(0) <= VNStageIntLLROutputS2xD(10)(2);
  CNStageIntLLRInputS3xD(233)(0) <= VNStageIntLLROutputS2xD(10)(3);
  CNStageIntLLRInputS3xD(349)(0) <= VNStageIntLLROutputS2xD(10)(4);
  CNStageIntLLRInputS3xD(42)(0) <= VNStageIntLLROutputS2xD(11)(0);
  CNStageIntLLRInputS3xD(84)(0) <= VNStageIntLLROutputS2xD(11)(1);
  CNStageIntLLRInputS3xD(130)(0) <= VNStageIntLLROutputS2xD(11)(2);
  CNStageIntLLRInputS3xD(214)(0) <= VNStageIntLLROutputS2xD(11)(3);
  CNStageIntLLRInputS3xD(232)(0) <= VNStageIntLLROutputS2xD(11)(4);
  CNStageIntLLRInputS3xD(348)(0) <= VNStageIntLLROutputS2xD(11)(5);
  CNStageIntLLRInputS3xD(41)(0) <= VNStageIntLLROutputS2xD(12)(0);
  CNStageIntLLRInputS3xD(83)(0) <= VNStageIntLLROutputS2xD(12)(1);
  CNStageIntLLRInputS3xD(129)(0) <= VNStageIntLLROutputS2xD(12)(2);
  CNStageIntLLRInputS3xD(213)(0) <= VNStageIntLLROutputS2xD(12)(3);
  CNStageIntLLRInputS3xD(231)(0) <= VNStageIntLLROutputS2xD(12)(4);
  CNStageIntLLRInputS3xD(299)(0) <= VNStageIntLLROutputS2xD(12)(5);
  CNStageIntLLRInputS3xD(347)(0) <= VNStageIntLLROutputS2xD(12)(6);
  CNStageIntLLRInputS3xD(82)(0) <= VNStageIntLLROutputS2xD(13)(0);
  CNStageIntLLRInputS3xD(128)(0) <= VNStageIntLLROutputS2xD(13)(1);
  CNStageIntLLRInputS3xD(212)(0) <= VNStageIntLLROutputS2xD(13)(2);
  CNStageIntLLRInputS3xD(230)(0) <= VNStageIntLLROutputS2xD(13)(3);
  CNStageIntLLRInputS3xD(298)(0) <= VNStageIntLLROutputS2xD(13)(4);
  CNStageIntLLRInputS3xD(346)(0) <= VNStageIntLLROutputS2xD(13)(5);
  CNStageIntLLRInputS3xD(40)(0) <= VNStageIntLLROutputS2xD(14)(0);
  CNStageIntLLRInputS3xD(81)(0) <= VNStageIntLLROutputS2xD(14)(1);
  CNStageIntLLRInputS3xD(127)(0) <= VNStageIntLLROutputS2xD(14)(2);
  CNStageIntLLRInputS3xD(211)(0) <= VNStageIntLLROutputS2xD(14)(3);
  CNStageIntLLRInputS3xD(229)(0) <= VNStageIntLLROutputS2xD(14)(4);
  CNStageIntLLRInputS3xD(297)(0) <= VNStageIntLLROutputS2xD(14)(5);
  CNStageIntLLRInputS3xD(345)(0) <= VNStageIntLLROutputS2xD(14)(6);
  CNStageIntLLRInputS3xD(39)(0) <= VNStageIntLLROutputS2xD(15)(0);
  CNStageIntLLRInputS3xD(80)(0) <= VNStageIntLLROutputS2xD(15)(1);
  CNStageIntLLRInputS3xD(126)(0) <= VNStageIntLLROutputS2xD(15)(2);
  CNStageIntLLRInputS3xD(210)(0) <= VNStageIntLLROutputS2xD(15)(3);
  CNStageIntLLRInputS3xD(228)(0) <= VNStageIntLLROutputS2xD(15)(4);
  CNStageIntLLRInputS3xD(296)(0) <= VNStageIntLLROutputS2xD(15)(5);
  CNStageIntLLRInputS3xD(344)(0) <= VNStageIntLLROutputS2xD(15)(6);
  CNStageIntLLRInputS3xD(38)(0) <= VNStageIntLLROutputS2xD(16)(0);
  CNStageIntLLRInputS3xD(125)(0) <= VNStageIntLLROutputS2xD(16)(1);
  CNStageIntLLRInputS3xD(209)(0) <= VNStageIntLLROutputS2xD(16)(2);
  CNStageIntLLRInputS3xD(227)(0) <= VNStageIntLLROutputS2xD(16)(3);
  CNStageIntLLRInputS3xD(295)(0) <= VNStageIntLLROutputS2xD(16)(4);
  CNStageIntLLRInputS3xD(343)(0) <= VNStageIntLLROutputS2xD(16)(5);
  CNStageIntLLRInputS3xD(37)(0) <= VNStageIntLLROutputS2xD(17)(0);
  CNStageIntLLRInputS3xD(79)(0) <= VNStageIntLLROutputS2xD(17)(1);
  CNStageIntLLRInputS3xD(124)(0) <= VNStageIntLLROutputS2xD(17)(2);
  CNStageIntLLRInputS3xD(208)(0) <= VNStageIntLLROutputS2xD(17)(3);
  CNStageIntLLRInputS3xD(226)(0) <= VNStageIntLLROutputS2xD(17)(4);
  CNStageIntLLRInputS3xD(294)(0) <= VNStageIntLLROutputS2xD(17)(5);
  CNStageIntLLRInputS3xD(342)(0) <= VNStageIntLLROutputS2xD(17)(6);
  CNStageIntLLRInputS3xD(36)(0) <= VNStageIntLLROutputS2xD(18)(0);
  CNStageIntLLRInputS3xD(78)(0) <= VNStageIntLLROutputS2xD(18)(1);
  CNStageIntLLRInputS3xD(123)(0) <= VNStageIntLLROutputS2xD(18)(2);
  CNStageIntLLRInputS3xD(207)(0) <= VNStageIntLLROutputS2xD(18)(3);
  CNStageIntLLRInputS3xD(225)(0) <= VNStageIntLLROutputS2xD(18)(4);
  CNStageIntLLRInputS3xD(293)(0) <= VNStageIntLLROutputS2xD(18)(5);
  CNStageIntLLRInputS3xD(341)(0) <= VNStageIntLLROutputS2xD(18)(6);
  CNStageIntLLRInputS3xD(35)(0) <= VNStageIntLLROutputS2xD(19)(0);
  CNStageIntLLRInputS3xD(77)(0) <= VNStageIntLLROutputS2xD(19)(1);
  CNStageIntLLRInputS3xD(122)(0) <= VNStageIntLLROutputS2xD(19)(2);
  CNStageIntLLRInputS3xD(278)(0) <= VNStageIntLLROutputS2xD(19)(3);
  CNStageIntLLRInputS3xD(340)(0) <= VNStageIntLLROutputS2xD(19)(4);
  CNStageIntLLRInputS3xD(34)(0) <= VNStageIntLLROutputS2xD(20)(0);
  CNStageIntLLRInputS3xD(76)(0) <= VNStageIntLLROutputS2xD(20)(1);
  CNStageIntLLRInputS3xD(277)(0) <= VNStageIntLLROutputS2xD(20)(2);
  CNStageIntLLRInputS3xD(292)(0) <= VNStageIntLLROutputS2xD(20)(3);
  CNStageIntLLRInputS3xD(339)(0) <= VNStageIntLLROutputS2xD(20)(4);
  CNStageIntLLRInputS3xD(33)(0) <= VNStageIntLLROutputS2xD(21)(0);
  CNStageIntLLRInputS3xD(75)(0) <= VNStageIntLLROutputS2xD(21)(1);
  CNStageIntLLRInputS3xD(121)(0) <= VNStageIntLLROutputS2xD(21)(2);
  CNStageIntLLRInputS3xD(206)(0) <= VNStageIntLLROutputS2xD(21)(3);
  CNStageIntLLRInputS3xD(276)(0) <= VNStageIntLLROutputS2xD(21)(4);
  CNStageIntLLRInputS3xD(291)(0) <= VNStageIntLLROutputS2xD(21)(5);
  CNStageIntLLRInputS3xD(338)(0) <= VNStageIntLLROutputS2xD(21)(6);
  CNStageIntLLRInputS3xD(32)(0) <= VNStageIntLLROutputS2xD(22)(0);
  CNStageIntLLRInputS3xD(74)(0) <= VNStageIntLLROutputS2xD(22)(1);
  CNStageIntLLRInputS3xD(120)(0) <= VNStageIntLLROutputS2xD(22)(2);
  CNStageIntLLRInputS3xD(205)(0) <= VNStageIntLLROutputS2xD(22)(3);
  CNStageIntLLRInputS3xD(275)(0) <= VNStageIntLLROutputS2xD(22)(4);
  CNStageIntLLRInputS3xD(290)(0) <= VNStageIntLLROutputS2xD(22)(5);
  CNStageIntLLRInputS3xD(337)(0) <= VNStageIntLLROutputS2xD(22)(6);
  CNStageIntLLRInputS3xD(31)(0) <= VNStageIntLLROutputS2xD(23)(0);
  CNStageIntLLRInputS3xD(73)(0) <= VNStageIntLLROutputS2xD(23)(1);
  CNStageIntLLRInputS3xD(119)(0) <= VNStageIntLLROutputS2xD(23)(2);
  CNStageIntLLRInputS3xD(204)(0) <= VNStageIntLLROutputS2xD(23)(3);
  CNStageIntLLRInputS3xD(274)(0) <= VNStageIntLLROutputS2xD(23)(4);
  CNStageIntLLRInputS3xD(289)(0) <= VNStageIntLLROutputS2xD(23)(5);
  CNStageIntLLRInputS3xD(336)(0) <= VNStageIntLLROutputS2xD(23)(6);
  CNStageIntLLRInputS3xD(30)(0) <= VNStageIntLLROutputS2xD(24)(0);
  CNStageIntLLRInputS3xD(72)(0) <= VNStageIntLLROutputS2xD(24)(1);
  CNStageIntLLRInputS3xD(118)(0) <= VNStageIntLLROutputS2xD(24)(2);
  CNStageIntLLRInputS3xD(203)(0) <= VNStageIntLLROutputS2xD(24)(3);
  CNStageIntLLRInputS3xD(273)(0) <= VNStageIntLLROutputS2xD(24)(4);
  CNStageIntLLRInputS3xD(288)(0) <= VNStageIntLLROutputS2xD(24)(5);
  CNStageIntLLRInputS3xD(335)(0) <= VNStageIntLLROutputS2xD(24)(6);
  CNStageIntLLRInputS3xD(29)(0) <= VNStageIntLLROutputS2xD(25)(0);
  CNStageIntLLRInputS3xD(71)(0) <= VNStageIntLLROutputS2xD(25)(1);
  CNStageIntLLRInputS3xD(117)(0) <= VNStageIntLLROutputS2xD(25)(2);
  CNStageIntLLRInputS3xD(202)(0) <= VNStageIntLLROutputS2xD(25)(3);
  CNStageIntLLRInputS3xD(287)(0) <= VNStageIntLLROutputS2xD(25)(4);
  CNStageIntLLRInputS3xD(28)(0) <= VNStageIntLLROutputS2xD(26)(0);
  CNStageIntLLRInputS3xD(70)(0) <= VNStageIntLLROutputS2xD(26)(1);
  CNStageIntLLRInputS3xD(116)(0) <= VNStageIntLLROutputS2xD(26)(2);
  CNStageIntLLRInputS3xD(201)(0) <= VNStageIntLLROutputS2xD(26)(3);
  CNStageIntLLRInputS3xD(272)(0) <= VNStageIntLLROutputS2xD(26)(4);
  CNStageIntLLRInputS3xD(286)(0) <= VNStageIntLLROutputS2xD(26)(5);
  CNStageIntLLRInputS3xD(334)(0) <= VNStageIntLLROutputS2xD(26)(6);
  CNStageIntLLRInputS3xD(27)(0) <= VNStageIntLLROutputS2xD(27)(0);
  CNStageIntLLRInputS3xD(69)(0) <= VNStageIntLLROutputS2xD(27)(1);
  CNStageIntLLRInputS3xD(115)(0) <= VNStageIntLLROutputS2xD(27)(2);
  CNStageIntLLRInputS3xD(200)(0) <= VNStageIntLLROutputS2xD(27)(3);
  CNStageIntLLRInputS3xD(285)(0) <= VNStageIntLLROutputS2xD(27)(4);
  CNStageIntLLRInputS3xD(26)(0) <= VNStageIntLLROutputS2xD(28)(0);
  CNStageIntLLRInputS3xD(68)(0) <= VNStageIntLLROutputS2xD(28)(1);
  CNStageIntLLRInputS3xD(114)(0) <= VNStageIntLLROutputS2xD(28)(2);
  CNStageIntLLRInputS3xD(199)(0) <= VNStageIntLLROutputS2xD(28)(3);
  CNStageIntLLRInputS3xD(271)(0) <= VNStageIntLLROutputS2xD(28)(4);
  CNStageIntLLRInputS3xD(333)(0) <= VNStageIntLLROutputS2xD(28)(5);
  CNStageIntLLRInputS3xD(25)(0) <= VNStageIntLLROutputS2xD(29)(0);
  CNStageIntLLRInputS3xD(67)(0) <= VNStageIntLLROutputS2xD(29)(1);
  CNStageIntLLRInputS3xD(113)(0) <= VNStageIntLLROutputS2xD(29)(2);
  CNStageIntLLRInputS3xD(270)(0) <= VNStageIntLLROutputS2xD(29)(3);
  CNStageIntLLRInputS3xD(24)(0) <= VNStageIntLLROutputS2xD(30)(0);
  CNStageIntLLRInputS3xD(66)(0) <= VNStageIntLLROutputS2xD(30)(1);
  CNStageIntLLRInputS3xD(112)(0) <= VNStageIntLLROutputS2xD(30)(2);
  CNStageIntLLRInputS3xD(198)(0) <= VNStageIntLLROutputS2xD(30)(3);
  CNStageIntLLRInputS3xD(269)(0) <= VNStageIntLLROutputS2xD(30)(4);
  CNStageIntLLRInputS3xD(284)(0) <= VNStageIntLLROutputS2xD(30)(5);
  CNStageIntLLRInputS3xD(23)(0) <= VNStageIntLLROutputS2xD(31)(0);
  CNStageIntLLRInputS3xD(65)(0) <= VNStageIntLLROutputS2xD(31)(1);
  CNStageIntLLRInputS3xD(197)(0) <= VNStageIntLLROutputS2xD(31)(2);
  CNStageIntLLRInputS3xD(283)(0) <= VNStageIntLLROutputS2xD(31)(3);
  CNStageIntLLRInputS3xD(22)(0) <= VNStageIntLLROutputS2xD(32)(0);
  CNStageIntLLRInputS3xD(64)(0) <= VNStageIntLLROutputS2xD(32)(1);
  CNStageIntLLRInputS3xD(111)(0) <= VNStageIntLLROutputS2xD(32)(2);
  CNStageIntLLRInputS3xD(268)(0) <= VNStageIntLLROutputS2xD(32)(3);
  CNStageIntLLRInputS3xD(21)(0) <= VNStageIntLLROutputS2xD(33)(0);
  CNStageIntLLRInputS3xD(63)(0) <= VNStageIntLLROutputS2xD(33)(1);
  CNStageIntLLRInputS3xD(169)(0) <= VNStageIntLLROutputS2xD(33)(2);
  CNStageIntLLRInputS3xD(196)(0) <= VNStageIntLLROutputS2xD(33)(3);
  CNStageIntLLRInputS3xD(267)(0) <= VNStageIntLLROutputS2xD(33)(4);
  CNStageIntLLRInputS3xD(282)(0) <= VNStageIntLLROutputS2xD(33)(5);
  CNStageIntLLRInputS3xD(20)(0) <= VNStageIntLLROutputS2xD(34)(0);
  CNStageIntLLRInputS3xD(62)(0) <= VNStageIntLLROutputS2xD(34)(1);
  CNStageIntLLRInputS3xD(168)(0) <= VNStageIntLLROutputS2xD(34)(2);
  CNStageIntLLRInputS3xD(195)(0) <= VNStageIntLLROutputS2xD(34)(3);
  CNStageIntLLRInputS3xD(266)(0) <= VNStageIntLLROutputS2xD(34)(4);
  CNStageIntLLRInputS3xD(281)(0) <= VNStageIntLLROutputS2xD(34)(5);
  CNStageIntLLRInputS3xD(19)(0) <= VNStageIntLLROutputS2xD(35)(0);
  CNStageIntLLRInputS3xD(61)(0) <= VNStageIntLLROutputS2xD(35)(1);
  CNStageIntLLRInputS3xD(167)(0) <= VNStageIntLLROutputS2xD(35)(2);
  CNStageIntLLRInputS3xD(194)(0) <= VNStageIntLLROutputS2xD(35)(3);
  CNStageIntLLRInputS3xD(265)(0) <= VNStageIntLLROutputS2xD(35)(4);
  CNStageIntLLRInputS3xD(280)(0) <= VNStageIntLLROutputS2xD(35)(5);
  CNStageIntLLRInputS3xD(18)(0) <= VNStageIntLLROutputS2xD(36)(0);
  CNStageIntLLRInputS3xD(60)(0) <= VNStageIntLLROutputS2xD(36)(1);
  CNStageIntLLRInputS3xD(166)(0) <= VNStageIntLLROutputS2xD(36)(2);
  CNStageIntLLRInputS3xD(264)(0) <= VNStageIntLLROutputS2xD(36)(3);
  CNStageIntLLRInputS3xD(17)(0) <= VNStageIntLLROutputS2xD(37)(0);
  CNStageIntLLRInputS3xD(59)(0) <= VNStageIntLLROutputS2xD(37)(1);
  CNStageIntLLRInputS3xD(165)(0) <= VNStageIntLLROutputS2xD(37)(2);
  CNStageIntLLRInputS3xD(193)(0) <= VNStageIntLLROutputS2xD(37)(3);
  CNStageIntLLRInputS3xD(263)(0) <= VNStageIntLLROutputS2xD(37)(4);
  CNStageIntLLRInputS3xD(331)(0) <= VNStageIntLLROutputS2xD(37)(5);
  CNStageIntLLRInputS3xD(383)(0) <= VNStageIntLLROutputS2xD(37)(6);
  CNStageIntLLRInputS3xD(16)(0) <= VNStageIntLLROutputS2xD(38)(0);
  CNStageIntLLRInputS3xD(58)(0) <= VNStageIntLLROutputS2xD(38)(1);
  CNStageIntLLRInputS3xD(164)(0) <= VNStageIntLLROutputS2xD(38)(2);
  CNStageIntLLRInputS3xD(192)(0) <= VNStageIntLLROutputS2xD(38)(3);
  CNStageIntLLRInputS3xD(262)(0) <= VNStageIntLLROutputS2xD(38)(4);
  CNStageIntLLRInputS3xD(330)(0) <= VNStageIntLLROutputS2xD(38)(5);
  CNStageIntLLRInputS3xD(382)(0) <= VNStageIntLLROutputS2xD(38)(6);
  CNStageIntLLRInputS3xD(15)(0) <= VNStageIntLLROutputS2xD(39)(0);
  CNStageIntLLRInputS3xD(57)(0) <= VNStageIntLLROutputS2xD(39)(1);
  CNStageIntLLRInputS3xD(163)(0) <= VNStageIntLLROutputS2xD(39)(2);
  CNStageIntLLRInputS3xD(191)(0) <= VNStageIntLLROutputS2xD(39)(3);
  CNStageIntLLRInputS3xD(261)(0) <= VNStageIntLLROutputS2xD(39)(4);
  CNStageIntLLRInputS3xD(329)(0) <= VNStageIntLLROutputS2xD(39)(5);
  CNStageIntLLRInputS3xD(381)(0) <= VNStageIntLLROutputS2xD(39)(6);
  CNStageIntLLRInputS3xD(14)(0) <= VNStageIntLLROutputS2xD(40)(0);
  CNStageIntLLRInputS3xD(56)(0) <= VNStageIntLLROutputS2xD(40)(1);
  CNStageIntLLRInputS3xD(162)(0) <= VNStageIntLLROutputS2xD(40)(2);
  CNStageIntLLRInputS3xD(260)(0) <= VNStageIntLLROutputS2xD(40)(3);
  CNStageIntLLRInputS3xD(380)(0) <= VNStageIntLLROutputS2xD(40)(4);
  CNStageIntLLRInputS3xD(13)(0) <= VNStageIntLLROutputS2xD(41)(0);
  CNStageIntLLRInputS3xD(55)(0) <= VNStageIntLLROutputS2xD(41)(1);
  CNStageIntLLRInputS3xD(161)(0) <= VNStageIntLLROutputS2xD(41)(2);
  CNStageIntLLRInputS3xD(190)(0) <= VNStageIntLLROutputS2xD(41)(3);
  CNStageIntLLRInputS3xD(259)(0) <= VNStageIntLLROutputS2xD(41)(4);
  CNStageIntLLRInputS3xD(328)(0) <= VNStageIntLLROutputS2xD(41)(5);
  CNStageIntLLRInputS3xD(379)(0) <= VNStageIntLLROutputS2xD(41)(6);
  CNStageIntLLRInputS3xD(12)(0) <= VNStageIntLLROutputS2xD(42)(0);
  CNStageIntLLRInputS3xD(54)(0) <= VNStageIntLLROutputS2xD(42)(1);
  CNStageIntLLRInputS3xD(160)(0) <= VNStageIntLLROutputS2xD(42)(2);
  CNStageIntLLRInputS3xD(189)(0) <= VNStageIntLLROutputS2xD(42)(3);
  CNStageIntLLRInputS3xD(258)(0) <= VNStageIntLLROutputS2xD(42)(4);
  CNStageIntLLRInputS3xD(327)(0) <= VNStageIntLLROutputS2xD(42)(5);
  CNStageIntLLRInputS3xD(378)(0) <= VNStageIntLLROutputS2xD(42)(6);
  CNStageIntLLRInputS3xD(109)(0) <= VNStageIntLLROutputS2xD(43)(0);
  CNStageIntLLRInputS3xD(159)(0) <= VNStageIntLLROutputS2xD(43)(1);
  CNStageIntLLRInputS3xD(188)(0) <= VNStageIntLLROutputS2xD(43)(2);
  CNStageIntLLRInputS3xD(257)(0) <= VNStageIntLLROutputS2xD(43)(3);
  CNStageIntLLRInputS3xD(326)(0) <= VNStageIntLLROutputS2xD(43)(4);
  CNStageIntLLRInputS3xD(377)(0) <= VNStageIntLLROutputS2xD(43)(5);
  CNStageIntLLRInputS3xD(11)(0) <= VNStageIntLLROutputS2xD(44)(0);
  CNStageIntLLRInputS3xD(108)(0) <= VNStageIntLLROutputS2xD(44)(1);
  CNStageIntLLRInputS3xD(158)(0) <= VNStageIntLLROutputS2xD(44)(2);
  CNStageIntLLRInputS3xD(187)(0) <= VNStageIntLLROutputS2xD(44)(3);
  CNStageIntLLRInputS3xD(256)(0) <= VNStageIntLLROutputS2xD(44)(4);
  CNStageIntLLRInputS3xD(325)(0) <= VNStageIntLLROutputS2xD(44)(5);
  CNStageIntLLRInputS3xD(376)(0) <= VNStageIntLLROutputS2xD(44)(6);
  CNStageIntLLRInputS3xD(10)(0) <= VNStageIntLLROutputS2xD(45)(0);
  CNStageIntLLRInputS3xD(107)(0) <= VNStageIntLLROutputS2xD(45)(1);
  CNStageIntLLRInputS3xD(157)(0) <= VNStageIntLLROutputS2xD(45)(2);
  CNStageIntLLRInputS3xD(186)(0) <= VNStageIntLLROutputS2xD(45)(3);
  CNStageIntLLRInputS3xD(255)(0) <= VNStageIntLLROutputS2xD(45)(4);
  CNStageIntLLRInputS3xD(324)(0) <= VNStageIntLLROutputS2xD(45)(5);
  CNStageIntLLRInputS3xD(375)(0) <= VNStageIntLLROutputS2xD(45)(6);
  CNStageIntLLRInputS3xD(9)(0) <= VNStageIntLLROutputS2xD(46)(0);
  CNStageIntLLRInputS3xD(106)(0) <= VNStageIntLLROutputS2xD(46)(1);
  CNStageIntLLRInputS3xD(156)(0) <= VNStageIntLLROutputS2xD(46)(2);
  CNStageIntLLRInputS3xD(185)(0) <= VNStageIntLLROutputS2xD(46)(3);
  CNStageIntLLRInputS3xD(254)(0) <= VNStageIntLLROutputS2xD(46)(4);
  CNStageIntLLRInputS3xD(323)(0) <= VNStageIntLLROutputS2xD(46)(5);
  CNStageIntLLRInputS3xD(374)(0) <= VNStageIntLLROutputS2xD(46)(6);
  CNStageIntLLRInputS3xD(8)(0) <= VNStageIntLLROutputS2xD(47)(0);
  CNStageIntLLRInputS3xD(155)(0) <= VNStageIntLLROutputS2xD(47)(1);
  CNStageIntLLRInputS3xD(253)(0) <= VNStageIntLLROutputS2xD(47)(2);
  CNStageIntLLRInputS3xD(373)(0) <= VNStageIntLLROutputS2xD(47)(3);
  CNStageIntLLRInputS3xD(7)(0) <= VNStageIntLLROutputS2xD(48)(0);
  CNStageIntLLRInputS3xD(154)(0) <= VNStageIntLLROutputS2xD(48)(1);
  CNStageIntLLRInputS3xD(322)(0) <= VNStageIntLLROutputS2xD(48)(2);
  CNStageIntLLRInputS3xD(372)(0) <= VNStageIntLLROutputS2xD(48)(3);
  CNStageIntLLRInputS3xD(6)(0) <= VNStageIntLLROutputS2xD(49)(0);
  CNStageIntLLRInputS3xD(105)(0) <= VNStageIntLLROutputS2xD(49)(1);
  CNStageIntLLRInputS3xD(153)(0) <= VNStageIntLLROutputS2xD(49)(2);
  CNStageIntLLRInputS3xD(184)(0) <= VNStageIntLLROutputS2xD(49)(3);
  CNStageIntLLRInputS3xD(252)(0) <= VNStageIntLLROutputS2xD(49)(4);
  CNStageIntLLRInputS3xD(321)(0) <= VNStageIntLLROutputS2xD(49)(5);
  CNStageIntLLRInputS3xD(371)(0) <= VNStageIntLLROutputS2xD(49)(6);
  CNStageIntLLRInputS3xD(5)(0) <= VNStageIntLLROutputS2xD(50)(0);
  CNStageIntLLRInputS3xD(104)(0) <= VNStageIntLLROutputS2xD(50)(1);
  CNStageIntLLRInputS3xD(152)(0) <= VNStageIntLLROutputS2xD(50)(2);
  CNStageIntLLRInputS3xD(183)(0) <= VNStageIntLLROutputS2xD(50)(3);
  CNStageIntLLRInputS3xD(251)(0) <= VNStageIntLLROutputS2xD(50)(4);
  CNStageIntLLRInputS3xD(320)(0) <= VNStageIntLLROutputS2xD(50)(5);
  CNStageIntLLRInputS3xD(370)(0) <= VNStageIntLLROutputS2xD(50)(6);
  CNStageIntLLRInputS3xD(4)(0) <= VNStageIntLLROutputS2xD(51)(0);
  CNStageIntLLRInputS3xD(103)(0) <= VNStageIntLLROutputS2xD(51)(1);
  CNStageIntLLRInputS3xD(182)(0) <= VNStageIntLLROutputS2xD(51)(2);
  CNStageIntLLRInputS3xD(250)(0) <= VNStageIntLLROutputS2xD(51)(3);
  CNStageIntLLRInputS3xD(319)(0) <= VNStageIntLLROutputS2xD(51)(4);
  CNStageIntLLRInputS3xD(369)(0) <= VNStageIntLLROutputS2xD(51)(5);
  CNStageIntLLRInputS3xD(102)(0) <= VNStageIntLLROutputS2xD(52)(0);
  CNStageIntLLRInputS3xD(151)(0) <= VNStageIntLLROutputS2xD(52)(1);
  CNStageIntLLRInputS3xD(181)(0) <= VNStageIntLLROutputS2xD(52)(2);
  CNStageIntLLRInputS3xD(318)(0) <= VNStageIntLLROutputS2xD(52)(3);
  CNStageIntLLRInputS3xD(368)(0) <= VNStageIntLLROutputS2xD(52)(4);
  CNStageIntLLRInputS3xD(3)(0) <= VNStageIntLLROutputS2xD(53)(0);
  CNStageIntLLRInputS3xD(150)(0) <= VNStageIntLLROutputS2xD(53)(1);
  CNStageIntLLRInputS3xD(180)(0) <= VNStageIntLLROutputS2xD(53)(2);
  CNStageIntLLRInputS3xD(249)(0) <= VNStageIntLLROutputS2xD(53)(3);
  CNStageIntLLRInputS3xD(317)(0) <= VNStageIntLLROutputS2xD(53)(4);
  CNStageIntLLRInputS3xD(367)(0) <= VNStageIntLLROutputS2xD(53)(5);
  CNStageIntLLRInputS3xD(2)(0) <= VNStageIntLLROutputS2xD(54)(0);
  CNStageIntLLRInputS3xD(101)(0) <= VNStageIntLLROutputS2xD(54)(1);
  CNStageIntLLRInputS3xD(149)(0) <= VNStageIntLLROutputS2xD(54)(2);
  CNStageIntLLRInputS3xD(179)(0) <= VNStageIntLLROutputS2xD(54)(3);
  CNStageIntLLRInputS3xD(316)(0) <= VNStageIntLLROutputS2xD(54)(4);
  CNStageIntLLRInputS3xD(366)(0) <= VNStageIntLLROutputS2xD(54)(5);
  CNStageIntLLRInputS3xD(1)(0) <= VNStageIntLLROutputS2xD(55)(0);
  CNStageIntLLRInputS3xD(100)(0) <= VNStageIntLLROutputS2xD(55)(1);
  CNStageIntLLRInputS3xD(148)(0) <= VNStageIntLLROutputS2xD(55)(2);
  CNStageIntLLRInputS3xD(178)(0) <= VNStageIntLLROutputS2xD(55)(3);
  CNStageIntLLRInputS3xD(248)(0) <= VNStageIntLLROutputS2xD(55)(4);
  CNStageIntLLRInputS3xD(315)(0) <= VNStageIntLLROutputS2xD(55)(5);
  CNStageIntLLRInputS3xD(365)(0) <= VNStageIntLLROutputS2xD(55)(6);
  CNStageIntLLRInputS3xD(0)(0) <= VNStageIntLLROutputS2xD(56)(0);
  CNStageIntLLRInputS3xD(99)(0) <= VNStageIntLLROutputS2xD(56)(1);
  CNStageIntLLRInputS3xD(147)(0) <= VNStageIntLLROutputS2xD(56)(2);
  CNStageIntLLRInputS3xD(177)(0) <= VNStageIntLLROutputS2xD(56)(3);
  CNStageIntLLRInputS3xD(247)(0) <= VNStageIntLLROutputS2xD(56)(4);
  CNStageIntLLRInputS3xD(314)(0) <= VNStageIntLLROutputS2xD(56)(5);
  CNStageIntLLRInputS3xD(364)(0) <= VNStageIntLLROutputS2xD(56)(6);
  CNStageIntLLRInputS3xD(98)(0) <= VNStageIntLLROutputS2xD(57)(0);
  CNStageIntLLRInputS3xD(146)(0) <= VNStageIntLLROutputS2xD(57)(1);
  CNStageIntLLRInputS3xD(176)(0) <= VNStageIntLLROutputS2xD(57)(2);
  CNStageIntLLRInputS3xD(246)(0) <= VNStageIntLLROutputS2xD(57)(3);
  CNStageIntLLRInputS3xD(313)(0) <= VNStageIntLLROutputS2xD(57)(4);
  CNStageIntLLRInputS3xD(363)(0) <= VNStageIntLLROutputS2xD(57)(5);
  CNStageIntLLRInputS3xD(97)(0) <= VNStageIntLLROutputS2xD(58)(0);
  CNStageIntLLRInputS3xD(145)(0) <= VNStageIntLLROutputS2xD(58)(1);
  CNStageIntLLRInputS3xD(175)(0) <= VNStageIntLLROutputS2xD(58)(2);
  CNStageIntLLRInputS3xD(312)(0) <= VNStageIntLLROutputS2xD(58)(3);
  CNStageIntLLRInputS3xD(362)(0) <= VNStageIntLLROutputS2xD(58)(4);
  CNStageIntLLRInputS3xD(144)(0) <= VNStageIntLLROutputS2xD(59)(0);
  CNStageIntLLRInputS3xD(174)(0) <= VNStageIntLLROutputS2xD(59)(1);
  CNStageIntLLRInputS3xD(245)(0) <= VNStageIntLLROutputS2xD(59)(2);
  CNStageIntLLRInputS3xD(311)(0) <= VNStageIntLLROutputS2xD(59)(3);
  CNStageIntLLRInputS3xD(361)(0) <= VNStageIntLLROutputS2xD(59)(4);
  CNStageIntLLRInputS3xD(96)(0) <= VNStageIntLLROutputS2xD(60)(0);
  CNStageIntLLRInputS3xD(143)(0) <= VNStageIntLLROutputS2xD(60)(1);
  CNStageIntLLRInputS3xD(173)(0) <= VNStageIntLLROutputS2xD(60)(2);
  CNStageIntLLRInputS3xD(244)(0) <= VNStageIntLLROutputS2xD(60)(3);
  CNStageIntLLRInputS3xD(310)(0) <= VNStageIntLLROutputS2xD(60)(4);
  CNStageIntLLRInputS3xD(360)(0) <= VNStageIntLLROutputS2xD(60)(5);
  CNStageIntLLRInputS3xD(95)(0) <= VNStageIntLLROutputS2xD(61)(0);
  CNStageIntLLRInputS3xD(142)(0) <= VNStageIntLLROutputS2xD(61)(1);
  CNStageIntLLRInputS3xD(172)(0) <= VNStageIntLLROutputS2xD(61)(2);
  CNStageIntLLRInputS3xD(243)(0) <= VNStageIntLLROutputS2xD(61)(3);
  CNStageIntLLRInputS3xD(309)(0) <= VNStageIntLLROutputS2xD(61)(4);
  CNStageIntLLRInputS3xD(359)(0) <= VNStageIntLLROutputS2xD(61)(5);
  CNStageIntLLRInputS3xD(94)(0) <= VNStageIntLLROutputS2xD(62)(0);
  CNStageIntLLRInputS3xD(141)(0) <= VNStageIntLLROutputS2xD(62)(1);
  CNStageIntLLRInputS3xD(171)(0) <= VNStageIntLLROutputS2xD(62)(2);
  CNStageIntLLRInputS3xD(242)(0) <= VNStageIntLLROutputS2xD(62)(3);
  CNStageIntLLRInputS3xD(308)(0) <= VNStageIntLLROutputS2xD(62)(4);
  CNStageIntLLRInputS3xD(358)(0) <= VNStageIntLLROutputS2xD(62)(5);
  CNStageIntLLRInputS3xD(52)(0) <= VNStageIntLLROutputS2xD(63)(0);
  CNStageIntLLRInputS3xD(93)(0) <= VNStageIntLLROutputS2xD(63)(1);
  CNStageIntLLRInputS3xD(140)(0) <= VNStageIntLLROutputS2xD(63)(2);
  CNStageIntLLRInputS3xD(357)(0) <= VNStageIntLLROutputS2xD(63)(3);
  CNStageIntLLRInputS3xD(53)(1) <= VNStageIntLLROutputS2xD(64)(0);
  CNStageIntLLRInputS3xD(109)(1) <= VNStageIntLLROutputS2xD(64)(1);
  CNStageIntLLRInputS3xD(130)(1) <= VNStageIntLLROutputS2xD(64)(2);
  CNStageIntLLRInputS3xD(245)(1) <= VNStageIntLLROutputS2xD(64)(3);
  CNStageIntLLRInputS3xD(299)(1) <= VNStageIntLLROutputS2xD(64)(4);
  CNStageIntLLRInputS3xD(342)(1) <= VNStageIntLLROutputS2xD(64)(5);
  CNStageIntLLRInputS3xD(51)(1) <= VNStageIntLLROutputS2xD(65)(0);
  CNStageIntLLRInputS3xD(74)(1) <= VNStageIntLLROutputS2xD(65)(1);
  CNStageIntLLRInputS3xD(141)(1) <= VNStageIntLLROutputS2xD(65)(2);
  CNStageIntLLRInputS3xD(189)(1) <= VNStageIntLLROutputS2xD(65)(3);
  CNStageIntLLRInputS3xD(286)(1) <= VNStageIntLLROutputS2xD(65)(4);
  CNStageIntLLRInputS3xD(50)(1) <= VNStageIntLLROutputS2xD(66)(0);
  CNStageIntLLRInputS3xD(66)(1) <= VNStageIntLLROutputS2xD(66)(1);
  CNStageIntLLRInputS3xD(155)(1) <= VNStageIntLLROutputS2xD(66)(2);
  CNStageIntLLRInputS3xD(244)(1) <= VNStageIntLLROutputS2xD(66)(3);
  CNStageIntLLRInputS3xD(97)(1) <= VNStageIntLLROutputS2xD(67)(0);
  CNStageIntLLRInputS3xD(275)(1) <= VNStageIntLLROutputS2xD(67)(1);
  CNStageIntLLRInputS3xD(322)(1) <= VNStageIntLLROutputS2xD(67)(2);
  CNStageIntLLRInputS3xD(365)(1) <= VNStageIntLLROutputS2xD(67)(3);
  CNStageIntLLRInputS3xD(49)(1) <= VNStageIntLLROutputS2xD(68)(0);
  CNStageIntLLRInputS3xD(112)(1) <= VNStageIntLLROutputS2xD(68)(1);
  CNStageIntLLRInputS3xD(210)(1) <= VNStageIntLLROutputS2xD(68)(2);
  CNStageIntLLRInputS3xD(256)(1) <= VNStageIntLLROutputS2xD(68)(3);
  CNStageIntLLRInputS3xD(318)(1) <= VNStageIntLLROutputS2xD(68)(4);
  CNStageIntLLRInputS3xD(381)(1) <= VNStageIntLLROutputS2xD(68)(5);
  CNStageIntLLRInputS3xD(48)(1) <= VNStageIntLLROutputS2xD(69)(0);
  CNStageIntLLRInputS3xD(101)(1) <= VNStageIntLLROutputS2xD(69)(1);
  CNStageIntLLRInputS3xD(135)(1) <= VNStageIntLLROutputS2xD(69)(2);
  CNStageIntLLRInputS3xD(215)(1) <= VNStageIntLLROutputS2xD(69)(3);
  CNStageIntLLRInputS3xD(259)(1) <= VNStageIntLLROutputS2xD(69)(4);
  CNStageIntLLRInputS3xD(283)(1) <= VNStageIntLLROutputS2xD(69)(5);
  CNStageIntLLRInputS3xD(351)(1) <= VNStageIntLLROutputS2xD(69)(6);
  CNStageIntLLRInputS3xD(47)(1) <= VNStageIntLLROutputS2xD(70)(0);
  CNStageIntLLRInputS3xD(104)(1) <= VNStageIntLLROutputS2xD(70)(1);
  CNStageIntLLRInputS3xD(136)(1) <= VNStageIntLLROutputS2xD(70)(2);
  CNStageIntLLRInputS3xD(206)(1) <= VNStageIntLLROutputS2xD(70)(3);
  CNStageIntLLRInputS3xD(246)(1) <= VNStageIntLLROutputS2xD(70)(4);
  CNStageIntLLRInputS3xD(301)(1) <= VNStageIntLLROutputS2xD(70)(5);
  CNStageIntLLRInputS3xD(46)(1) <= VNStageIntLLROutputS2xD(71)(0);
  CNStageIntLLRInputS3xD(95)(1) <= VNStageIntLLROutputS2xD(71)(1);
  CNStageIntLLRInputS3xD(176)(1) <= VNStageIntLLROutputS2xD(71)(2);
  CNStageIntLLRInputS3xD(276)(1) <= VNStageIntLLROutputS2xD(71)(3);
  CNStageIntLLRInputS3xD(302)(1) <= VNStageIntLLROutputS2xD(71)(4);
  CNStageIntLLRInputS3xD(353)(1) <= VNStageIntLLROutputS2xD(71)(5);
  CNStageIntLLRInputS3xD(45)(1) <= VNStageIntLLROutputS2xD(72)(0);
  CNStageIntLLRInputS3xD(75)(1) <= VNStageIntLLROutputS2xD(72)(1);
  CNStageIntLLRInputS3xD(162)(1) <= VNStageIntLLROutputS2xD(72)(2);
  CNStageIntLLRInputS3xD(183)(1) <= VNStageIntLLROutputS2xD(72)(3);
  CNStageIntLLRInputS3xD(243)(1) <= VNStageIntLLROutputS2xD(72)(4);
  CNStageIntLLRInputS3xD(367)(1) <= VNStageIntLLROutputS2xD(72)(5);
  CNStageIntLLRInputS3xD(44)(1) <= VNStageIntLLROutputS2xD(73)(0);
  CNStageIntLLRInputS3xD(56)(1) <= VNStageIntLLROutputS2xD(73)(1);
  CNStageIntLLRInputS3xD(121)(1) <= VNStageIntLLROutputS2xD(73)(2);
  CNStageIntLLRInputS3xD(219)(1) <= VNStageIntLLROutputS2xD(73)(3);
  CNStageIntLLRInputS3xD(328)(1) <= VNStageIntLLROutputS2xD(73)(4);
  CNStageIntLLRInputS3xD(363)(1) <= VNStageIntLLROutputS2xD(73)(5);
  CNStageIntLLRInputS3xD(43)(1) <= VNStageIntLLROutputS2xD(74)(0);
  CNStageIntLLRInputS3xD(70)(1) <= VNStageIntLLROutputS2xD(74)(1);
  CNStageIntLLRInputS3xD(125)(1) <= VNStageIntLLROutputS2xD(74)(2);
  CNStageIntLLRInputS3xD(221)(1) <= VNStageIntLLROutputS2xD(74)(3);
  CNStageIntLLRInputS3xD(290)(1) <= VNStageIntLLROutputS2xD(74)(4);
  CNStageIntLLRInputS3xD(42)(1) <= VNStageIntLLROutputS2xD(75)(0);
  CNStageIntLLRInputS3xD(81)(1) <= VNStageIntLLROutputS2xD(75)(1);
  CNStageIntLLRInputS3xD(170)(1) <= VNStageIntLLROutputS2xD(75)(2);
  CNStageIntLLRInputS3xD(192)(1) <= VNStageIntLLROutputS2xD(75)(3);
  CNStageIntLLRInputS3xD(278)(1) <= VNStageIntLLROutputS2xD(75)(4);
  CNStageIntLLRInputS3xD(294)(1) <= VNStageIntLLROutputS2xD(75)(5);
  CNStageIntLLRInputS3xD(347)(1) <= VNStageIntLLROutputS2xD(75)(6);
  CNStageIntLLRInputS3xD(41)(1) <= VNStageIntLLROutputS2xD(76)(0);
  CNStageIntLLRInputS3xD(106)(1) <= VNStageIntLLROutputS2xD(76)(1);
  CNStageIntLLRInputS3xD(124)(1) <= VNStageIntLLROutputS2xD(76)(2);
  CNStageIntLLRInputS3xD(174)(1) <= VNStageIntLLROutputS2xD(76)(3);
  CNStageIntLLRInputS3xD(270)(1) <= VNStageIntLLROutputS2xD(76)(4);
  CNStageIntLLRInputS3xD(332)(1) <= VNStageIntLLROutputS2xD(76)(5);
  CNStageIntLLRInputS3xD(348)(1) <= VNStageIntLLROutputS2xD(76)(6);
  CNStageIntLLRInputS3xD(119)(1) <= VNStageIntLLROutputS2xD(77)(0);
  CNStageIntLLRInputS3xD(185)(1) <= VNStageIntLLROutputS2xD(77)(1);
  CNStageIntLLRInputS3xD(257)(1) <= VNStageIntLLROutputS2xD(77)(2);
  CNStageIntLLRInputS3xD(293)(1) <= VNStageIntLLROutputS2xD(77)(3);
  CNStageIntLLRInputS3xD(383)(1) <= VNStageIntLLROutputS2xD(77)(4);
  CNStageIntLLRInputS3xD(40)(1) <= VNStageIntLLROutputS2xD(78)(0);
  CNStageIntLLRInputS3xD(84)(1) <= VNStageIntLLROutputS2xD(78)(1);
  CNStageIntLLRInputS3xD(159)(1) <= VNStageIntLLROutputS2xD(78)(2);
  CNStageIntLLRInputS3xD(193)(1) <= VNStageIntLLROutputS2xD(78)(3);
  CNStageIntLLRInputS3xD(274)(1) <= VNStageIntLLROutputS2xD(78)(4);
  CNStageIntLLRInputS3xD(288)(1) <= VNStageIntLLROutputS2xD(78)(5);
  CNStageIntLLRInputS3xD(374)(1) <= VNStageIntLLROutputS2xD(78)(6);
  CNStageIntLLRInputS3xD(39)(1) <= VNStageIntLLROutputS2xD(79)(0);
  CNStageIntLLRInputS3xD(99)(1) <= VNStageIntLLROutputS2xD(79)(1);
  CNStageIntLLRInputS3xD(167)(1) <= VNStageIntLLROutputS2xD(79)(2);
  CNStageIntLLRInputS3xD(220)(1) <= VNStageIntLLROutputS2xD(79)(3);
  CNStageIntLLRInputS3xD(325)(1) <= VNStageIntLLROutputS2xD(79)(4);
  CNStageIntLLRInputS3xD(38)(1) <= VNStageIntLLROutputS2xD(80)(0);
  CNStageIntLLRInputS3xD(62)(1) <= VNStageIntLLROutputS2xD(80)(1);
  CNStageIntLLRInputS3xD(131)(1) <= VNStageIntLLROutputS2xD(80)(2);
  CNStageIntLLRInputS3xD(182)(1) <= VNStageIntLLROutputS2xD(80)(3);
  CNStageIntLLRInputS3xD(248)(1) <= VNStageIntLLROutputS2xD(80)(4);
  CNStageIntLLRInputS3xD(337)(1) <= VNStageIntLLROutputS2xD(80)(5);
  CNStageIntLLRInputS3xD(37)(1) <= VNStageIntLLROutputS2xD(81)(0);
  CNStageIntLLRInputS3xD(72)(1) <= VNStageIntLLROutputS2xD(81)(1);
  CNStageIntLLRInputS3xD(129)(1) <= VNStageIntLLROutputS2xD(81)(2);
  CNStageIntLLRInputS3xD(262)(1) <= VNStageIntLLROutputS2xD(81)(3);
  CNStageIntLLRInputS3xD(36)(1) <= VNStageIntLLROutputS2xD(82)(0);
  CNStageIntLLRInputS3xD(67)(1) <= VNStageIntLLROutputS2xD(82)(1);
  CNStageIntLLRInputS3xD(165)(1) <= VNStageIntLLROutputS2xD(82)(2);
  CNStageIntLLRInputS3xD(188)(1) <= VNStageIntLLROutputS2xD(82)(3);
  CNStageIntLLRInputS3xD(254)(1) <= VNStageIntLLROutputS2xD(82)(4);
  CNStageIntLLRInputS3xD(298)(1) <= VNStageIntLLROutputS2xD(82)(5);
  CNStageIntLLRInputS3xD(336)(1) <= VNStageIntLLROutputS2xD(82)(6);
  CNStageIntLLRInputS3xD(35)(1) <= VNStageIntLLROutputS2xD(83)(0);
  CNStageIntLLRInputS3xD(73)(1) <= VNStageIntLLROutputS2xD(83)(1);
  CNStageIntLLRInputS3xD(144)(1) <= VNStageIntLLROutputS2xD(83)(2);
  CNStageIntLLRInputS3xD(208)(1) <= VNStageIntLLROutputS2xD(83)(3);
  CNStageIntLLRInputS3xD(232)(1) <= VNStageIntLLROutputS2xD(83)(4);
  CNStageIntLLRInputS3xD(330)(1) <= VNStageIntLLROutputS2xD(83)(5);
  CNStageIntLLRInputS3xD(34)(1) <= VNStageIntLLROutputS2xD(84)(0);
  CNStageIntLLRInputS3xD(61)(1) <= VNStageIntLLROutputS2xD(84)(1);
  CNStageIntLLRInputS3xD(147)(1) <= VNStageIntLLROutputS2xD(84)(2);
  CNStageIntLLRInputS3xD(222)(1) <= VNStageIntLLROutputS2xD(84)(3);
  CNStageIntLLRInputS3xD(310)(1) <= VNStageIntLLROutputS2xD(84)(4);
  CNStageIntLLRInputS3xD(371)(1) <= VNStageIntLLROutputS2xD(84)(5);
  CNStageIntLLRInputS3xD(33)(1) <= VNStageIntLLROutputS2xD(85)(0);
  CNStageIntLLRInputS3xD(132)(1) <= VNStageIntLLROutputS2xD(85)(1);
  CNStageIntLLRInputS3xD(218)(1) <= VNStageIntLLROutputS2xD(85)(2);
  CNStageIntLLRInputS3xD(235)(1) <= VNStageIntLLROutputS2xD(85)(3);
  CNStageIntLLRInputS3xD(313)(1) <= VNStageIntLLROutputS2xD(85)(4);
  CNStageIntLLRInputS3xD(379)(1) <= VNStageIntLLROutputS2xD(85)(5);
  CNStageIntLLRInputS3xD(32)(1) <= VNStageIntLLROutputS2xD(86)(0);
  CNStageIntLLRInputS3xD(166)(1) <= VNStageIntLLROutputS2xD(86)(1);
  CNStageIntLLRInputS3xD(239)(1) <= VNStageIntLLROutputS2xD(86)(2);
  CNStageIntLLRInputS3xD(343)(1) <= VNStageIntLLROutputS2xD(86)(3);
  CNStageIntLLRInputS3xD(31)(1) <= VNStageIntLLROutputS2xD(87)(0);
  CNStageIntLLRInputS3xD(77)(1) <= VNStageIntLLROutputS2xD(87)(1);
  CNStageIntLLRInputS3xD(128)(1) <= VNStageIntLLROutputS2xD(87)(2);
  CNStageIntLLRInputS3xD(203)(1) <= VNStageIntLLROutputS2xD(87)(3);
  CNStageIntLLRInputS3xD(229)(1) <= VNStageIntLLROutputS2xD(87)(4);
  CNStageIntLLRInputS3xD(331)(1) <= VNStageIntLLROutputS2xD(87)(5);
  CNStageIntLLRInputS3xD(341)(1) <= VNStageIntLLROutputS2xD(87)(6);
  CNStageIntLLRInputS3xD(30)(1) <= VNStageIntLLROutputS2xD(88)(0);
  CNStageIntLLRInputS3xD(79)(1) <= VNStageIntLLROutputS2xD(88)(1);
  CNStageIntLLRInputS3xD(156)(1) <= VNStageIntLLROutputS2xD(88)(2);
  CNStageIntLLRInputS3xD(204)(1) <= VNStageIntLLROutputS2xD(88)(3);
  CNStageIntLLRInputS3xD(263)(1) <= VNStageIntLLROutputS2xD(88)(4);
  CNStageIntLLRInputS3xD(297)(1) <= VNStageIntLLROutputS2xD(88)(5);
  CNStageIntLLRInputS3xD(377)(1) <= VNStageIntLLROutputS2xD(88)(6);
  CNStageIntLLRInputS3xD(29)(1) <= VNStageIntLLROutputS2xD(89)(0);
  CNStageIntLLRInputS3xD(102)(1) <= VNStageIntLLROutputS2xD(89)(1);
  CNStageIntLLRInputS3xD(140)(1) <= VNStageIntLLROutputS2xD(89)(2);
  CNStageIntLLRInputS3xD(184)(1) <= VNStageIntLLROutputS2xD(89)(3);
  CNStageIntLLRInputS3xD(247)(1) <= VNStageIntLLROutputS2xD(89)(4);
  CNStageIntLLRInputS3xD(355)(1) <= VNStageIntLLROutputS2xD(89)(5);
  CNStageIntLLRInputS3xD(28)(1) <= VNStageIntLLROutputS2xD(90)(0);
  CNStageIntLLRInputS3xD(85)(1) <= VNStageIntLLROutputS2xD(90)(1);
  CNStageIntLLRInputS3xD(168)(1) <= VNStageIntLLROutputS2xD(90)(2);
  CNStageIntLLRInputS3xD(175)(1) <= VNStageIntLLROutputS2xD(90)(3);
  CNStageIntLLRInputS3xD(258)(1) <= VNStageIntLLROutputS2xD(90)(4);
  CNStageIntLLRInputS3xD(307)(1) <= VNStageIntLLROutputS2xD(90)(5);
  CNStageIntLLRInputS3xD(358)(1) <= VNStageIntLLROutputS2xD(90)(6);
  CNStageIntLLRInputS3xD(27)(1) <= VNStageIntLLROutputS2xD(91)(0);
  CNStageIntLLRInputS3xD(96)(1) <= VNStageIntLLROutputS2xD(91)(1);
  CNStageIntLLRInputS3xD(158)(1) <= VNStageIntLLROutputS2xD(91)(2);
  CNStageIntLLRInputS3xD(191)(1) <= VNStageIntLLROutputS2xD(91)(3);
  CNStageIntLLRInputS3xD(269)(1) <= VNStageIntLLROutputS2xD(91)(4);
  CNStageIntLLRInputS3xD(280)(1) <= VNStageIntLLROutputS2xD(91)(5);
  CNStageIntLLRInputS3xD(344)(1) <= VNStageIntLLROutputS2xD(91)(6);
  CNStageIntLLRInputS3xD(26)(1) <= VNStageIntLLROutputS2xD(92)(0);
  CNStageIntLLRInputS3xD(103)(1) <= VNStageIntLLROutputS2xD(92)(1);
  CNStageIntLLRInputS3xD(145)(1) <= VNStageIntLLROutputS2xD(92)(2);
  CNStageIntLLRInputS3xD(195)(1) <= VNStageIntLLROutputS2xD(92)(3);
  CNStageIntLLRInputS3xD(242)(1) <= VNStageIntLLROutputS2xD(92)(4);
  CNStageIntLLRInputS3xD(324)(1) <= VNStageIntLLROutputS2xD(92)(5);
  CNStageIntLLRInputS3xD(378)(1) <= VNStageIntLLROutputS2xD(92)(6);
  CNStageIntLLRInputS3xD(25)(1) <= VNStageIntLLROutputS2xD(93)(0);
  CNStageIntLLRInputS3xD(78)(1) <= VNStageIntLLROutputS2xD(93)(1);
  CNStageIntLLRInputS3xD(164)(1) <= VNStageIntLLROutputS2xD(93)(2);
  CNStageIntLLRInputS3xD(224)(1) <= VNStageIntLLROutputS2xD(93)(3);
  CNStageIntLLRInputS3xD(231)(1) <= VNStageIntLLROutputS2xD(93)(4);
  CNStageIntLLRInputS3xD(311)(1) <= VNStageIntLLROutputS2xD(93)(5);
  CNStageIntLLRInputS3xD(340)(1) <= VNStageIntLLROutputS2xD(93)(6);
  CNStageIntLLRInputS3xD(24)(1) <= VNStageIntLLROutputS2xD(94)(0);
  CNStageIntLLRInputS3xD(92)(1) <= VNStageIntLLROutputS2xD(94)(1);
  CNStageIntLLRInputS3xD(194)(1) <= VNStageIntLLROutputS2xD(94)(2);
  CNStageIntLLRInputS3xD(329)(1) <= VNStageIntLLROutputS2xD(94)(3);
  CNStageIntLLRInputS3xD(368)(1) <= VNStageIntLLROutputS2xD(94)(4);
  CNStageIntLLRInputS3xD(23)(1) <= VNStageIntLLROutputS2xD(95)(0);
  CNStageIntLLRInputS3xD(63)(1) <= VNStageIntLLROutputS2xD(95)(1);
  CNStageIntLLRInputS3xD(134)(1) <= VNStageIntLLROutputS2xD(95)(2);
  CNStageIntLLRInputS3xD(190)(1) <= VNStageIntLLROutputS2xD(95)(3);
  CNStageIntLLRInputS3xD(234)(1) <= VNStageIntLLROutputS2xD(95)(4);
  CNStageIntLLRInputS3xD(303)(1) <= VNStageIntLLROutputS2xD(95)(5);
  CNStageIntLLRInputS3xD(352)(1) <= VNStageIntLLROutputS2xD(95)(6);
  CNStageIntLLRInputS3xD(22)(1) <= VNStageIntLLROutputS2xD(96)(0);
  CNStageIntLLRInputS3xD(98)(1) <= VNStageIntLLROutputS2xD(96)(1);
  CNStageIntLLRInputS3xD(150)(1) <= VNStageIntLLROutputS2xD(96)(2);
  CNStageIntLLRInputS3xD(172)(1) <= VNStageIntLLROutputS2xD(96)(3);
  CNStageIntLLRInputS3xD(251)(1) <= VNStageIntLLROutputS2xD(96)(4);
  CNStageIntLLRInputS3xD(380)(1) <= VNStageIntLLROutputS2xD(96)(5);
  CNStageIntLLRInputS3xD(21)(1) <= VNStageIntLLROutputS2xD(97)(0);
  CNStageIntLLRInputS3xD(65)(1) <= VNStageIntLLROutputS2xD(97)(1);
  CNStageIntLLRInputS3xD(142)(1) <= VNStageIntLLROutputS2xD(97)(2);
  CNStageIntLLRInputS3xD(180)(1) <= VNStageIntLLROutputS2xD(97)(3);
  CNStageIntLLRInputS3xD(260)(1) <= VNStageIntLLROutputS2xD(97)(4);
  CNStageIntLLRInputS3xD(316)(1) <= VNStageIntLLROutputS2xD(97)(5);
  CNStageIntLLRInputS3xD(370)(1) <= VNStageIntLLROutputS2xD(97)(6);
  CNStageIntLLRInputS3xD(20)(1) <= VNStageIntLLROutputS2xD(98)(0);
  CNStageIntLLRInputS3xD(116)(1) <= VNStageIntLLROutputS2xD(98)(1);
  CNStageIntLLRInputS3xD(199)(1) <= VNStageIntLLROutputS2xD(98)(2);
  CNStageIntLLRInputS3xD(255)(1) <= VNStageIntLLROutputS2xD(98)(3);
  CNStageIntLLRInputS3xD(308)(1) <= VNStageIntLLROutputS2xD(98)(4);
  CNStageIntLLRInputS3xD(356)(1) <= VNStageIntLLROutputS2xD(98)(5);
  CNStageIntLLRInputS3xD(19)(1) <= VNStageIntLLROutputS2xD(99)(0);
  CNStageIntLLRInputS3xD(76)(1) <= VNStageIntLLROutputS2xD(99)(1);
  CNStageIntLLRInputS3xD(126)(1) <= VNStageIntLLROutputS2xD(99)(2);
  CNStageIntLLRInputS3xD(198)(1) <= VNStageIntLLROutputS2xD(99)(3);
  CNStageIntLLRInputS3xD(261)(1) <= VNStageIntLLROutputS2xD(99)(4);
  CNStageIntLLRInputS3xD(285)(1) <= VNStageIntLLROutputS2xD(99)(5);
  CNStageIntLLRInputS3xD(376)(1) <= VNStageIntLLROutputS2xD(99)(6);
  CNStageIntLLRInputS3xD(18)(1) <= VNStageIntLLROutputS2xD(100)(0);
  CNStageIntLLRInputS3xD(94)(1) <= VNStageIntLLROutputS2xD(100)(1);
  CNStageIntLLRInputS3xD(120)(1) <= VNStageIntLLROutputS2xD(100)(2);
  CNStageIntLLRInputS3xD(178)(1) <= VNStageIntLLROutputS2xD(100)(3);
  CNStageIntLLRInputS3xD(250)(1) <= VNStageIntLLROutputS2xD(100)(4);
  CNStageIntLLRInputS3xD(295)(1) <= VNStageIntLLROutputS2xD(100)(5);
  CNStageIntLLRInputS3xD(349)(1) <= VNStageIntLLROutputS2xD(100)(6);
  CNStageIntLLRInputS3xD(17)(1) <= VNStageIntLLROutputS2xD(101)(0);
  CNStageIntLLRInputS3xD(58)(1) <= VNStageIntLLROutputS2xD(101)(1);
  CNStageIntLLRInputS3xD(123)(1) <= VNStageIntLLROutputS2xD(101)(2);
  CNStageIntLLRInputS3xD(211)(1) <= VNStageIntLLROutputS2xD(101)(3);
  CNStageIntLLRInputS3xD(273)(1) <= VNStageIntLLROutputS2xD(101)(4);
  CNStageIntLLRInputS3xD(289)(1) <= VNStageIntLLROutputS2xD(101)(5);
  CNStageIntLLRInputS3xD(346)(1) <= VNStageIntLLROutputS2xD(101)(6);
  CNStageIntLLRInputS3xD(16)(1) <= VNStageIntLLROutputS2xD(102)(0);
  CNStageIntLLRInputS3xD(59)(1) <= VNStageIntLLROutputS2xD(102)(1);
  CNStageIntLLRInputS3xD(113)(1) <= VNStageIntLLROutputS2xD(102)(2);
  CNStageIntLLRInputS3xD(214)(1) <= VNStageIntLLROutputS2xD(102)(3);
  CNStageIntLLRInputS3xD(226)(1) <= VNStageIntLLROutputS2xD(102)(4);
  CNStageIntLLRInputS3xD(361)(1) <= VNStageIntLLROutputS2xD(102)(5);
  CNStageIntLLRInputS3xD(15)(1) <= VNStageIntLLROutputS2xD(103)(0);
  CNStageIntLLRInputS3xD(93)(1) <= VNStageIntLLROutputS2xD(103)(1);
  CNStageIntLLRInputS3xD(151)(1) <= VNStageIntLLROutputS2xD(103)(2);
  CNStageIntLLRInputS3xD(200)(1) <= VNStageIntLLROutputS2xD(103)(3);
  CNStageIntLLRInputS3xD(265)(1) <= VNStageIntLLROutputS2xD(103)(4);
  CNStageIntLLRInputS3xD(284)(1) <= VNStageIntLLROutputS2xD(103)(5);
  CNStageIntLLRInputS3xD(354)(1) <= VNStageIntLLROutputS2xD(103)(6);
  CNStageIntLLRInputS3xD(14)(1) <= VNStageIntLLROutputS2xD(104)(0);
  CNStageIntLLRInputS3xD(86)(1) <= VNStageIntLLROutputS2xD(104)(1);
  CNStageIntLLRInputS3xD(133)(1) <= VNStageIntLLROutputS2xD(104)(2);
  CNStageIntLLRInputS3xD(179)(1) <= VNStageIntLLROutputS2xD(104)(3);
  CNStageIntLLRInputS3xD(267)(1) <= VNStageIntLLROutputS2xD(104)(4);
  CNStageIntLLRInputS3xD(317)(1) <= VNStageIntLLROutputS2xD(104)(5);
  CNStageIntLLRInputS3xD(13)(1) <= VNStageIntLLROutputS2xD(105)(0);
  CNStageIntLLRInputS3xD(146)(1) <= VNStageIntLLROutputS2xD(105)(1);
  CNStageIntLLRInputS3xD(197)(1) <= VNStageIntLLROutputS2xD(105)(2);
  CNStageIntLLRInputS3xD(237)(1) <= VNStageIntLLROutputS2xD(105)(3);
  CNStageIntLLRInputS3xD(300)(1) <= VNStageIntLLROutputS2xD(105)(4);
  CNStageIntLLRInputS3xD(338)(1) <= VNStageIntLLROutputS2xD(105)(5);
  CNStageIntLLRInputS3xD(12)(1) <= VNStageIntLLROutputS2xD(106)(0);
  CNStageIntLLRInputS3xD(157)(1) <= VNStageIntLLROutputS2xD(106)(1);
  CNStageIntLLRInputS3xD(223)(1) <= VNStageIntLLROutputS2xD(106)(2);
  CNStageIntLLRInputS3xD(272)(1) <= VNStageIntLLROutputS2xD(106)(3);
  CNStageIntLLRInputS3xD(312)(1) <= VNStageIntLLROutputS2xD(106)(4);
  CNStageIntLLRInputS3xD(333)(1) <= VNStageIntLLROutputS2xD(106)(5);
  CNStageIntLLRInputS3xD(110)(1) <= VNStageIntLLROutputS2xD(107)(0);
  CNStageIntLLRInputS3xD(127)(1) <= VNStageIntLLROutputS2xD(107)(1);
  CNStageIntLLRInputS3xD(207)(1) <= VNStageIntLLROutputS2xD(107)(2);
  CNStageIntLLRInputS3xD(230)(1) <= VNStageIntLLROutputS2xD(107)(3);
  CNStageIntLLRInputS3xD(323)(1) <= VNStageIntLLROutputS2xD(107)(4);
  CNStageIntLLRInputS3xD(335)(1) <= VNStageIntLLROutputS2xD(107)(5);
  CNStageIntLLRInputS3xD(11)(1) <= VNStageIntLLROutputS2xD(108)(0);
  CNStageIntLLRInputS3xD(105)(1) <= VNStageIntLLROutputS2xD(108)(1);
  CNStageIntLLRInputS3xD(115)(1) <= VNStageIntLLROutputS2xD(108)(2);
  CNStageIntLLRInputS3xD(181)(1) <= VNStageIntLLROutputS2xD(108)(3);
  CNStageIntLLRInputS3xD(238)(1) <= VNStageIntLLROutputS2xD(108)(4);
  CNStageIntLLRInputS3xD(296)(1) <= VNStageIntLLROutputS2xD(108)(5);
  CNStageIntLLRInputS3xD(10)(1) <= VNStageIntLLROutputS2xD(109)(0);
  CNStageIntLLRInputS3xD(100)(1) <= VNStageIntLLROutputS2xD(109)(1);
  CNStageIntLLRInputS3xD(160)(1) <= VNStageIntLLROutputS2xD(109)(2);
  CNStageIntLLRInputS3xD(171)(1) <= VNStageIntLLROutputS2xD(109)(3);
  CNStageIntLLRInputS3xD(266)(1) <= VNStageIntLLROutputS2xD(109)(4);
  CNStageIntLLRInputS3xD(362)(1) <= VNStageIntLLROutputS2xD(109)(5);
  CNStageIntLLRInputS3xD(9)(1) <= VNStageIntLLROutputS2xD(110)(0);
  CNStageIntLLRInputS3xD(83)(1) <= VNStageIntLLROutputS2xD(110)(1);
  CNStageIntLLRInputS3xD(118)(1) <= VNStageIntLLROutputS2xD(110)(2);
  CNStageIntLLRInputS3xD(212)(1) <= VNStageIntLLROutputS2xD(110)(3);
  CNStageIntLLRInputS3xD(225)(1) <= VNStageIntLLROutputS2xD(110)(4);
  CNStageIntLLRInputS3xD(326)(1) <= VNStageIntLLROutputS2xD(110)(5);
  CNStageIntLLRInputS3xD(345)(1) <= VNStageIntLLROutputS2xD(110)(6);
  CNStageIntLLRInputS3xD(8)(1) <= VNStageIntLLROutputS2xD(111)(0);
  CNStageIntLLRInputS3xD(90)(1) <= VNStageIntLLROutputS2xD(111)(1);
  CNStageIntLLRInputS3xD(138)(1) <= VNStageIntLLROutputS2xD(111)(2);
  CNStageIntLLRInputS3xD(177)(1) <= VNStageIntLLROutputS2xD(111)(3);
  CNStageIntLLRInputS3xD(252)(1) <= VNStageIntLLROutputS2xD(111)(4);
  CNStageIntLLRInputS3xD(287)(1) <= VNStageIntLLROutputS2xD(111)(5);
  CNStageIntLLRInputS3xD(357)(1) <= VNStageIntLLROutputS2xD(111)(6);
  CNStageIntLLRInputS3xD(7)(1) <= VNStageIntLLROutputS2xD(112)(0);
  CNStageIntLLRInputS3xD(54)(1) <= VNStageIntLLROutputS2xD(112)(1);
  CNStageIntLLRInputS3xD(148)(1) <= VNStageIntLLROutputS2xD(112)(2);
  CNStageIntLLRInputS3xD(205)(1) <= VNStageIntLLROutputS2xD(112)(3);
  CNStageIntLLRInputS3xD(233)(1) <= VNStageIntLLROutputS2xD(112)(4);
  CNStageIntLLRInputS3xD(305)(1) <= VNStageIntLLROutputS2xD(112)(5);
  CNStageIntLLRInputS3xD(369)(1) <= VNStageIntLLROutputS2xD(112)(6);
  CNStageIntLLRInputS3xD(6)(1) <= VNStageIntLLROutputS2xD(113)(0);
  CNStageIntLLRInputS3xD(108)(1) <= VNStageIntLLROutputS2xD(113)(1);
  CNStageIntLLRInputS3xD(143)(1) <= VNStageIntLLROutputS2xD(113)(2);
  CNStageIntLLRInputS3xD(202)(1) <= VNStageIntLLROutputS2xD(113)(3);
  CNStageIntLLRInputS3xD(253)(1) <= VNStageIntLLROutputS2xD(113)(4);
  CNStageIntLLRInputS3xD(314)(1) <= VNStageIntLLROutputS2xD(113)(5);
  CNStageIntLLRInputS3xD(339)(1) <= VNStageIntLLROutputS2xD(113)(6);
  CNStageIntLLRInputS3xD(5)(1) <= VNStageIntLLROutputS2xD(114)(0);
  CNStageIntLLRInputS3xD(88)(1) <= VNStageIntLLROutputS2xD(114)(1);
  CNStageIntLLRInputS3xD(149)(1) <= VNStageIntLLROutputS2xD(114)(2);
  CNStageIntLLRInputS3xD(216)(1) <= VNStageIntLLROutputS2xD(114)(3);
  CNStageIntLLRInputS3xD(268)(1) <= VNStageIntLLROutputS2xD(114)(4);
  CNStageIntLLRInputS3xD(309)(1) <= VNStageIntLLROutputS2xD(114)(5);
  CNStageIntLLRInputS3xD(4)(1) <= VNStageIntLLROutputS2xD(115)(0);
  CNStageIntLLRInputS3xD(68)(1) <= VNStageIntLLROutputS2xD(115)(1);
  CNStageIntLLRInputS3xD(137)(1) <= VNStageIntLLROutputS2xD(115)(2);
  CNStageIntLLRInputS3xD(209)(1) <= VNStageIntLLROutputS2xD(115)(3);
  CNStageIntLLRInputS3xD(264)(1) <= VNStageIntLLROutputS2xD(115)(4);
  CNStageIntLLRInputS3xD(315)(1) <= VNStageIntLLROutputS2xD(115)(5);
  CNStageIntLLRInputS3xD(372)(1) <= VNStageIntLLROutputS2xD(115)(6);
  CNStageIntLLRInputS3xD(71)(1) <= VNStageIntLLROutputS2xD(116)(0);
  CNStageIntLLRInputS3xD(163)(1) <= VNStageIntLLROutputS2xD(116)(1);
  CNStageIntLLRInputS3xD(187)(1) <= VNStageIntLLROutputS2xD(116)(2);
  CNStageIntLLRInputS3xD(228)(1) <= VNStageIntLLROutputS2xD(116)(3);
  CNStageIntLLRInputS3xD(304)(1) <= VNStageIntLLROutputS2xD(116)(4);
  CNStageIntLLRInputS3xD(3)(1) <= VNStageIntLLROutputS2xD(117)(0);
  CNStageIntLLRInputS3xD(55)(1) <= VNStageIntLLROutputS2xD(117)(1);
  CNStageIntLLRInputS3xD(111)(1) <= VNStageIntLLROutputS2xD(117)(2);
  CNStageIntLLRInputS3xD(196)(1) <= VNStageIntLLROutputS2xD(117)(3);
  CNStageIntLLRInputS3xD(2)(1) <= VNStageIntLLROutputS2xD(118)(0);
  CNStageIntLLRInputS3xD(89)(1) <= VNStageIntLLROutputS2xD(118)(1);
  CNStageIntLLRInputS3xD(152)(1) <= VNStageIntLLROutputS2xD(118)(2);
  CNStageIntLLRInputS3xD(249)(1) <= VNStageIntLLROutputS2xD(118)(3);
  CNStageIntLLRInputS3xD(282)(1) <= VNStageIntLLROutputS2xD(118)(4);
  CNStageIntLLRInputS3xD(359)(1) <= VNStageIntLLROutputS2xD(118)(5);
  CNStageIntLLRInputS3xD(1)(1) <= VNStageIntLLROutputS2xD(119)(0);
  CNStageIntLLRInputS3xD(107)(1) <= VNStageIntLLROutputS2xD(119)(1);
  CNStageIntLLRInputS3xD(154)(1) <= VNStageIntLLROutputS2xD(119)(2);
  CNStageIntLLRInputS3xD(227)(1) <= VNStageIntLLROutputS2xD(119)(3);
  CNStageIntLLRInputS3xD(319)(1) <= VNStageIntLLROutputS2xD(119)(4);
  CNStageIntLLRInputS3xD(0)(1) <= VNStageIntLLROutputS2xD(120)(0);
  CNStageIntLLRInputS3xD(80)(1) <= VNStageIntLLROutputS2xD(120)(1);
  CNStageIntLLRInputS3xD(321)(1) <= VNStageIntLLROutputS2xD(120)(2);
  CNStageIntLLRInputS3xD(360)(1) <= VNStageIntLLROutputS2xD(120)(3);
  CNStageIntLLRInputS3xD(64)(1) <= VNStageIntLLROutputS2xD(121)(0);
  CNStageIntLLRInputS3xD(161)(1) <= VNStageIntLLROutputS2xD(121)(1);
  CNStageIntLLRInputS3xD(217)(1) <= VNStageIntLLROutputS2xD(121)(2);
  CNStageIntLLRInputS3xD(236)(1) <= VNStageIntLLROutputS2xD(121)(3);
  CNStageIntLLRInputS3xD(291)(1) <= VNStageIntLLROutputS2xD(121)(4);
  CNStageIntLLRInputS3xD(350)(1) <= VNStageIntLLROutputS2xD(121)(5);
  CNStageIntLLRInputS3xD(91)(1) <= VNStageIntLLROutputS2xD(122)(0);
  CNStageIntLLRInputS3xD(114)(1) <= VNStageIntLLROutputS2xD(122)(1);
  CNStageIntLLRInputS3xD(201)(1) <= VNStageIntLLROutputS2xD(122)(2);
  CNStageIntLLRInputS3xD(241)(1) <= VNStageIntLLROutputS2xD(122)(3);
  CNStageIntLLRInputS3xD(327)(1) <= VNStageIntLLROutputS2xD(122)(4);
  CNStageIntLLRInputS3xD(375)(1) <= VNStageIntLLROutputS2xD(122)(5);
  CNStageIntLLRInputS3xD(82)(1) <= VNStageIntLLROutputS2xD(123)(0);
  CNStageIntLLRInputS3xD(122)(1) <= VNStageIntLLROutputS2xD(123)(1);
  CNStageIntLLRInputS3xD(213)(1) <= VNStageIntLLROutputS2xD(123)(2);
  CNStageIntLLRInputS3xD(279)(1) <= VNStageIntLLROutputS2xD(123)(3);
  CNStageIntLLRInputS3xD(382)(1) <= VNStageIntLLROutputS2xD(123)(4);
  CNStageIntLLRInputS3xD(69)(1) <= VNStageIntLLROutputS2xD(124)(0);
  CNStageIntLLRInputS3xD(153)(1) <= VNStageIntLLROutputS2xD(124)(1);
  CNStageIntLLRInputS3xD(240)(1) <= VNStageIntLLROutputS2xD(124)(2);
  CNStageIntLLRInputS3xD(292)(1) <= VNStageIntLLROutputS2xD(124)(3);
  CNStageIntLLRInputS3xD(364)(1) <= VNStageIntLLROutputS2xD(124)(4);
  CNStageIntLLRInputS3xD(87)(1) <= VNStageIntLLROutputS2xD(125)(0);
  CNStageIntLLRInputS3xD(169)(1) <= VNStageIntLLROutputS2xD(125)(1);
  CNStageIntLLRInputS3xD(320)(1) <= VNStageIntLLROutputS2xD(125)(2);
  CNStageIntLLRInputS3xD(366)(1) <= VNStageIntLLROutputS2xD(125)(3);
  CNStageIntLLRInputS3xD(60)(1) <= VNStageIntLLROutputS2xD(126)(0);
  CNStageIntLLRInputS3xD(139)(1) <= VNStageIntLLROutputS2xD(126)(1);
  CNStageIntLLRInputS3xD(186)(1) <= VNStageIntLLROutputS2xD(126)(2);
  CNStageIntLLRInputS3xD(271)(1) <= VNStageIntLLROutputS2xD(126)(3);
  CNStageIntLLRInputS3xD(281)(1) <= VNStageIntLLROutputS2xD(126)(4);
  CNStageIntLLRInputS3xD(334)(1) <= VNStageIntLLROutputS2xD(126)(5);
  CNStageIntLLRInputS3xD(52)(1) <= VNStageIntLLROutputS2xD(127)(0);
  CNStageIntLLRInputS3xD(57)(1) <= VNStageIntLLROutputS2xD(127)(1);
  CNStageIntLLRInputS3xD(117)(1) <= VNStageIntLLROutputS2xD(127)(2);
  CNStageIntLLRInputS3xD(173)(1) <= VNStageIntLLROutputS2xD(127)(3);
  CNStageIntLLRInputS3xD(277)(1) <= VNStageIntLLROutputS2xD(127)(4);
  CNStageIntLLRInputS3xD(306)(1) <= VNStageIntLLROutputS2xD(127)(5);
  CNStageIntLLRInputS3xD(373)(1) <= VNStageIntLLROutputS2xD(127)(6);
  CNStageIntLLRInputS3xD(53)(2) <= VNStageIntLLROutputS2xD(128)(0);
  CNStageIntLLRInputS3xD(108)(2) <= VNStageIntLLROutputS2xD(128)(1);
  CNStageIntLLRInputS3xD(129)(2) <= VNStageIntLLROutputS2xD(128)(2);
  CNStageIntLLRInputS3xD(198)(2) <= VNStageIntLLROutputS2xD(128)(3);
  CNStageIntLLRInputS3xD(244)(2) <= VNStageIntLLROutputS2xD(128)(4);
  CNStageIntLLRInputS3xD(298)(2) <= VNStageIntLLROutputS2xD(128)(5);
  CNStageIntLLRInputS3xD(341)(2) <= VNStageIntLLROutputS2xD(128)(6);
  CNStageIntLLRInputS3xD(51)(2) <= VNStageIntLLROutputS2xD(129)(0);
  CNStageIntLLRInputS3xD(56)(2) <= VNStageIntLLROutputS2xD(129)(1);
  CNStageIntLLRInputS3xD(116)(2) <= VNStageIntLLROutputS2xD(129)(2);
  CNStageIntLLRInputS3xD(172)(2) <= VNStageIntLLROutputS2xD(129)(3);
  CNStageIntLLRInputS3xD(276)(2) <= VNStageIntLLROutputS2xD(129)(4);
  CNStageIntLLRInputS3xD(305)(2) <= VNStageIntLLROutputS2xD(129)(5);
  CNStageIntLLRInputS3xD(372)(2) <= VNStageIntLLROutputS2xD(129)(6);
  CNStageIntLLRInputS3xD(50)(2) <= VNStageIntLLROutputS2xD(130)(0);
  CNStageIntLLRInputS3xD(73)(2) <= VNStageIntLLROutputS2xD(130)(1);
  CNStageIntLLRInputS3xD(140)(2) <= VNStageIntLLROutputS2xD(130)(2);
  CNStageIntLLRInputS3xD(188)(2) <= VNStageIntLLROutputS2xD(130)(3);
  CNStageIntLLRInputS3xD(245)(2) <= VNStageIntLLROutputS2xD(130)(4);
  CNStageIntLLRInputS3xD(285)(2) <= VNStageIntLLROutputS2xD(130)(5);
  CNStageIntLLRInputS3xD(65)(2) <= VNStageIntLLROutputS2xD(131)(0);
  CNStageIntLLRInputS3xD(154)(2) <= VNStageIntLLROutputS2xD(131)(1);
  CNStageIntLLRInputS3xD(206)(2) <= VNStageIntLLROutputS2xD(131)(2);
  CNStageIntLLRInputS3xD(243)(2) <= VNStageIntLLROutputS2xD(131)(3);
  CNStageIntLLRInputS3xD(307)(2) <= VNStageIntLLROutputS2xD(131)(4);
  CNStageIntLLRInputS3xD(334)(2) <= VNStageIntLLROutputS2xD(131)(5);
  CNStageIntLLRInputS3xD(49)(2) <= VNStageIntLLROutputS2xD(132)(0);
  CNStageIntLLRInputS3xD(151)(2) <= VNStageIntLLROutputS2xD(132)(1);
  CNStageIntLLRInputS3xD(214)(2) <= VNStageIntLLROutputS2xD(132)(2);
  CNStageIntLLRInputS3xD(274)(2) <= VNStageIntLLROutputS2xD(132)(3);
  CNStageIntLLRInputS3xD(321)(2) <= VNStageIntLLROutputS2xD(132)(4);
  CNStageIntLLRInputS3xD(364)(2) <= VNStageIntLLROutputS2xD(132)(5);
  CNStageIntLLRInputS3xD(48)(2) <= VNStageIntLLROutputS2xD(133)(0);
  CNStageIntLLRInputS3xD(209)(2) <= VNStageIntLLROutputS2xD(133)(1);
  CNStageIntLLRInputS3xD(255)(2) <= VNStageIntLLROutputS2xD(133)(2);
  CNStageIntLLRInputS3xD(317)(2) <= VNStageIntLLROutputS2xD(133)(3);
  CNStageIntLLRInputS3xD(380)(2) <= VNStageIntLLROutputS2xD(133)(4);
  CNStageIntLLRInputS3xD(47)(2) <= VNStageIntLLROutputS2xD(134)(0);
  CNStageIntLLRInputS3xD(100)(2) <= VNStageIntLLROutputS2xD(134)(1);
  CNStageIntLLRInputS3xD(134)(2) <= VNStageIntLLROutputS2xD(134)(2);
  CNStageIntLLRInputS3xD(258)(2) <= VNStageIntLLROutputS2xD(134)(3);
  CNStageIntLLRInputS3xD(46)(2) <= VNStageIntLLROutputS2xD(135)(0);
  CNStageIntLLRInputS3xD(103)(2) <= VNStageIntLLROutputS2xD(135)(1);
  CNStageIntLLRInputS3xD(135)(2) <= VNStageIntLLROutputS2xD(135)(2);
  CNStageIntLLRInputS3xD(205)(2) <= VNStageIntLLROutputS2xD(135)(3);
  CNStageIntLLRInputS3xD(45)(2) <= VNStageIntLLROutputS2xD(136)(0);
  CNStageIntLLRInputS3xD(94)(2) <= VNStageIntLLROutputS2xD(136)(1);
  CNStageIntLLRInputS3xD(111)(2) <= VNStageIntLLROutputS2xD(136)(2);
  CNStageIntLLRInputS3xD(175)(2) <= VNStageIntLLROutputS2xD(136)(3);
  CNStageIntLLRInputS3xD(275)(2) <= VNStageIntLLROutputS2xD(136)(4);
  CNStageIntLLRInputS3xD(301)(2) <= VNStageIntLLROutputS2xD(136)(5);
  CNStageIntLLRInputS3xD(352)(2) <= VNStageIntLLROutputS2xD(136)(6);
  CNStageIntLLRInputS3xD(44)(2) <= VNStageIntLLROutputS2xD(137)(0);
  CNStageIntLLRInputS3xD(74)(2) <= VNStageIntLLROutputS2xD(137)(1);
  CNStageIntLLRInputS3xD(161)(2) <= VNStageIntLLROutputS2xD(137)(2);
  CNStageIntLLRInputS3xD(182)(2) <= VNStageIntLLROutputS2xD(137)(3);
  CNStageIntLLRInputS3xD(242)(2) <= VNStageIntLLROutputS2xD(137)(4);
  CNStageIntLLRInputS3xD(282)(2) <= VNStageIntLLROutputS2xD(137)(5);
  CNStageIntLLRInputS3xD(366)(2) <= VNStageIntLLROutputS2xD(137)(6);
  CNStageIntLLRInputS3xD(43)(2) <= VNStageIntLLROutputS2xD(138)(0);
  CNStageIntLLRInputS3xD(55)(2) <= VNStageIntLLROutputS2xD(138)(1);
  CNStageIntLLRInputS3xD(120)(2) <= VNStageIntLLROutputS2xD(138)(2);
  CNStageIntLLRInputS3xD(218)(2) <= VNStageIntLLROutputS2xD(138)(3);
  CNStageIntLLRInputS3xD(268)(2) <= VNStageIntLLROutputS2xD(138)(4);
  CNStageIntLLRInputS3xD(327)(2) <= VNStageIntLLROutputS2xD(138)(5);
  CNStageIntLLRInputS3xD(362)(2) <= VNStageIntLLROutputS2xD(138)(6);
  CNStageIntLLRInputS3xD(42)(2) <= VNStageIntLLROutputS2xD(139)(0);
  CNStageIntLLRInputS3xD(69)(2) <= VNStageIntLLROutputS2xD(139)(1);
  CNStageIntLLRInputS3xD(124)(2) <= VNStageIntLLROutputS2xD(139)(2);
  CNStageIntLLRInputS3xD(220)(2) <= VNStageIntLLROutputS2xD(139)(3);
  CNStageIntLLRInputS3xD(252)(2) <= VNStageIntLLROutputS2xD(139)(4);
  CNStageIntLLRInputS3xD(289)(2) <= VNStageIntLLROutputS2xD(139)(5);
  CNStageIntLLRInputS3xD(383)(2) <= VNStageIntLLROutputS2xD(139)(6);
  CNStageIntLLRInputS3xD(41)(2) <= VNStageIntLLROutputS2xD(140)(0);
  CNStageIntLLRInputS3xD(80)(2) <= VNStageIntLLROutputS2xD(140)(1);
  CNStageIntLLRInputS3xD(170)(2) <= VNStageIntLLROutputS2xD(140)(2);
  CNStageIntLLRInputS3xD(191)(2) <= VNStageIntLLROutputS2xD(140)(3);
  CNStageIntLLRInputS3xD(277)(2) <= VNStageIntLLROutputS2xD(140)(4);
  CNStageIntLLRInputS3xD(293)(2) <= VNStageIntLLROutputS2xD(140)(5);
  CNStageIntLLRInputS3xD(346)(2) <= VNStageIntLLROutputS2xD(140)(6);
  CNStageIntLLRInputS3xD(123)(2) <= VNStageIntLLROutputS2xD(141)(0);
  CNStageIntLLRInputS3xD(173)(2) <= VNStageIntLLROutputS2xD(141)(1);
  CNStageIntLLRInputS3xD(269)(2) <= VNStageIntLLROutputS2xD(141)(2);
  CNStageIntLLRInputS3xD(332)(2) <= VNStageIntLLROutputS2xD(141)(3);
  CNStageIntLLRInputS3xD(347)(2) <= VNStageIntLLROutputS2xD(141)(4);
  CNStageIntLLRInputS3xD(40)(2) <= VNStageIntLLROutputS2xD(142)(0);
  CNStageIntLLRInputS3xD(96)(2) <= VNStageIntLLROutputS2xD(142)(1);
  CNStageIntLLRInputS3xD(118)(2) <= VNStageIntLLROutputS2xD(142)(2);
  CNStageIntLLRInputS3xD(256)(2) <= VNStageIntLLROutputS2xD(142)(3);
  CNStageIntLLRInputS3xD(382)(2) <= VNStageIntLLROutputS2xD(142)(4);
  CNStageIntLLRInputS3xD(39)(2) <= VNStageIntLLROutputS2xD(143)(0);
  CNStageIntLLRInputS3xD(83)(2) <= VNStageIntLLROutputS2xD(143)(1);
  CNStageIntLLRInputS3xD(158)(2) <= VNStageIntLLROutputS2xD(143)(2);
  CNStageIntLLRInputS3xD(192)(2) <= VNStageIntLLROutputS2xD(143)(3);
  CNStageIntLLRInputS3xD(273)(2) <= VNStageIntLLROutputS2xD(143)(4);
  CNStageIntLLRInputS3xD(287)(2) <= VNStageIntLLROutputS2xD(143)(5);
  CNStageIntLLRInputS3xD(373)(2) <= VNStageIntLLROutputS2xD(143)(6);
  CNStageIntLLRInputS3xD(38)(2) <= VNStageIntLLROutputS2xD(144)(0);
  CNStageIntLLRInputS3xD(98)(2) <= VNStageIntLLROutputS2xD(144)(1);
  CNStageIntLLRInputS3xD(166)(2) <= VNStageIntLLROutputS2xD(144)(2);
  CNStageIntLLRInputS3xD(219)(2) <= VNStageIntLLROutputS2xD(144)(3);
  CNStageIntLLRInputS3xD(249)(2) <= VNStageIntLLROutputS2xD(144)(4);
  CNStageIntLLRInputS3xD(324)(2) <= VNStageIntLLROutputS2xD(144)(5);
  CNStageIntLLRInputS3xD(333)(2) <= VNStageIntLLROutputS2xD(144)(6);
  CNStageIntLLRInputS3xD(37)(2) <= VNStageIntLLROutputS2xD(145)(0);
  CNStageIntLLRInputS3xD(61)(2) <= VNStageIntLLROutputS2xD(145)(1);
  CNStageIntLLRInputS3xD(130)(2) <= VNStageIntLLROutputS2xD(145)(2);
  CNStageIntLLRInputS3xD(181)(2) <= VNStageIntLLROutputS2xD(145)(3);
  CNStageIntLLRInputS3xD(247)(2) <= VNStageIntLLROutputS2xD(145)(4);
  CNStageIntLLRInputS3xD(331)(2) <= VNStageIntLLROutputS2xD(145)(5);
  CNStageIntLLRInputS3xD(336)(2) <= VNStageIntLLROutputS2xD(145)(6);
  CNStageIntLLRInputS3xD(36)(2) <= VNStageIntLLROutputS2xD(146)(0);
  CNStageIntLLRInputS3xD(71)(2) <= VNStageIntLLROutputS2xD(146)(1);
  CNStageIntLLRInputS3xD(128)(2) <= VNStageIntLLROutputS2xD(146)(2);
  CNStageIntLLRInputS3xD(261)(2) <= VNStageIntLLROutputS2xD(146)(3);
  CNStageIntLLRInputS3xD(299)(2) <= VNStageIntLLROutputS2xD(146)(4);
  CNStageIntLLRInputS3xD(35)(2) <= VNStageIntLLROutputS2xD(147)(0);
  CNStageIntLLRInputS3xD(66)(2) <= VNStageIntLLROutputS2xD(147)(1);
  CNStageIntLLRInputS3xD(164)(2) <= VNStageIntLLROutputS2xD(147)(2);
  CNStageIntLLRInputS3xD(187)(2) <= VNStageIntLLROutputS2xD(147)(3);
  CNStageIntLLRInputS3xD(253)(2) <= VNStageIntLLROutputS2xD(147)(4);
  CNStageIntLLRInputS3xD(297)(2) <= VNStageIntLLROutputS2xD(147)(5);
  CNStageIntLLRInputS3xD(335)(2) <= VNStageIntLLROutputS2xD(147)(6);
  CNStageIntLLRInputS3xD(34)(2) <= VNStageIntLLROutputS2xD(148)(0);
  CNStageIntLLRInputS3xD(72)(2) <= VNStageIntLLROutputS2xD(148)(1);
  CNStageIntLLRInputS3xD(143)(2) <= VNStageIntLLROutputS2xD(148)(2);
  CNStageIntLLRInputS3xD(207)(2) <= VNStageIntLLROutputS2xD(148)(3);
  CNStageIntLLRInputS3xD(231)(2) <= VNStageIntLLROutputS2xD(148)(4);
  CNStageIntLLRInputS3xD(329)(2) <= VNStageIntLLROutputS2xD(148)(5);
  CNStageIntLLRInputS3xD(33)(2) <= VNStageIntLLROutputS2xD(149)(0);
  CNStageIntLLRInputS3xD(60)(2) <= VNStageIntLLROutputS2xD(149)(1);
  CNStageIntLLRInputS3xD(146)(2) <= VNStageIntLLROutputS2xD(149)(2);
  CNStageIntLLRInputS3xD(221)(2) <= VNStageIntLLROutputS2xD(149)(3);
  CNStageIntLLRInputS3xD(241)(2) <= VNStageIntLLROutputS2xD(149)(4);
  CNStageIntLLRInputS3xD(309)(2) <= VNStageIntLLROutputS2xD(149)(5);
  CNStageIntLLRInputS3xD(370)(2) <= VNStageIntLLROutputS2xD(149)(6);
  CNStageIntLLRInputS3xD(32)(2) <= VNStageIntLLROutputS2xD(150)(0);
  CNStageIntLLRInputS3xD(86)(2) <= VNStageIntLLROutputS2xD(150)(1);
  CNStageIntLLRInputS3xD(131)(2) <= VNStageIntLLROutputS2xD(150)(2);
  CNStageIntLLRInputS3xD(217)(2) <= VNStageIntLLROutputS2xD(150)(3);
  CNStageIntLLRInputS3xD(312)(2) <= VNStageIntLLROutputS2xD(150)(4);
  CNStageIntLLRInputS3xD(378)(2) <= VNStageIntLLROutputS2xD(150)(5);
  CNStageIntLLRInputS3xD(31)(2) <= VNStageIntLLROutputS2xD(151)(0);
  CNStageIntLLRInputS3xD(92)(2) <= VNStageIntLLROutputS2xD(151)(1);
  CNStageIntLLRInputS3xD(165)(2) <= VNStageIntLLROutputS2xD(151)(2);
  CNStageIntLLRInputS3xD(184)(2) <= VNStageIntLLROutputS2xD(151)(3);
  CNStageIntLLRInputS3xD(238)(2) <= VNStageIntLLROutputS2xD(151)(4);
  CNStageIntLLRInputS3xD(342)(2) <= VNStageIntLLROutputS2xD(151)(5);
  CNStageIntLLRInputS3xD(30)(2) <= VNStageIntLLROutputS2xD(152)(0);
  CNStageIntLLRInputS3xD(76)(2) <= VNStageIntLLROutputS2xD(152)(1);
  CNStageIntLLRInputS3xD(127)(2) <= VNStageIntLLROutputS2xD(152)(2);
  CNStageIntLLRInputS3xD(202)(2) <= VNStageIntLLROutputS2xD(152)(3);
  CNStageIntLLRInputS3xD(228)(2) <= VNStageIntLLROutputS2xD(152)(4);
  CNStageIntLLRInputS3xD(330)(2) <= VNStageIntLLROutputS2xD(152)(5);
  CNStageIntLLRInputS3xD(340)(2) <= VNStageIntLLROutputS2xD(152)(6);
  CNStageIntLLRInputS3xD(29)(2) <= VNStageIntLLROutputS2xD(153)(0);
  CNStageIntLLRInputS3xD(78)(2) <= VNStageIntLLROutputS2xD(153)(1);
  CNStageIntLLRInputS3xD(155)(2) <= VNStageIntLLROutputS2xD(153)(2);
  CNStageIntLLRInputS3xD(203)(2) <= VNStageIntLLROutputS2xD(153)(3);
  CNStageIntLLRInputS3xD(262)(2) <= VNStageIntLLROutputS2xD(153)(4);
  CNStageIntLLRInputS3xD(296)(2) <= VNStageIntLLROutputS2xD(153)(5);
  CNStageIntLLRInputS3xD(376)(2) <= VNStageIntLLROutputS2xD(153)(6);
  CNStageIntLLRInputS3xD(28)(2) <= VNStageIntLLROutputS2xD(154)(0);
  CNStageIntLLRInputS3xD(139)(2) <= VNStageIntLLROutputS2xD(154)(1);
  CNStageIntLLRInputS3xD(183)(2) <= VNStageIntLLROutputS2xD(154)(2);
  CNStageIntLLRInputS3xD(246)(2) <= VNStageIntLLROutputS2xD(154)(3);
  CNStageIntLLRInputS3xD(322)(2) <= VNStageIntLLROutputS2xD(154)(4);
  CNStageIntLLRInputS3xD(27)(2) <= VNStageIntLLROutputS2xD(155)(0);
  CNStageIntLLRInputS3xD(84)(2) <= VNStageIntLLROutputS2xD(155)(1);
  CNStageIntLLRInputS3xD(167)(2) <= VNStageIntLLROutputS2xD(155)(2);
  CNStageIntLLRInputS3xD(174)(2) <= VNStageIntLLROutputS2xD(155)(3);
  CNStageIntLLRInputS3xD(257)(2) <= VNStageIntLLROutputS2xD(155)(4);
  CNStageIntLLRInputS3xD(306)(2) <= VNStageIntLLROutputS2xD(155)(5);
  CNStageIntLLRInputS3xD(357)(2) <= VNStageIntLLROutputS2xD(155)(6);
  CNStageIntLLRInputS3xD(26)(2) <= VNStageIntLLROutputS2xD(156)(0);
  CNStageIntLLRInputS3xD(95)(2) <= VNStageIntLLROutputS2xD(156)(1);
  CNStageIntLLRInputS3xD(157)(2) <= VNStageIntLLROutputS2xD(156)(2);
  CNStageIntLLRInputS3xD(343)(2) <= VNStageIntLLROutputS2xD(156)(3);
  CNStageIntLLRInputS3xD(25)(2) <= VNStageIntLLROutputS2xD(157)(0);
  CNStageIntLLRInputS3xD(102)(2) <= VNStageIntLLROutputS2xD(157)(1);
  CNStageIntLLRInputS3xD(144)(2) <= VNStageIntLLROutputS2xD(157)(2);
  CNStageIntLLRInputS3xD(194)(2) <= VNStageIntLLROutputS2xD(157)(3);
  CNStageIntLLRInputS3xD(323)(2) <= VNStageIntLLROutputS2xD(157)(4);
  CNStageIntLLRInputS3xD(377)(2) <= VNStageIntLLROutputS2xD(157)(5);
  CNStageIntLLRInputS3xD(24)(2) <= VNStageIntLLROutputS2xD(158)(0);
  CNStageIntLLRInputS3xD(77)(2) <= VNStageIntLLROutputS2xD(158)(1);
  CNStageIntLLRInputS3xD(163)(2) <= VNStageIntLLROutputS2xD(158)(2);
  CNStageIntLLRInputS3xD(224)(2) <= VNStageIntLLROutputS2xD(158)(3);
  CNStageIntLLRInputS3xD(230)(2) <= VNStageIntLLROutputS2xD(158)(4);
  CNStageIntLLRInputS3xD(310)(2) <= VNStageIntLLROutputS2xD(158)(5);
  CNStageIntLLRInputS3xD(339)(2) <= VNStageIntLLROutputS2xD(158)(6);
  CNStageIntLLRInputS3xD(23)(2) <= VNStageIntLLROutputS2xD(159)(0);
  CNStageIntLLRInputS3xD(91)(2) <= VNStageIntLLROutputS2xD(159)(1);
  CNStageIntLLRInputS3xD(136)(2) <= VNStageIntLLROutputS2xD(159)(2);
  CNStageIntLLRInputS3xD(271)(2) <= VNStageIntLLROutputS2xD(159)(3);
  CNStageIntLLRInputS3xD(367)(2) <= VNStageIntLLROutputS2xD(159)(4);
  CNStageIntLLRInputS3xD(22)(2) <= VNStageIntLLROutputS2xD(160)(0);
  CNStageIntLLRInputS3xD(62)(2) <= VNStageIntLLROutputS2xD(160)(1);
  CNStageIntLLRInputS3xD(133)(2) <= VNStageIntLLROutputS2xD(160)(2);
  CNStageIntLLRInputS3xD(189)(2) <= VNStageIntLLROutputS2xD(160)(3);
  CNStageIntLLRInputS3xD(233)(2) <= VNStageIntLLROutputS2xD(160)(4);
  CNStageIntLLRInputS3xD(302)(2) <= VNStageIntLLROutputS2xD(160)(5);
  CNStageIntLLRInputS3xD(351)(2) <= VNStageIntLLROutputS2xD(160)(6);
  CNStageIntLLRInputS3xD(21)(2) <= VNStageIntLLROutputS2xD(161)(0);
  CNStageIntLLRInputS3xD(97)(2) <= VNStageIntLLROutputS2xD(161)(1);
  CNStageIntLLRInputS3xD(149)(2) <= VNStageIntLLROutputS2xD(161)(2);
  CNStageIntLLRInputS3xD(171)(2) <= VNStageIntLLROutputS2xD(161)(3);
  CNStageIntLLRInputS3xD(250)(2) <= VNStageIntLLROutputS2xD(161)(4);
  CNStageIntLLRInputS3xD(300)(2) <= VNStageIntLLROutputS2xD(161)(5);
  CNStageIntLLRInputS3xD(379)(2) <= VNStageIntLLROutputS2xD(161)(6);
  CNStageIntLLRInputS3xD(20)(2) <= VNStageIntLLROutputS2xD(162)(0);
  CNStageIntLLRInputS3xD(64)(2) <= VNStageIntLLROutputS2xD(162)(1);
  CNStageIntLLRInputS3xD(141)(2) <= VNStageIntLLROutputS2xD(162)(2);
  CNStageIntLLRInputS3xD(179)(2) <= VNStageIntLLROutputS2xD(162)(3);
  CNStageIntLLRInputS3xD(259)(2) <= VNStageIntLLROutputS2xD(162)(4);
  CNStageIntLLRInputS3xD(315)(2) <= VNStageIntLLROutputS2xD(162)(5);
  CNStageIntLLRInputS3xD(369)(2) <= VNStageIntLLROutputS2xD(162)(6);
  CNStageIntLLRInputS3xD(19)(2) <= VNStageIntLLROutputS2xD(163)(0);
  CNStageIntLLRInputS3xD(79)(2) <= VNStageIntLLROutputS2xD(163)(1);
  CNStageIntLLRInputS3xD(115)(2) <= VNStageIntLLROutputS2xD(163)(2);
  CNStageIntLLRInputS3xD(254)(2) <= VNStageIntLLROutputS2xD(163)(3);
  CNStageIntLLRInputS3xD(355)(2) <= VNStageIntLLROutputS2xD(163)(4);
  CNStageIntLLRInputS3xD(18)(2) <= VNStageIntLLROutputS2xD(164)(0);
  CNStageIntLLRInputS3xD(75)(2) <= VNStageIntLLROutputS2xD(164)(1);
  CNStageIntLLRInputS3xD(125)(2) <= VNStageIntLLROutputS2xD(164)(2);
  CNStageIntLLRInputS3xD(197)(2) <= VNStageIntLLROutputS2xD(164)(3);
  CNStageIntLLRInputS3xD(260)(2) <= VNStageIntLLROutputS2xD(164)(4);
  CNStageIntLLRInputS3xD(375)(2) <= VNStageIntLLROutputS2xD(164)(5);
  CNStageIntLLRInputS3xD(17)(2) <= VNStageIntLLROutputS2xD(165)(0);
  CNStageIntLLRInputS3xD(93)(2) <= VNStageIntLLROutputS2xD(165)(1);
  CNStageIntLLRInputS3xD(119)(2) <= VNStageIntLLROutputS2xD(165)(2);
  CNStageIntLLRInputS3xD(177)(2) <= VNStageIntLLROutputS2xD(165)(3);
  CNStageIntLLRInputS3xD(294)(2) <= VNStageIntLLROutputS2xD(165)(4);
  CNStageIntLLRInputS3xD(348)(2) <= VNStageIntLLROutputS2xD(165)(5);
  CNStageIntLLRInputS3xD(16)(2) <= VNStageIntLLROutputS2xD(166)(0);
  CNStageIntLLRInputS3xD(57)(2) <= VNStageIntLLROutputS2xD(166)(1);
  CNStageIntLLRInputS3xD(122)(2) <= VNStageIntLLROutputS2xD(166)(2);
  CNStageIntLLRInputS3xD(210)(2) <= VNStageIntLLROutputS2xD(166)(3);
  CNStageIntLLRInputS3xD(288)(2) <= VNStageIntLLROutputS2xD(166)(4);
  CNStageIntLLRInputS3xD(345)(2) <= VNStageIntLLROutputS2xD(166)(5);
  CNStageIntLLRInputS3xD(15)(2) <= VNStageIntLLROutputS2xD(167)(0);
  CNStageIntLLRInputS3xD(58)(2) <= VNStageIntLLROutputS2xD(167)(1);
  CNStageIntLLRInputS3xD(112)(2) <= VNStageIntLLROutputS2xD(167)(2);
  CNStageIntLLRInputS3xD(213)(2) <= VNStageIntLLROutputS2xD(167)(3);
  CNStageIntLLRInputS3xD(225)(2) <= VNStageIntLLROutputS2xD(167)(4);
  CNStageIntLLRInputS3xD(292)(2) <= VNStageIntLLROutputS2xD(167)(5);
  CNStageIntLLRInputS3xD(360)(2) <= VNStageIntLLROutputS2xD(167)(6);
  CNStageIntLLRInputS3xD(14)(2) <= VNStageIntLLROutputS2xD(168)(0);
  CNStageIntLLRInputS3xD(150)(2) <= VNStageIntLLROutputS2xD(168)(1);
  CNStageIntLLRInputS3xD(199)(2) <= VNStageIntLLROutputS2xD(168)(2);
  CNStageIntLLRInputS3xD(264)(2) <= VNStageIntLLROutputS2xD(168)(3);
  CNStageIntLLRInputS3xD(283)(2) <= VNStageIntLLROutputS2xD(168)(4);
  CNStageIntLLRInputS3xD(353)(2) <= VNStageIntLLROutputS2xD(168)(5);
  CNStageIntLLRInputS3xD(13)(2) <= VNStageIntLLROutputS2xD(169)(0);
  CNStageIntLLRInputS3xD(85)(2) <= VNStageIntLLROutputS2xD(169)(1);
  CNStageIntLLRInputS3xD(132)(2) <= VNStageIntLLROutputS2xD(169)(2);
  CNStageIntLLRInputS3xD(178)(2) <= VNStageIntLLROutputS2xD(169)(3);
  CNStageIntLLRInputS3xD(266)(2) <= VNStageIntLLROutputS2xD(169)(4);
  CNStageIntLLRInputS3xD(316)(2) <= VNStageIntLLROutputS2xD(169)(5);
  CNStageIntLLRInputS3xD(12)(2) <= VNStageIntLLROutputS2xD(170)(0);
  CNStageIntLLRInputS3xD(101)(2) <= VNStageIntLLROutputS2xD(170)(1);
  CNStageIntLLRInputS3xD(145)(2) <= VNStageIntLLROutputS2xD(170)(2);
  CNStageIntLLRInputS3xD(236)(2) <= VNStageIntLLROutputS2xD(170)(3);
  CNStageIntLLRInputS3xD(337)(2) <= VNStageIntLLROutputS2xD(170)(4);
  CNStageIntLLRInputS3xD(105)(2) <= VNStageIntLLROutputS2xD(171)(0);
  CNStageIntLLRInputS3xD(156)(2) <= VNStageIntLLROutputS2xD(171)(1);
  CNStageIntLLRInputS3xD(222)(2) <= VNStageIntLLROutputS2xD(171)(2);
  CNStageIntLLRInputS3xD(311)(2) <= VNStageIntLLROutputS2xD(171)(3);
  CNStageIntLLRInputS3xD(11)(2) <= VNStageIntLLROutputS2xD(172)(0);
  CNStageIntLLRInputS3xD(110)(2) <= VNStageIntLLROutputS2xD(172)(1);
  CNStageIntLLRInputS3xD(126)(2) <= VNStageIntLLROutputS2xD(172)(2);
  CNStageIntLLRInputS3xD(229)(2) <= VNStageIntLLROutputS2xD(172)(3);
  CNStageIntLLRInputS3xD(10)(2) <= VNStageIntLLROutputS2xD(173)(0);
  CNStageIntLLRInputS3xD(104)(2) <= VNStageIntLLROutputS2xD(173)(1);
  CNStageIntLLRInputS3xD(114)(2) <= VNStageIntLLROutputS2xD(173)(2);
  CNStageIntLLRInputS3xD(180)(2) <= VNStageIntLLROutputS2xD(173)(3);
  CNStageIntLLRInputS3xD(237)(2) <= VNStageIntLLROutputS2xD(173)(4);
  CNStageIntLLRInputS3xD(295)(2) <= VNStageIntLLROutputS2xD(173)(5);
  CNStageIntLLRInputS3xD(9)(2) <= VNStageIntLLROutputS2xD(174)(0);
  CNStageIntLLRInputS3xD(99)(2) <= VNStageIntLLROutputS2xD(174)(1);
  CNStageIntLLRInputS3xD(159)(2) <= VNStageIntLLROutputS2xD(174)(2);
  CNStageIntLLRInputS3xD(265)(2) <= VNStageIntLLROutputS2xD(174)(3);
  CNStageIntLLRInputS3xD(361)(2) <= VNStageIntLLROutputS2xD(174)(4);
  CNStageIntLLRInputS3xD(8)(2) <= VNStageIntLLROutputS2xD(175)(0);
  CNStageIntLLRInputS3xD(82)(2) <= VNStageIntLLROutputS2xD(175)(1);
  CNStageIntLLRInputS3xD(117)(2) <= VNStageIntLLROutputS2xD(175)(2);
  CNStageIntLLRInputS3xD(211)(2) <= VNStageIntLLROutputS2xD(175)(3);
  CNStageIntLLRInputS3xD(278)(2) <= VNStageIntLLROutputS2xD(175)(4);
  CNStageIntLLRInputS3xD(325)(2) <= VNStageIntLLROutputS2xD(175)(5);
  CNStageIntLLRInputS3xD(344)(2) <= VNStageIntLLROutputS2xD(175)(6);
  CNStageIntLLRInputS3xD(7)(2) <= VNStageIntLLROutputS2xD(176)(0);
  CNStageIntLLRInputS3xD(89)(2) <= VNStageIntLLROutputS2xD(176)(1);
  CNStageIntLLRInputS3xD(137)(2) <= VNStageIntLLROutputS2xD(176)(2);
  CNStageIntLLRInputS3xD(176)(2) <= VNStageIntLLROutputS2xD(176)(3);
  CNStageIntLLRInputS3xD(251)(2) <= VNStageIntLLROutputS2xD(176)(4);
  CNStageIntLLRInputS3xD(286)(2) <= VNStageIntLLROutputS2xD(176)(5);
  CNStageIntLLRInputS3xD(356)(2) <= VNStageIntLLROutputS2xD(176)(6);
  CNStageIntLLRInputS3xD(6)(2) <= VNStageIntLLROutputS2xD(177)(0);
  CNStageIntLLRInputS3xD(109)(2) <= VNStageIntLLROutputS2xD(177)(1);
  CNStageIntLLRInputS3xD(147)(2) <= VNStageIntLLROutputS2xD(177)(2);
  CNStageIntLLRInputS3xD(204)(2) <= VNStageIntLLROutputS2xD(177)(3);
  CNStageIntLLRInputS3xD(232)(2) <= VNStageIntLLROutputS2xD(177)(4);
  CNStageIntLLRInputS3xD(304)(2) <= VNStageIntLLROutputS2xD(177)(5);
  CNStageIntLLRInputS3xD(368)(2) <= VNStageIntLLROutputS2xD(177)(6);
  CNStageIntLLRInputS3xD(5)(2) <= VNStageIntLLROutputS2xD(178)(0);
  CNStageIntLLRInputS3xD(107)(2) <= VNStageIntLLROutputS2xD(178)(1);
  CNStageIntLLRInputS3xD(142)(2) <= VNStageIntLLROutputS2xD(178)(2);
  CNStageIntLLRInputS3xD(201)(2) <= VNStageIntLLROutputS2xD(178)(3);
  CNStageIntLLRInputS3xD(313)(2) <= VNStageIntLLROutputS2xD(178)(4);
  CNStageIntLLRInputS3xD(338)(2) <= VNStageIntLLROutputS2xD(178)(5);
  CNStageIntLLRInputS3xD(4)(2) <= VNStageIntLLROutputS2xD(179)(0);
  CNStageIntLLRInputS3xD(87)(2) <= VNStageIntLLROutputS2xD(179)(1);
  CNStageIntLLRInputS3xD(148)(2) <= VNStageIntLLROutputS2xD(179)(2);
  CNStageIntLLRInputS3xD(215)(2) <= VNStageIntLLROutputS2xD(179)(3);
  CNStageIntLLRInputS3xD(267)(2) <= VNStageIntLLROutputS2xD(179)(4);
  CNStageIntLLRInputS3xD(308)(2) <= VNStageIntLLROutputS2xD(179)(5);
  CNStageIntLLRInputS3xD(67)(2) <= VNStageIntLLROutputS2xD(180)(0);
  CNStageIntLLRInputS3xD(208)(2) <= VNStageIntLLROutputS2xD(180)(1);
  CNStageIntLLRInputS3xD(263)(2) <= VNStageIntLLROutputS2xD(180)(2);
  CNStageIntLLRInputS3xD(314)(2) <= VNStageIntLLROutputS2xD(180)(3);
  CNStageIntLLRInputS3xD(371)(2) <= VNStageIntLLROutputS2xD(180)(4);
  CNStageIntLLRInputS3xD(3)(2) <= VNStageIntLLROutputS2xD(181)(0);
  CNStageIntLLRInputS3xD(70)(2) <= VNStageIntLLROutputS2xD(181)(1);
  CNStageIntLLRInputS3xD(162)(2) <= VNStageIntLLROutputS2xD(181)(2);
  CNStageIntLLRInputS3xD(186)(2) <= VNStageIntLLROutputS2xD(181)(3);
  CNStageIntLLRInputS3xD(227)(2) <= VNStageIntLLROutputS2xD(181)(4);
  CNStageIntLLRInputS3xD(303)(2) <= VNStageIntLLROutputS2xD(181)(5);
  CNStageIntLLRInputS3xD(2)(2) <= VNStageIntLLROutputS2xD(182)(0);
  CNStageIntLLRInputS3xD(54)(2) <= VNStageIntLLROutputS2xD(182)(1);
  CNStageIntLLRInputS3xD(169)(2) <= VNStageIntLLROutputS2xD(182)(2);
  CNStageIntLLRInputS3xD(195)(2) <= VNStageIntLLROutputS2xD(182)(3);
  CNStageIntLLRInputS3xD(248)(2) <= VNStageIntLLROutputS2xD(182)(4);
  CNStageIntLLRInputS3xD(328)(2) <= VNStageIntLLROutputS2xD(182)(5);
  CNStageIntLLRInputS3xD(350)(2) <= VNStageIntLLROutputS2xD(182)(6);
  CNStageIntLLRInputS3xD(1)(2) <= VNStageIntLLROutputS2xD(183)(0);
  CNStageIntLLRInputS3xD(88)(2) <= VNStageIntLLROutputS2xD(183)(1);
  CNStageIntLLRInputS3xD(190)(2) <= VNStageIntLLROutputS2xD(183)(2);
  CNStageIntLLRInputS3xD(281)(2) <= VNStageIntLLROutputS2xD(183)(3);
  CNStageIntLLRInputS3xD(358)(2) <= VNStageIntLLROutputS2xD(183)(4);
  CNStageIntLLRInputS3xD(0)(2) <= VNStageIntLLROutputS2xD(184)(0);
  CNStageIntLLRInputS3xD(106)(2) <= VNStageIntLLROutputS2xD(184)(1);
  CNStageIntLLRInputS3xD(153)(2) <= VNStageIntLLROutputS2xD(184)(2);
  CNStageIntLLRInputS3xD(193)(2) <= VNStageIntLLROutputS2xD(184)(3);
  CNStageIntLLRInputS3xD(226)(2) <= VNStageIntLLROutputS2xD(184)(4);
  CNStageIntLLRInputS3xD(318)(2) <= VNStageIntLLROutputS2xD(184)(5);
  CNStageIntLLRInputS3xD(354)(2) <= VNStageIntLLROutputS2xD(184)(6);
  CNStageIntLLRInputS3xD(121)(2) <= VNStageIntLLROutputS2xD(185)(0);
  CNStageIntLLRInputS3xD(272)(2) <= VNStageIntLLROutputS2xD(185)(1);
  CNStageIntLLRInputS3xD(320)(2) <= VNStageIntLLROutputS2xD(185)(2);
  CNStageIntLLRInputS3xD(359)(2) <= VNStageIntLLROutputS2xD(185)(3);
  CNStageIntLLRInputS3xD(63)(2) <= VNStageIntLLROutputS2xD(186)(0);
  CNStageIntLLRInputS3xD(160)(2) <= VNStageIntLLROutputS2xD(186)(1);
  CNStageIntLLRInputS3xD(216)(2) <= VNStageIntLLROutputS2xD(186)(2);
  CNStageIntLLRInputS3xD(235)(2) <= VNStageIntLLROutputS2xD(186)(3);
  CNStageIntLLRInputS3xD(290)(2) <= VNStageIntLLROutputS2xD(186)(4);
  CNStageIntLLRInputS3xD(349)(2) <= VNStageIntLLROutputS2xD(186)(5);
  CNStageIntLLRInputS3xD(90)(2) <= VNStageIntLLROutputS2xD(187)(0);
  CNStageIntLLRInputS3xD(113)(2) <= VNStageIntLLROutputS2xD(187)(1);
  CNStageIntLLRInputS3xD(200)(2) <= VNStageIntLLROutputS2xD(187)(2);
  CNStageIntLLRInputS3xD(240)(2) <= VNStageIntLLROutputS2xD(187)(3);
  CNStageIntLLRInputS3xD(326)(2) <= VNStageIntLLROutputS2xD(187)(4);
  CNStageIntLLRInputS3xD(374)(2) <= VNStageIntLLROutputS2xD(187)(5);
  CNStageIntLLRInputS3xD(81)(2) <= VNStageIntLLROutputS2xD(188)(0);
  CNStageIntLLRInputS3xD(212)(2) <= VNStageIntLLROutputS2xD(188)(1);
  CNStageIntLLRInputS3xD(279)(2) <= VNStageIntLLROutputS2xD(188)(2);
  CNStageIntLLRInputS3xD(284)(2) <= VNStageIntLLROutputS2xD(188)(3);
  CNStageIntLLRInputS3xD(381)(2) <= VNStageIntLLROutputS2xD(188)(4);
  CNStageIntLLRInputS3xD(68)(2) <= VNStageIntLLROutputS2xD(189)(0);
  CNStageIntLLRInputS3xD(152)(2) <= VNStageIntLLROutputS2xD(189)(1);
  CNStageIntLLRInputS3xD(223)(2) <= VNStageIntLLROutputS2xD(189)(2);
  CNStageIntLLRInputS3xD(239)(2) <= VNStageIntLLROutputS2xD(189)(3);
  CNStageIntLLRInputS3xD(291)(2) <= VNStageIntLLROutputS2xD(189)(4);
  CNStageIntLLRInputS3xD(363)(2) <= VNStageIntLLROutputS2xD(189)(5);
  CNStageIntLLRInputS3xD(168)(2) <= VNStageIntLLROutputS2xD(190)(0);
  CNStageIntLLRInputS3xD(196)(2) <= VNStageIntLLROutputS2xD(190)(1);
  CNStageIntLLRInputS3xD(234)(2) <= VNStageIntLLROutputS2xD(190)(2);
  CNStageIntLLRInputS3xD(319)(2) <= VNStageIntLLROutputS2xD(190)(3);
  CNStageIntLLRInputS3xD(365)(2) <= VNStageIntLLROutputS2xD(190)(4);
  CNStageIntLLRInputS3xD(52)(2) <= VNStageIntLLROutputS2xD(191)(0);
  CNStageIntLLRInputS3xD(59)(2) <= VNStageIntLLROutputS2xD(191)(1);
  CNStageIntLLRInputS3xD(138)(2) <= VNStageIntLLROutputS2xD(191)(2);
  CNStageIntLLRInputS3xD(185)(2) <= VNStageIntLLROutputS2xD(191)(3);
  CNStageIntLLRInputS3xD(270)(2) <= VNStageIntLLROutputS2xD(191)(4);
  CNStageIntLLRInputS3xD(280)(2) <= VNStageIntLLROutputS2xD(191)(5);
  CNStageIntLLRInputS3xD(53)(3) <= VNStageIntLLROutputS2xD(192)(0);
  CNStageIntLLRInputS3xD(107)(3) <= VNStageIntLLROutputS2xD(192)(1);
  CNStageIntLLRInputS3xD(128)(3) <= VNStageIntLLROutputS2xD(192)(2);
  CNStageIntLLRInputS3xD(197)(3) <= VNStageIntLLROutputS2xD(192)(3);
  CNStageIntLLRInputS3xD(243)(3) <= VNStageIntLLROutputS2xD(192)(4);
  CNStageIntLLRInputS3xD(297)(3) <= VNStageIntLLROutputS2xD(192)(5);
  CNStageIntLLRInputS3xD(340)(3) <= VNStageIntLLROutputS2xD(192)(6);
  CNStageIntLLRInputS3xD(51)(3) <= VNStageIntLLROutputS2xD(193)(0);
  CNStageIntLLRInputS3xD(58)(3) <= VNStageIntLLROutputS2xD(193)(1);
  CNStageIntLLRInputS3xD(137)(3) <= VNStageIntLLROutputS2xD(193)(2);
  CNStageIntLLRInputS3xD(269)(3) <= VNStageIntLLROutputS2xD(193)(3);
  CNStageIntLLRInputS3xD(333)(3) <= VNStageIntLLROutputS2xD(193)(4);
  CNStageIntLLRInputS3xD(50)(3) <= VNStageIntLLROutputS2xD(194)(0);
  CNStageIntLLRInputS3xD(55)(3) <= VNStageIntLLROutputS2xD(194)(1);
  CNStageIntLLRInputS3xD(115)(3) <= VNStageIntLLROutputS2xD(194)(2);
  CNStageIntLLRInputS3xD(171)(3) <= VNStageIntLLROutputS2xD(194)(3);
  CNStageIntLLRInputS3xD(275)(3) <= VNStageIntLLROutputS2xD(194)(4);
  CNStageIntLLRInputS3xD(304)(3) <= VNStageIntLLROutputS2xD(194)(5);
  CNStageIntLLRInputS3xD(371)(3) <= VNStageIntLLROutputS2xD(194)(6);
  CNStageIntLLRInputS3xD(72)(3) <= VNStageIntLLROutputS2xD(195)(0);
  CNStageIntLLRInputS3xD(139)(3) <= VNStageIntLLROutputS2xD(195)(1);
  CNStageIntLLRInputS3xD(187)(3) <= VNStageIntLLROutputS2xD(195)(2);
  CNStageIntLLRInputS3xD(244)(3) <= VNStageIntLLROutputS2xD(195)(3);
  CNStageIntLLRInputS3xD(49)(3) <= VNStageIntLLROutputS2xD(196)(0);
  CNStageIntLLRInputS3xD(64)(3) <= VNStageIntLLROutputS2xD(196)(1);
  CNStageIntLLRInputS3xD(153)(3) <= VNStageIntLLROutputS2xD(196)(2);
  CNStageIntLLRInputS3xD(205)(3) <= VNStageIntLLROutputS2xD(196)(3);
  CNStageIntLLRInputS3xD(242)(3) <= VNStageIntLLROutputS2xD(196)(4);
  CNStageIntLLRInputS3xD(306)(3) <= VNStageIntLLROutputS2xD(196)(5);
  CNStageIntLLRInputS3xD(48)(3) <= VNStageIntLLROutputS2xD(197)(0);
  CNStageIntLLRInputS3xD(96)(3) <= VNStageIntLLROutputS2xD(197)(1);
  CNStageIntLLRInputS3xD(150)(3) <= VNStageIntLLROutputS2xD(197)(2);
  CNStageIntLLRInputS3xD(213)(3) <= VNStageIntLLROutputS2xD(197)(3);
  CNStageIntLLRInputS3xD(273)(3) <= VNStageIntLLROutputS2xD(197)(4);
  CNStageIntLLRInputS3xD(320)(3) <= VNStageIntLLROutputS2xD(197)(5);
  CNStageIntLLRInputS3xD(363)(3) <= VNStageIntLLROutputS2xD(197)(6);
  CNStageIntLLRInputS3xD(47)(3) <= VNStageIntLLROutputS2xD(198)(0);
  CNStageIntLLRInputS3xD(105)(3) <= VNStageIntLLROutputS2xD(198)(1);
  CNStageIntLLRInputS3xD(111)(3) <= VNStageIntLLROutputS2xD(198)(2);
  CNStageIntLLRInputS3xD(208)(3) <= VNStageIntLLROutputS2xD(198)(3);
  CNStageIntLLRInputS3xD(254)(3) <= VNStageIntLLROutputS2xD(198)(4);
  CNStageIntLLRInputS3xD(316)(3) <= VNStageIntLLROutputS2xD(198)(5);
  CNStageIntLLRInputS3xD(379)(3) <= VNStageIntLLROutputS2xD(198)(6);
  CNStageIntLLRInputS3xD(46)(3) <= VNStageIntLLROutputS2xD(199)(0);
  CNStageIntLLRInputS3xD(99)(3) <= VNStageIntLLROutputS2xD(199)(1);
  CNStageIntLLRInputS3xD(133)(3) <= VNStageIntLLROutputS2xD(199)(2);
  CNStageIntLLRInputS3xD(214)(3) <= VNStageIntLLROutputS2xD(199)(3);
  CNStageIntLLRInputS3xD(257)(3) <= VNStageIntLLROutputS2xD(199)(4);
  CNStageIntLLRInputS3xD(282)(3) <= VNStageIntLLROutputS2xD(199)(5);
  CNStageIntLLRInputS3xD(350)(3) <= VNStageIntLLROutputS2xD(199)(6);
  CNStageIntLLRInputS3xD(45)(3) <= VNStageIntLLROutputS2xD(200)(0);
  CNStageIntLLRInputS3xD(102)(3) <= VNStageIntLLROutputS2xD(200)(1);
  CNStageIntLLRInputS3xD(134)(3) <= VNStageIntLLROutputS2xD(200)(2);
  CNStageIntLLRInputS3xD(204)(3) <= VNStageIntLLROutputS2xD(200)(3);
  CNStageIntLLRInputS3xD(245)(3) <= VNStageIntLLROutputS2xD(200)(4);
  CNStageIntLLRInputS3xD(300)(3) <= VNStageIntLLROutputS2xD(200)(5);
  CNStageIntLLRInputS3xD(44)(3) <= VNStageIntLLROutputS2xD(201)(0);
  CNStageIntLLRInputS3xD(93)(3) <= VNStageIntLLROutputS2xD(201)(1);
  CNStageIntLLRInputS3xD(169)(3) <= VNStageIntLLROutputS2xD(201)(2);
  CNStageIntLLRInputS3xD(174)(3) <= VNStageIntLLROutputS2xD(201)(3);
  CNStageIntLLRInputS3xD(274)(3) <= VNStageIntLLROutputS2xD(201)(4);
  CNStageIntLLRInputS3xD(351)(3) <= VNStageIntLLROutputS2xD(201)(5);
  CNStageIntLLRInputS3xD(43)(3) <= VNStageIntLLROutputS2xD(202)(0);
  CNStageIntLLRInputS3xD(73)(3) <= VNStageIntLLROutputS2xD(202)(1);
  CNStageIntLLRInputS3xD(160)(3) <= VNStageIntLLROutputS2xD(202)(2);
  CNStageIntLLRInputS3xD(181)(3) <= VNStageIntLLROutputS2xD(202)(3);
  CNStageIntLLRInputS3xD(281)(3) <= VNStageIntLLROutputS2xD(202)(4);
  CNStageIntLLRInputS3xD(365)(3) <= VNStageIntLLROutputS2xD(202)(5);
  CNStageIntLLRInputS3xD(42)(3) <= VNStageIntLLROutputS2xD(203)(0);
  CNStageIntLLRInputS3xD(54)(3) <= VNStageIntLLROutputS2xD(203)(1);
  CNStageIntLLRInputS3xD(119)(3) <= VNStageIntLLROutputS2xD(203)(2);
  CNStageIntLLRInputS3xD(217)(3) <= VNStageIntLLROutputS2xD(203)(3);
  CNStageIntLLRInputS3xD(267)(3) <= VNStageIntLLROutputS2xD(203)(4);
  CNStageIntLLRInputS3xD(326)(3) <= VNStageIntLLROutputS2xD(203)(5);
  CNStageIntLLRInputS3xD(361)(3) <= VNStageIntLLROutputS2xD(203)(6);
  CNStageIntLLRInputS3xD(41)(3) <= VNStageIntLLROutputS2xD(204)(0);
  CNStageIntLLRInputS3xD(68)(3) <= VNStageIntLLROutputS2xD(204)(1);
  CNStageIntLLRInputS3xD(123)(3) <= VNStageIntLLROutputS2xD(204)(2);
  CNStageIntLLRInputS3xD(219)(3) <= VNStageIntLLROutputS2xD(204)(3);
  CNStageIntLLRInputS3xD(251)(3) <= VNStageIntLLROutputS2xD(204)(4);
  CNStageIntLLRInputS3xD(288)(3) <= VNStageIntLLROutputS2xD(204)(5);
  CNStageIntLLRInputS3xD(382)(3) <= VNStageIntLLROutputS2xD(204)(6);
  CNStageIntLLRInputS3xD(170)(3) <= VNStageIntLLROutputS2xD(205)(0);
  CNStageIntLLRInputS3xD(276)(3) <= VNStageIntLLROutputS2xD(205)(1);
  CNStageIntLLRInputS3xD(345)(3) <= VNStageIntLLROutputS2xD(205)(2);
  CNStageIntLLRInputS3xD(40)(3) <= VNStageIntLLROutputS2xD(206)(0);
  CNStageIntLLRInputS3xD(122)(3) <= VNStageIntLLROutputS2xD(206)(1);
  CNStageIntLLRInputS3xD(172)(3) <= VNStageIntLLROutputS2xD(206)(2);
  CNStageIntLLRInputS3xD(332)(3) <= VNStageIntLLROutputS2xD(206)(3);
  CNStageIntLLRInputS3xD(346)(3) <= VNStageIntLLROutputS2xD(206)(4);
  CNStageIntLLRInputS3xD(39)(3) <= VNStageIntLLROutputS2xD(207)(0);
  CNStageIntLLRInputS3xD(95)(3) <= VNStageIntLLROutputS2xD(207)(1);
  CNStageIntLLRInputS3xD(117)(3) <= VNStageIntLLROutputS2xD(207)(2);
  CNStageIntLLRInputS3xD(255)(3) <= VNStageIntLLROutputS2xD(207)(3);
  CNStageIntLLRInputS3xD(292)(3) <= VNStageIntLLROutputS2xD(207)(4);
  CNStageIntLLRInputS3xD(381)(3) <= VNStageIntLLROutputS2xD(207)(5);
  CNStageIntLLRInputS3xD(38)(3) <= VNStageIntLLROutputS2xD(208)(0);
  CNStageIntLLRInputS3xD(82)(3) <= VNStageIntLLROutputS2xD(208)(1);
  CNStageIntLLRInputS3xD(157)(3) <= VNStageIntLLROutputS2xD(208)(2);
  CNStageIntLLRInputS3xD(191)(3) <= VNStageIntLLROutputS2xD(208)(3);
  CNStageIntLLRInputS3xD(286)(3) <= VNStageIntLLROutputS2xD(208)(4);
  CNStageIntLLRInputS3xD(372)(3) <= VNStageIntLLROutputS2xD(208)(5);
  CNStageIntLLRInputS3xD(37)(3) <= VNStageIntLLROutputS2xD(209)(0);
  CNStageIntLLRInputS3xD(97)(3) <= VNStageIntLLROutputS2xD(209)(1);
  CNStageIntLLRInputS3xD(165)(3) <= VNStageIntLLROutputS2xD(209)(2);
  CNStageIntLLRInputS3xD(218)(3) <= VNStageIntLLROutputS2xD(209)(3);
  CNStageIntLLRInputS3xD(323)(3) <= VNStageIntLLROutputS2xD(209)(4);
  CNStageIntLLRInputS3xD(36)(3) <= VNStageIntLLROutputS2xD(210)(0);
  CNStageIntLLRInputS3xD(60)(3) <= VNStageIntLLROutputS2xD(210)(1);
  CNStageIntLLRInputS3xD(129)(3) <= VNStageIntLLROutputS2xD(210)(2);
  CNStageIntLLRInputS3xD(180)(3) <= VNStageIntLLROutputS2xD(210)(3);
  CNStageIntLLRInputS3xD(246)(3) <= VNStageIntLLROutputS2xD(210)(4);
  CNStageIntLLRInputS3xD(330)(3) <= VNStageIntLLROutputS2xD(210)(5);
  CNStageIntLLRInputS3xD(335)(3) <= VNStageIntLLROutputS2xD(210)(6);
  CNStageIntLLRInputS3xD(35)(3) <= VNStageIntLLROutputS2xD(211)(0);
  CNStageIntLLRInputS3xD(70)(3) <= VNStageIntLLROutputS2xD(211)(1);
  CNStageIntLLRInputS3xD(127)(3) <= VNStageIntLLROutputS2xD(211)(2);
  CNStageIntLLRInputS3xD(206)(3) <= VNStageIntLLROutputS2xD(211)(3);
  CNStageIntLLRInputS3xD(260)(3) <= VNStageIntLLROutputS2xD(211)(4);
  CNStageIntLLRInputS3xD(298)(3) <= VNStageIntLLROutputS2xD(211)(5);
  CNStageIntLLRInputS3xD(34)(3) <= VNStageIntLLROutputS2xD(212)(0);
  CNStageIntLLRInputS3xD(65)(3) <= VNStageIntLLROutputS2xD(212)(1);
  CNStageIntLLRInputS3xD(163)(3) <= VNStageIntLLROutputS2xD(212)(2);
  CNStageIntLLRInputS3xD(186)(3) <= VNStageIntLLROutputS2xD(212)(3);
  CNStageIntLLRInputS3xD(296)(3) <= VNStageIntLLROutputS2xD(212)(4);
  CNStageIntLLRInputS3xD(33)(3) <= VNStageIntLLROutputS2xD(213)(0);
  CNStageIntLLRInputS3xD(71)(3) <= VNStageIntLLROutputS2xD(213)(1);
  CNStageIntLLRInputS3xD(142)(3) <= VNStageIntLLROutputS2xD(213)(2);
  CNStageIntLLRInputS3xD(230)(3) <= VNStageIntLLROutputS2xD(213)(3);
  CNStageIntLLRInputS3xD(32)(3) <= VNStageIntLLROutputS2xD(214)(0);
  CNStageIntLLRInputS3xD(59)(3) <= VNStageIntLLROutputS2xD(214)(1);
  CNStageIntLLRInputS3xD(145)(3) <= VNStageIntLLROutputS2xD(214)(2);
  CNStageIntLLRInputS3xD(220)(3) <= VNStageIntLLROutputS2xD(214)(3);
  CNStageIntLLRInputS3xD(240)(3) <= VNStageIntLLROutputS2xD(214)(4);
  CNStageIntLLRInputS3xD(308)(3) <= VNStageIntLLROutputS2xD(214)(5);
  CNStageIntLLRInputS3xD(369)(3) <= VNStageIntLLROutputS2xD(214)(6);
  CNStageIntLLRInputS3xD(31)(3) <= VNStageIntLLROutputS2xD(215)(0);
  CNStageIntLLRInputS3xD(85)(3) <= VNStageIntLLROutputS2xD(215)(1);
  CNStageIntLLRInputS3xD(130)(3) <= VNStageIntLLROutputS2xD(215)(2);
  CNStageIntLLRInputS3xD(216)(3) <= VNStageIntLLROutputS2xD(215)(3);
  CNStageIntLLRInputS3xD(234)(3) <= VNStageIntLLROutputS2xD(215)(4);
  CNStageIntLLRInputS3xD(311)(3) <= VNStageIntLLROutputS2xD(215)(5);
  CNStageIntLLRInputS3xD(377)(3) <= VNStageIntLLROutputS2xD(215)(6);
  CNStageIntLLRInputS3xD(30)(3) <= VNStageIntLLROutputS2xD(216)(0);
  CNStageIntLLRInputS3xD(91)(3) <= VNStageIntLLROutputS2xD(216)(1);
  CNStageIntLLRInputS3xD(164)(3) <= VNStageIntLLROutputS2xD(216)(2);
  CNStageIntLLRInputS3xD(183)(3) <= VNStageIntLLROutputS2xD(216)(3);
  CNStageIntLLRInputS3xD(237)(3) <= VNStageIntLLROutputS2xD(216)(4);
  CNStageIntLLRInputS3xD(299)(3) <= VNStageIntLLROutputS2xD(216)(5);
  CNStageIntLLRInputS3xD(341)(3) <= VNStageIntLLROutputS2xD(216)(6);
  CNStageIntLLRInputS3xD(29)(3) <= VNStageIntLLROutputS2xD(217)(0);
  CNStageIntLLRInputS3xD(75)(3) <= VNStageIntLLROutputS2xD(217)(1);
  CNStageIntLLRInputS3xD(126)(3) <= VNStageIntLLROutputS2xD(217)(2);
  CNStageIntLLRInputS3xD(201)(3) <= VNStageIntLLROutputS2xD(217)(3);
  CNStageIntLLRInputS3xD(227)(3) <= VNStageIntLLROutputS2xD(217)(4);
  CNStageIntLLRInputS3xD(329)(3) <= VNStageIntLLROutputS2xD(217)(5);
  CNStageIntLLRInputS3xD(339)(3) <= VNStageIntLLROutputS2xD(217)(6);
  CNStageIntLLRInputS3xD(28)(3) <= VNStageIntLLROutputS2xD(218)(0);
  CNStageIntLLRInputS3xD(77)(3) <= VNStageIntLLROutputS2xD(218)(1);
  CNStageIntLLRInputS3xD(154)(3) <= VNStageIntLLROutputS2xD(218)(2);
  CNStageIntLLRInputS3xD(202)(3) <= VNStageIntLLROutputS2xD(218)(3);
  CNStageIntLLRInputS3xD(261)(3) <= VNStageIntLLROutputS2xD(218)(4);
  CNStageIntLLRInputS3xD(295)(3) <= VNStageIntLLROutputS2xD(218)(5);
  CNStageIntLLRInputS3xD(375)(3) <= VNStageIntLLROutputS2xD(218)(6);
  CNStageIntLLRInputS3xD(27)(3) <= VNStageIntLLROutputS2xD(219)(0);
  CNStageIntLLRInputS3xD(101)(3) <= VNStageIntLLROutputS2xD(219)(1);
  CNStageIntLLRInputS3xD(138)(3) <= VNStageIntLLROutputS2xD(219)(2);
  CNStageIntLLRInputS3xD(182)(3) <= VNStageIntLLROutputS2xD(219)(3);
  CNStageIntLLRInputS3xD(321)(3) <= VNStageIntLLROutputS2xD(219)(4);
  CNStageIntLLRInputS3xD(354)(3) <= VNStageIntLLROutputS2xD(219)(5);
  CNStageIntLLRInputS3xD(26)(3) <= VNStageIntLLROutputS2xD(220)(0);
  CNStageIntLLRInputS3xD(83)(3) <= VNStageIntLLROutputS2xD(220)(1);
  CNStageIntLLRInputS3xD(166)(3) <= VNStageIntLLROutputS2xD(220)(2);
  CNStageIntLLRInputS3xD(173)(3) <= VNStageIntLLROutputS2xD(220)(3);
  CNStageIntLLRInputS3xD(256)(3) <= VNStageIntLLROutputS2xD(220)(4);
  CNStageIntLLRInputS3xD(305)(3) <= VNStageIntLLROutputS2xD(220)(5);
  CNStageIntLLRInputS3xD(356)(3) <= VNStageIntLLROutputS2xD(220)(6);
  CNStageIntLLRInputS3xD(25)(3) <= VNStageIntLLROutputS2xD(221)(0);
  CNStageIntLLRInputS3xD(94)(3) <= VNStageIntLLROutputS2xD(221)(1);
  CNStageIntLLRInputS3xD(156)(3) <= VNStageIntLLROutputS2xD(221)(2);
  CNStageIntLLRInputS3xD(190)(3) <= VNStageIntLLROutputS2xD(221)(3);
  CNStageIntLLRInputS3xD(268)(3) <= VNStageIntLLROutputS2xD(221)(4);
  CNStageIntLLRInputS3xD(331)(3) <= VNStageIntLLROutputS2xD(221)(5);
  CNStageIntLLRInputS3xD(342)(3) <= VNStageIntLLROutputS2xD(221)(6);
  CNStageIntLLRInputS3xD(24)(3) <= VNStageIntLLROutputS2xD(222)(0);
  CNStageIntLLRInputS3xD(143)(3) <= VNStageIntLLROutputS2xD(222)(1);
  CNStageIntLLRInputS3xD(241)(3) <= VNStageIntLLROutputS2xD(222)(2);
  CNStageIntLLRInputS3xD(376)(3) <= VNStageIntLLROutputS2xD(222)(3);
  CNStageIntLLRInputS3xD(23)(3) <= VNStageIntLLROutputS2xD(223)(0);
  CNStageIntLLRInputS3xD(76)(3) <= VNStageIntLLROutputS2xD(223)(1);
  CNStageIntLLRInputS3xD(162)(3) <= VNStageIntLLROutputS2xD(223)(2);
  CNStageIntLLRInputS3xD(224)(3) <= VNStageIntLLROutputS2xD(223)(3);
  CNStageIntLLRInputS3xD(229)(3) <= VNStageIntLLROutputS2xD(223)(4);
  CNStageIntLLRInputS3xD(309)(3) <= VNStageIntLLROutputS2xD(223)(5);
  CNStageIntLLRInputS3xD(338)(3) <= VNStageIntLLROutputS2xD(223)(6);
  CNStageIntLLRInputS3xD(22)(3) <= VNStageIntLLROutputS2xD(224)(0);
  CNStageIntLLRInputS3xD(90)(3) <= VNStageIntLLROutputS2xD(224)(1);
  CNStageIntLLRInputS3xD(135)(3) <= VNStageIntLLROutputS2xD(224)(2);
  CNStageIntLLRInputS3xD(193)(3) <= VNStageIntLLROutputS2xD(224)(3);
  CNStageIntLLRInputS3xD(270)(3) <= VNStageIntLLROutputS2xD(224)(4);
  CNStageIntLLRInputS3xD(328)(3) <= VNStageIntLLROutputS2xD(224)(5);
  CNStageIntLLRInputS3xD(366)(3) <= VNStageIntLLROutputS2xD(224)(6);
  CNStageIntLLRInputS3xD(21)(3) <= VNStageIntLLROutputS2xD(225)(0);
  CNStageIntLLRInputS3xD(61)(3) <= VNStageIntLLROutputS2xD(225)(1);
  CNStageIntLLRInputS3xD(132)(3) <= VNStageIntLLROutputS2xD(225)(2);
  CNStageIntLLRInputS3xD(188)(3) <= VNStageIntLLROutputS2xD(225)(3);
  CNStageIntLLRInputS3xD(232)(3) <= VNStageIntLLROutputS2xD(225)(4);
  CNStageIntLLRInputS3xD(301)(3) <= VNStageIntLLROutputS2xD(225)(5);
  CNStageIntLLRInputS3xD(20)(3) <= VNStageIntLLROutputS2xD(226)(0);
  CNStageIntLLRInputS3xD(148)(3) <= VNStageIntLLROutputS2xD(226)(1);
  CNStageIntLLRInputS3xD(378)(3) <= VNStageIntLLROutputS2xD(226)(2);
  CNStageIntLLRInputS3xD(19)(3) <= VNStageIntLLROutputS2xD(227)(0);
  CNStageIntLLRInputS3xD(63)(3) <= VNStageIntLLROutputS2xD(227)(1);
  CNStageIntLLRInputS3xD(140)(3) <= VNStageIntLLROutputS2xD(227)(2);
  CNStageIntLLRInputS3xD(178)(3) <= VNStageIntLLROutputS2xD(227)(3);
  CNStageIntLLRInputS3xD(258)(3) <= VNStageIntLLROutputS2xD(227)(4);
  CNStageIntLLRInputS3xD(314)(3) <= VNStageIntLLROutputS2xD(227)(5);
  CNStageIntLLRInputS3xD(368)(3) <= VNStageIntLLROutputS2xD(227)(6);
  CNStageIntLLRInputS3xD(18)(3) <= VNStageIntLLROutputS2xD(228)(0);
  CNStageIntLLRInputS3xD(78)(3) <= VNStageIntLLROutputS2xD(228)(1);
  CNStageIntLLRInputS3xD(114)(3) <= VNStageIntLLROutputS2xD(228)(2);
  CNStageIntLLRInputS3xD(198)(3) <= VNStageIntLLROutputS2xD(228)(3);
  CNStageIntLLRInputS3xD(253)(3) <= VNStageIntLLROutputS2xD(228)(4);
  CNStageIntLLRInputS3xD(307)(3) <= VNStageIntLLROutputS2xD(228)(5);
  CNStageIntLLRInputS3xD(17)(3) <= VNStageIntLLROutputS2xD(229)(0);
  CNStageIntLLRInputS3xD(74)(3) <= VNStageIntLLROutputS2xD(229)(1);
  CNStageIntLLRInputS3xD(124)(3) <= VNStageIntLLROutputS2xD(229)(2);
  CNStageIntLLRInputS3xD(259)(3) <= VNStageIntLLROutputS2xD(229)(3);
  CNStageIntLLRInputS3xD(374)(3) <= VNStageIntLLROutputS2xD(229)(4);
  CNStageIntLLRInputS3xD(16)(3) <= VNStageIntLLROutputS2xD(230)(0);
  CNStageIntLLRInputS3xD(118)(3) <= VNStageIntLLROutputS2xD(230)(1);
  CNStageIntLLRInputS3xD(176)(3) <= VNStageIntLLROutputS2xD(230)(2);
  CNStageIntLLRInputS3xD(249)(3) <= VNStageIntLLROutputS2xD(230)(3);
  CNStageIntLLRInputS3xD(293)(3) <= VNStageIntLLROutputS2xD(230)(4);
  CNStageIntLLRInputS3xD(347)(3) <= VNStageIntLLROutputS2xD(230)(5);
  CNStageIntLLRInputS3xD(15)(3) <= VNStageIntLLROutputS2xD(231)(0);
  CNStageIntLLRInputS3xD(56)(3) <= VNStageIntLLROutputS2xD(231)(1);
  CNStageIntLLRInputS3xD(209)(3) <= VNStageIntLLROutputS2xD(231)(2);
  CNStageIntLLRInputS3xD(272)(3) <= VNStageIntLLROutputS2xD(231)(3);
  CNStageIntLLRInputS3xD(287)(3) <= VNStageIntLLROutputS2xD(231)(4);
  CNStageIntLLRInputS3xD(344)(3) <= VNStageIntLLROutputS2xD(231)(5);
  CNStageIntLLRInputS3xD(14)(3) <= VNStageIntLLROutputS2xD(232)(0);
  CNStageIntLLRInputS3xD(57)(3) <= VNStageIntLLROutputS2xD(232)(1);
  CNStageIntLLRInputS3xD(212)(3) <= VNStageIntLLROutputS2xD(232)(2);
  CNStageIntLLRInputS3xD(278)(3) <= VNStageIntLLROutputS2xD(232)(3);
  CNStageIntLLRInputS3xD(291)(3) <= VNStageIntLLROutputS2xD(232)(4);
  CNStageIntLLRInputS3xD(359)(3) <= VNStageIntLLROutputS2xD(232)(5);
  CNStageIntLLRInputS3xD(13)(3) <= VNStageIntLLROutputS2xD(233)(0);
  CNStageIntLLRInputS3xD(92)(3) <= VNStageIntLLROutputS2xD(233)(1);
  CNStageIntLLRInputS3xD(149)(3) <= VNStageIntLLROutputS2xD(233)(2);
  CNStageIntLLRInputS3xD(263)(3) <= VNStageIntLLROutputS2xD(233)(3);
  CNStageIntLLRInputS3xD(352)(3) <= VNStageIntLLROutputS2xD(233)(4);
  CNStageIntLLRInputS3xD(12)(3) <= VNStageIntLLROutputS2xD(234)(0);
  CNStageIntLLRInputS3xD(84)(3) <= VNStageIntLLROutputS2xD(234)(1);
  CNStageIntLLRInputS3xD(131)(3) <= VNStageIntLLROutputS2xD(234)(2);
  CNStageIntLLRInputS3xD(177)(3) <= VNStageIntLLROutputS2xD(234)(3);
  CNStageIntLLRInputS3xD(265)(3) <= VNStageIntLLROutputS2xD(234)(4);
  CNStageIntLLRInputS3xD(315)(3) <= VNStageIntLLROutputS2xD(234)(5);
  CNStageIntLLRInputS3xD(100)(3) <= VNStageIntLLROutputS2xD(235)(0);
  CNStageIntLLRInputS3xD(144)(3) <= VNStageIntLLROutputS2xD(235)(1);
  CNStageIntLLRInputS3xD(196)(3) <= VNStageIntLLROutputS2xD(235)(2);
  CNStageIntLLRInputS3xD(235)(3) <= VNStageIntLLROutputS2xD(235)(3);
  CNStageIntLLRInputS3xD(336)(3) <= VNStageIntLLROutputS2xD(235)(4);
  CNStageIntLLRInputS3xD(11)(3) <= VNStageIntLLROutputS2xD(236)(0);
  CNStageIntLLRInputS3xD(104)(3) <= VNStageIntLLROutputS2xD(236)(1);
  CNStageIntLLRInputS3xD(155)(3) <= VNStageIntLLROutputS2xD(236)(2);
  CNStageIntLLRInputS3xD(221)(3) <= VNStageIntLLROutputS2xD(236)(3);
  CNStageIntLLRInputS3xD(271)(3) <= VNStageIntLLROutputS2xD(236)(4);
  CNStageIntLLRInputS3xD(310)(3) <= VNStageIntLLROutputS2xD(236)(5);
  CNStageIntLLRInputS3xD(10)(3) <= VNStageIntLLROutputS2xD(237)(0);
  CNStageIntLLRInputS3xD(110)(3) <= VNStageIntLLROutputS2xD(237)(1);
  CNStageIntLLRInputS3xD(125)(3) <= VNStageIntLLROutputS2xD(237)(2);
  CNStageIntLLRInputS3xD(228)(3) <= VNStageIntLLROutputS2xD(237)(3);
  CNStageIntLLRInputS3xD(322)(3) <= VNStageIntLLROutputS2xD(237)(4);
  CNStageIntLLRInputS3xD(334)(3) <= VNStageIntLLROutputS2xD(237)(5);
  CNStageIntLLRInputS3xD(9)(3) <= VNStageIntLLROutputS2xD(238)(0);
  CNStageIntLLRInputS3xD(103)(3) <= VNStageIntLLROutputS2xD(238)(1);
  CNStageIntLLRInputS3xD(113)(3) <= VNStageIntLLROutputS2xD(238)(2);
  CNStageIntLLRInputS3xD(179)(3) <= VNStageIntLLROutputS2xD(238)(3);
  CNStageIntLLRInputS3xD(236)(3) <= VNStageIntLLROutputS2xD(238)(4);
  CNStageIntLLRInputS3xD(294)(3) <= VNStageIntLLROutputS2xD(238)(5);
  CNStageIntLLRInputS3xD(383)(3) <= VNStageIntLLROutputS2xD(238)(6);
  CNStageIntLLRInputS3xD(8)(3) <= VNStageIntLLROutputS2xD(239)(0);
  CNStageIntLLRInputS3xD(98)(3) <= VNStageIntLLROutputS2xD(239)(1);
  CNStageIntLLRInputS3xD(158)(3) <= VNStageIntLLROutputS2xD(239)(2);
  CNStageIntLLRInputS3xD(223)(3) <= VNStageIntLLROutputS2xD(239)(3);
  CNStageIntLLRInputS3xD(264)(3) <= VNStageIntLLROutputS2xD(239)(4);
  CNStageIntLLRInputS3xD(284)(3) <= VNStageIntLLROutputS2xD(239)(5);
  CNStageIntLLRInputS3xD(360)(3) <= VNStageIntLLROutputS2xD(239)(6);
  CNStageIntLLRInputS3xD(7)(3) <= VNStageIntLLROutputS2xD(240)(0);
  CNStageIntLLRInputS3xD(81)(3) <= VNStageIntLLROutputS2xD(240)(1);
  CNStageIntLLRInputS3xD(116)(3) <= VNStageIntLLROutputS2xD(240)(2);
  CNStageIntLLRInputS3xD(210)(3) <= VNStageIntLLROutputS2xD(240)(3);
  CNStageIntLLRInputS3xD(277)(3) <= VNStageIntLLROutputS2xD(240)(4);
  CNStageIntLLRInputS3xD(324)(3) <= VNStageIntLLROutputS2xD(240)(5);
  CNStageIntLLRInputS3xD(343)(3) <= VNStageIntLLROutputS2xD(240)(6);
  CNStageIntLLRInputS3xD(6)(3) <= VNStageIntLLROutputS2xD(241)(0);
  CNStageIntLLRInputS3xD(88)(3) <= VNStageIntLLROutputS2xD(241)(1);
  CNStageIntLLRInputS3xD(175)(3) <= VNStageIntLLROutputS2xD(241)(2);
  CNStageIntLLRInputS3xD(250)(3) <= VNStageIntLLROutputS2xD(241)(3);
  CNStageIntLLRInputS3xD(285)(3) <= VNStageIntLLROutputS2xD(241)(4);
  CNStageIntLLRInputS3xD(355)(3) <= VNStageIntLLROutputS2xD(241)(5);
  CNStageIntLLRInputS3xD(5)(3) <= VNStageIntLLROutputS2xD(242)(0);
  CNStageIntLLRInputS3xD(108)(3) <= VNStageIntLLROutputS2xD(242)(1);
  CNStageIntLLRInputS3xD(146)(3) <= VNStageIntLLROutputS2xD(242)(2);
  CNStageIntLLRInputS3xD(203)(3) <= VNStageIntLLROutputS2xD(242)(3);
  CNStageIntLLRInputS3xD(231)(3) <= VNStageIntLLROutputS2xD(242)(4);
  CNStageIntLLRInputS3xD(303)(3) <= VNStageIntLLROutputS2xD(242)(5);
  CNStageIntLLRInputS3xD(367)(3) <= VNStageIntLLROutputS2xD(242)(6);
  CNStageIntLLRInputS3xD(4)(3) <= VNStageIntLLROutputS2xD(243)(0);
  CNStageIntLLRInputS3xD(106)(3) <= VNStageIntLLROutputS2xD(243)(1);
  CNStageIntLLRInputS3xD(141)(3) <= VNStageIntLLROutputS2xD(243)(2);
  CNStageIntLLRInputS3xD(200)(3) <= VNStageIntLLROutputS2xD(243)(3);
  CNStageIntLLRInputS3xD(252)(3) <= VNStageIntLLROutputS2xD(243)(4);
  CNStageIntLLRInputS3xD(312)(3) <= VNStageIntLLROutputS2xD(243)(5);
  CNStageIntLLRInputS3xD(337)(3) <= VNStageIntLLROutputS2xD(243)(6);
  CNStageIntLLRInputS3xD(147)(3) <= VNStageIntLLROutputS2xD(244)(0);
  CNStageIntLLRInputS3xD(266)(3) <= VNStageIntLLROutputS2xD(244)(1);
  CNStageIntLLRInputS3xD(3)(3) <= VNStageIntLLROutputS2xD(245)(0);
  CNStageIntLLRInputS3xD(66)(3) <= VNStageIntLLROutputS2xD(245)(1);
  CNStageIntLLRInputS3xD(136)(3) <= VNStageIntLLROutputS2xD(245)(2);
  CNStageIntLLRInputS3xD(207)(3) <= VNStageIntLLROutputS2xD(245)(3);
  CNStageIntLLRInputS3xD(262)(3) <= VNStageIntLLROutputS2xD(245)(4);
  CNStageIntLLRInputS3xD(313)(3) <= VNStageIntLLROutputS2xD(245)(5);
  CNStageIntLLRInputS3xD(370)(3) <= VNStageIntLLROutputS2xD(245)(6);
  CNStageIntLLRInputS3xD(2)(3) <= VNStageIntLLROutputS2xD(246)(0);
  CNStageIntLLRInputS3xD(69)(3) <= VNStageIntLLROutputS2xD(246)(1);
  CNStageIntLLRInputS3xD(161)(3) <= VNStageIntLLROutputS2xD(246)(2);
  CNStageIntLLRInputS3xD(185)(3) <= VNStageIntLLROutputS2xD(246)(3);
  CNStageIntLLRInputS3xD(226)(3) <= VNStageIntLLROutputS2xD(246)(4);
  CNStageIntLLRInputS3xD(302)(3) <= VNStageIntLLROutputS2xD(246)(5);
  CNStageIntLLRInputS3xD(1)(3) <= VNStageIntLLROutputS2xD(247)(0);
  CNStageIntLLRInputS3xD(109)(3) <= VNStageIntLLROutputS2xD(247)(1);
  CNStageIntLLRInputS3xD(168)(3) <= VNStageIntLLROutputS2xD(247)(2);
  CNStageIntLLRInputS3xD(194)(3) <= VNStageIntLLROutputS2xD(247)(3);
  CNStageIntLLRInputS3xD(247)(3) <= VNStageIntLLROutputS2xD(247)(4);
  CNStageIntLLRInputS3xD(327)(3) <= VNStageIntLLROutputS2xD(247)(5);
  CNStageIntLLRInputS3xD(349)(3) <= VNStageIntLLROutputS2xD(247)(6);
  CNStageIntLLRInputS3xD(0)(3) <= VNStageIntLLROutputS2xD(248)(0);
  CNStageIntLLRInputS3xD(87)(3) <= VNStageIntLLROutputS2xD(248)(1);
  CNStageIntLLRInputS3xD(151)(3) <= VNStageIntLLROutputS2xD(248)(2);
  CNStageIntLLRInputS3xD(189)(3) <= VNStageIntLLROutputS2xD(248)(3);
  CNStageIntLLRInputS3xD(248)(3) <= VNStageIntLLROutputS2xD(248)(4);
  CNStageIntLLRInputS3xD(280)(3) <= VNStageIntLLROutputS2xD(248)(5);
  CNStageIntLLRInputS3xD(357)(3) <= VNStageIntLLROutputS2xD(248)(6);
  CNStageIntLLRInputS3xD(152)(3) <= VNStageIntLLROutputS2xD(249)(0);
  CNStageIntLLRInputS3xD(192)(3) <= VNStageIntLLROutputS2xD(249)(1);
  CNStageIntLLRInputS3xD(225)(3) <= VNStageIntLLROutputS2xD(249)(2);
  CNStageIntLLRInputS3xD(317)(3) <= VNStageIntLLROutputS2xD(249)(3);
  CNStageIntLLRInputS3xD(353)(3) <= VNStageIntLLROutputS2xD(249)(4);
  CNStageIntLLRInputS3xD(79)(3) <= VNStageIntLLROutputS2xD(250)(0);
  CNStageIntLLRInputS3xD(120)(3) <= VNStageIntLLROutputS2xD(250)(1);
  CNStageIntLLRInputS3xD(184)(3) <= VNStageIntLLROutputS2xD(250)(2);
  CNStageIntLLRInputS3xD(319)(3) <= VNStageIntLLROutputS2xD(250)(3);
  CNStageIntLLRInputS3xD(358)(3) <= VNStageIntLLROutputS2xD(250)(4);
  CNStageIntLLRInputS3xD(62)(3) <= VNStageIntLLROutputS2xD(251)(0);
  CNStageIntLLRInputS3xD(159)(3) <= VNStageIntLLROutputS2xD(251)(1);
  CNStageIntLLRInputS3xD(215)(3) <= VNStageIntLLROutputS2xD(251)(2);
  CNStageIntLLRInputS3xD(289)(3) <= VNStageIntLLROutputS2xD(251)(3);
  CNStageIntLLRInputS3xD(348)(3) <= VNStageIntLLROutputS2xD(251)(4);
  CNStageIntLLRInputS3xD(89)(3) <= VNStageIntLLROutputS2xD(252)(0);
  CNStageIntLLRInputS3xD(112)(3) <= VNStageIntLLROutputS2xD(252)(1);
  CNStageIntLLRInputS3xD(199)(3) <= VNStageIntLLROutputS2xD(252)(2);
  CNStageIntLLRInputS3xD(239)(3) <= VNStageIntLLROutputS2xD(252)(3);
  CNStageIntLLRInputS3xD(325)(3) <= VNStageIntLLROutputS2xD(252)(4);
  CNStageIntLLRInputS3xD(373)(3) <= VNStageIntLLROutputS2xD(252)(5);
  CNStageIntLLRInputS3xD(80)(3) <= VNStageIntLLROutputS2xD(253)(0);
  CNStageIntLLRInputS3xD(121)(3) <= VNStageIntLLROutputS2xD(253)(1);
  CNStageIntLLRInputS3xD(211)(3) <= VNStageIntLLROutputS2xD(253)(2);
  CNStageIntLLRInputS3xD(279)(3) <= VNStageIntLLROutputS2xD(253)(3);
  CNStageIntLLRInputS3xD(283)(3) <= VNStageIntLLROutputS2xD(253)(4);
  CNStageIntLLRInputS3xD(380)(3) <= VNStageIntLLROutputS2xD(253)(5);
  CNStageIntLLRInputS3xD(67)(3) <= VNStageIntLLROutputS2xD(254)(0);
  CNStageIntLLRInputS3xD(222)(3) <= VNStageIntLLROutputS2xD(254)(1);
  CNStageIntLLRInputS3xD(238)(3) <= VNStageIntLLROutputS2xD(254)(2);
  CNStageIntLLRInputS3xD(290)(3) <= VNStageIntLLROutputS2xD(254)(3);
  CNStageIntLLRInputS3xD(362)(3) <= VNStageIntLLROutputS2xD(254)(4);
  CNStageIntLLRInputS3xD(52)(3) <= VNStageIntLLROutputS2xD(255)(0);
  CNStageIntLLRInputS3xD(86)(3) <= VNStageIntLLROutputS2xD(255)(1);
  CNStageIntLLRInputS3xD(167)(3) <= VNStageIntLLROutputS2xD(255)(2);
  CNStageIntLLRInputS3xD(195)(3) <= VNStageIntLLROutputS2xD(255)(3);
  CNStageIntLLRInputS3xD(233)(3) <= VNStageIntLLROutputS2xD(255)(4);
  CNStageIntLLRInputS3xD(318)(3) <= VNStageIntLLROutputS2xD(255)(5);
  CNStageIntLLRInputS3xD(364)(3) <= VNStageIntLLROutputS2xD(255)(6);
  CNStageIntLLRInputS3xD(53)(4) <= VNStageIntLLROutputS2xD(256)(0);
  CNStageIntLLRInputS3xD(106)(4) <= VNStageIntLLROutputS2xD(256)(1);
  CNStageIntLLRInputS3xD(127)(4) <= VNStageIntLLROutputS2xD(256)(2);
  CNStageIntLLRInputS3xD(242)(4) <= VNStageIntLLROutputS2xD(256)(3);
  CNStageIntLLRInputS3xD(296)(4) <= VNStageIntLLROutputS2xD(256)(4);
  CNStageIntLLRInputS3xD(339)(4) <= VNStageIntLLROutputS2xD(256)(5);
  CNStageIntLLRInputS3xD(51)(4) <= VNStageIntLLROutputS2xD(257)(0);
  CNStageIntLLRInputS3xD(85)(4) <= VNStageIntLLROutputS2xD(257)(1);
  CNStageIntLLRInputS3xD(166)(4) <= VNStageIntLLROutputS2xD(257)(2);
  CNStageIntLLRInputS3xD(194)(4) <= VNStageIntLLROutputS2xD(257)(3);
  CNStageIntLLRInputS3xD(232)(4) <= VNStageIntLLROutputS2xD(257)(4);
  CNStageIntLLRInputS3xD(317)(4) <= VNStageIntLLROutputS2xD(257)(5);
  CNStageIntLLRInputS3xD(363)(4) <= VNStageIntLLROutputS2xD(257)(6);
  CNStageIntLLRInputS3xD(50)(4) <= VNStageIntLLROutputS2xD(258)(0);
  CNStageIntLLRInputS3xD(57)(4) <= VNStageIntLLROutputS2xD(258)(1);
  CNStageIntLLRInputS3xD(331)(4) <= VNStageIntLLROutputS2xD(258)(2);
  CNStageIntLLRInputS3xD(54)(4) <= VNStageIntLLROutputS2xD(259)(0);
  CNStageIntLLRInputS3xD(114)(4) <= VNStageIntLLROutputS2xD(259)(1);
  CNStageIntLLRInputS3xD(274)(4) <= VNStageIntLLROutputS2xD(259)(2);
  CNStageIntLLRInputS3xD(303)(4) <= VNStageIntLLROutputS2xD(259)(3);
  CNStageIntLLRInputS3xD(370)(4) <= VNStageIntLLROutputS2xD(259)(4);
  CNStageIntLLRInputS3xD(49)(4) <= VNStageIntLLROutputS2xD(260)(0);
  CNStageIntLLRInputS3xD(71)(4) <= VNStageIntLLROutputS2xD(260)(1);
  CNStageIntLLRInputS3xD(138)(4) <= VNStageIntLLROutputS2xD(260)(2);
  CNStageIntLLRInputS3xD(186)(4) <= VNStageIntLLROutputS2xD(260)(3);
  CNStageIntLLRInputS3xD(243)(4) <= VNStageIntLLROutputS2xD(260)(4);
  CNStageIntLLRInputS3xD(383)(4) <= VNStageIntLLROutputS2xD(260)(5);
  CNStageIntLLRInputS3xD(48)(4) <= VNStageIntLLROutputS2xD(261)(0);
  CNStageIntLLRInputS3xD(63)(4) <= VNStageIntLLROutputS2xD(261)(1);
  CNStageIntLLRInputS3xD(152)(4) <= VNStageIntLLROutputS2xD(261)(2);
  CNStageIntLLRInputS3xD(204)(4) <= VNStageIntLLROutputS2xD(261)(3);
  CNStageIntLLRInputS3xD(305)(4) <= VNStageIntLLROutputS2xD(261)(4);
  CNStageIntLLRInputS3xD(333)(4) <= VNStageIntLLROutputS2xD(261)(5);
  CNStageIntLLRInputS3xD(47)(4) <= VNStageIntLLROutputS2xD(262)(0);
  CNStageIntLLRInputS3xD(95)(4) <= VNStageIntLLROutputS2xD(262)(1);
  CNStageIntLLRInputS3xD(149)(4) <= VNStageIntLLROutputS2xD(262)(2);
  CNStageIntLLRInputS3xD(212)(4) <= VNStageIntLLROutputS2xD(262)(3);
  CNStageIntLLRInputS3xD(319)(4) <= VNStageIntLLROutputS2xD(262)(4);
  CNStageIntLLRInputS3xD(362)(4) <= VNStageIntLLROutputS2xD(262)(5);
  CNStageIntLLRInputS3xD(46)(4) <= VNStageIntLLROutputS2xD(263)(0);
  CNStageIntLLRInputS3xD(104)(4) <= VNStageIntLLROutputS2xD(263)(1);
  CNStageIntLLRInputS3xD(169)(4) <= VNStageIntLLROutputS2xD(263)(2);
  CNStageIntLLRInputS3xD(207)(4) <= VNStageIntLLROutputS2xD(263)(3);
  CNStageIntLLRInputS3xD(253)(4) <= VNStageIntLLROutputS2xD(263)(4);
  CNStageIntLLRInputS3xD(315)(4) <= VNStageIntLLROutputS2xD(263)(5);
  CNStageIntLLRInputS3xD(378)(4) <= VNStageIntLLROutputS2xD(263)(6);
  CNStageIntLLRInputS3xD(45)(4) <= VNStageIntLLROutputS2xD(264)(0);
  CNStageIntLLRInputS3xD(98)(4) <= VNStageIntLLROutputS2xD(264)(1);
  CNStageIntLLRInputS3xD(132)(4) <= VNStageIntLLROutputS2xD(264)(2);
  CNStageIntLLRInputS3xD(213)(4) <= VNStageIntLLROutputS2xD(264)(3);
  CNStageIntLLRInputS3xD(256)(4) <= VNStageIntLLROutputS2xD(264)(4);
  CNStageIntLLRInputS3xD(281)(4) <= VNStageIntLLROutputS2xD(264)(5);
  CNStageIntLLRInputS3xD(349)(4) <= VNStageIntLLROutputS2xD(264)(6);
  CNStageIntLLRInputS3xD(44)(4) <= VNStageIntLLROutputS2xD(265)(0);
  CNStageIntLLRInputS3xD(133)(4) <= VNStageIntLLROutputS2xD(265)(1);
  CNStageIntLLRInputS3xD(203)(4) <= VNStageIntLLROutputS2xD(265)(2);
  CNStageIntLLRInputS3xD(244)(4) <= VNStageIntLLROutputS2xD(265)(3);
  CNStageIntLLRInputS3xD(43)(4) <= VNStageIntLLROutputS2xD(266)(0);
  CNStageIntLLRInputS3xD(168)(4) <= VNStageIntLLROutputS2xD(266)(1);
  CNStageIntLLRInputS3xD(173)(4) <= VNStageIntLLROutputS2xD(266)(2);
  CNStageIntLLRInputS3xD(273)(4) <= VNStageIntLLROutputS2xD(266)(3);
  CNStageIntLLRInputS3xD(300)(4) <= VNStageIntLLROutputS2xD(266)(4);
  CNStageIntLLRInputS3xD(42)(4) <= VNStageIntLLROutputS2xD(267)(0);
  CNStageIntLLRInputS3xD(72)(4) <= VNStageIntLLROutputS2xD(267)(1);
  CNStageIntLLRInputS3xD(159)(4) <= VNStageIntLLROutputS2xD(267)(2);
  CNStageIntLLRInputS3xD(180)(4) <= VNStageIntLLROutputS2xD(267)(3);
  CNStageIntLLRInputS3xD(241)(4) <= VNStageIntLLROutputS2xD(267)(4);
  CNStageIntLLRInputS3xD(280)(4) <= VNStageIntLLROutputS2xD(267)(5);
  CNStageIntLLRInputS3xD(364)(4) <= VNStageIntLLROutputS2xD(267)(6);
  CNStageIntLLRInputS3xD(41)(4) <= VNStageIntLLROutputS2xD(268)(0);
  CNStageIntLLRInputS3xD(109)(4) <= VNStageIntLLROutputS2xD(268)(1);
  CNStageIntLLRInputS3xD(118)(4) <= VNStageIntLLROutputS2xD(268)(2);
  CNStageIntLLRInputS3xD(216)(4) <= VNStageIntLLROutputS2xD(268)(3);
  CNStageIntLLRInputS3xD(266)(4) <= VNStageIntLLROutputS2xD(268)(4);
  CNStageIntLLRInputS3xD(325)(4) <= VNStageIntLLROutputS2xD(268)(5);
  CNStageIntLLRInputS3xD(360)(4) <= VNStageIntLLROutputS2xD(268)(6);
  CNStageIntLLRInputS3xD(67)(4) <= VNStageIntLLROutputS2xD(269)(0);
  CNStageIntLLRInputS3xD(122)(4) <= VNStageIntLLROutputS2xD(269)(1);
  CNStageIntLLRInputS3xD(218)(4) <= VNStageIntLLROutputS2xD(269)(2);
  CNStageIntLLRInputS3xD(250)(4) <= VNStageIntLLROutputS2xD(269)(3);
  CNStageIntLLRInputS3xD(287)(4) <= VNStageIntLLROutputS2xD(269)(4);
  CNStageIntLLRInputS3xD(381)(4) <= VNStageIntLLROutputS2xD(269)(5);
  CNStageIntLLRInputS3xD(40)(4) <= VNStageIntLLROutputS2xD(270)(0);
  CNStageIntLLRInputS3xD(79)(4) <= VNStageIntLLROutputS2xD(270)(1);
  CNStageIntLLRInputS3xD(170)(4) <= VNStageIntLLROutputS2xD(270)(2);
  CNStageIntLLRInputS3xD(190)(4) <= VNStageIntLLROutputS2xD(270)(3);
  CNStageIntLLRInputS3xD(275)(4) <= VNStageIntLLROutputS2xD(270)(4);
  CNStageIntLLRInputS3xD(292)(4) <= VNStageIntLLROutputS2xD(270)(5);
  CNStageIntLLRInputS3xD(344)(4) <= VNStageIntLLROutputS2xD(270)(6);
  CNStageIntLLRInputS3xD(39)(4) <= VNStageIntLLROutputS2xD(271)(0);
  CNStageIntLLRInputS3xD(105)(4) <= VNStageIntLLROutputS2xD(271)(1);
  CNStageIntLLRInputS3xD(171)(4) <= VNStageIntLLROutputS2xD(271)(2);
  CNStageIntLLRInputS3xD(268)(4) <= VNStageIntLLROutputS2xD(271)(3);
  CNStageIntLLRInputS3xD(332)(4) <= VNStageIntLLROutputS2xD(271)(4);
  CNStageIntLLRInputS3xD(345)(4) <= VNStageIntLLROutputS2xD(271)(5);
  CNStageIntLLRInputS3xD(38)(4) <= VNStageIntLLROutputS2xD(272)(0);
  CNStageIntLLRInputS3xD(94)(4) <= VNStageIntLLROutputS2xD(272)(1);
  CNStageIntLLRInputS3xD(116)(4) <= VNStageIntLLROutputS2xD(272)(2);
  CNStageIntLLRInputS3xD(184)(4) <= VNStageIntLLROutputS2xD(272)(3);
  CNStageIntLLRInputS3xD(254)(4) <= VNStageIntLLROutputS2xD(272)(4);
  CNStageIntLLRInputS3xD(291)(4) <= VNStageIntLLROutputS2xD(272)(5);
  CNStageIntLLRInputS3xD(380)(4) <= VNStageIntLLROutputS2xD(272)(6);
  CNStageIntLLRInputS3xD(37)(4) <= VNStageIntLLROutputS2xD(273)(0);
  CNStageIntLLRInputS3xD(81)(4) <= VNStageIntLLROutputS2xD(273)(1);
  CNStageIntLLRInputS3xD(156)(4) <= VNStageIntLLROutputS2xD(273)(2);
  CNStageIntLLRInputS3xD(272)(4) <= VNStageIntLLROutputS2xD(273)(3);
  CNStageIntLLRInputS3xD(285)(4) <= VNStageIntLLROutputS2xD(273)(4);
  CNStageIntLLRInputS3xD(371)(4) <= VNStageIntLLROutputS2xD(273)(5);
  CNStageIntLLRInputS3xD(36)(4) <= VNStageIntLLROutputS2xD(274)(0);
  CNStageIntLLRInputS3xD(164)(4) <= VNStageIntLLROutputS2xD(274)(1);
  CNStageIntLLRInputS3xD(217)(4) <= VNStageIntLLROutputS2xD(274)(2);
  CNStageIntLLRInputS3xD(248)(4) <= VNStageIntLLROutputS2xD(274)(3);
  CNStageIntLLRInputS3xD(35)(4) <= VNStageIntLLROutputS2xD(275)(0);
  CNStageIntLLRInputS3xD(59)(4) <= VNStageIntLLROutputS2xD(275)(1);
  CNStageIntLLRInputS3xD(128)(4) <= VNStageIntLLROutputS2xD(275)(2);
  CNStageIntLLRInputS3xD(179)(4) <= VNStageIntLLROutputS2xD(275)(3);
  CNStageIntLLRInputS3xD(329)(4) <= VNStageIntLLROutputS2xD(275)(4);
  CNStageIntLLRInputS3xD(34)(4) <= VNStageIntLLROutputS2xD(276)(0);
  CNStageIntLLRInputS3xD(69)(4) <= VNStageIntLLROutputS2xD(276)(1);
  CNStageIntLLRInputS3xD(126)(4) <= VNStageIntLLROutputS2xD(276)(2);
  CNStageIntLLRInputS3xD(205)(4) <= VNStageIntLLROutputS2xD(276)(3);
  CNStageIntLLRInputS3xD(259)(4) <= VNStageIntLLROutputS2xD(276)(4);
  CNStageIntLLRInputS3xD(297)(4) <= VNStageIntLLROutputS2xD(276)(5);
  CNStageIntLLRInputS3xD(33)(4) <= VNStageIntLLROutputS2xD(277)(0);
  CNStageIntLLRInputS3xD(64)(4) <= VNStageIntLLROutputS2xD(277)(1);
  CNStageIntLLRInputS3xD(162)(4) <= VNStageIntLLROutputS2xD(277)(2);
  CNStageIntLLRInputS3xD(185)(4) <= VNStageIntLLROutputS2xD(277)(3);
  CNStageIntLLRInputS3xD(252)(4) <= VNStageIntLLROutputS2xD(277)(4);
  CNStageIntLLRInputS3xD(295)(4) <= VNStageIntLLROutputS2xD(277)(5);
  CNStageIntLLRInputS3xD(334)(4) <= VNStageIntLLROutputS2xD(277)(6);
  CNStageIntLLRInputS3xD(32)(4) <= VNStageIntLLROutputS2xD(278)(0);
  CNStageIntLLRInputS3xD(70)(4) <= VNStageIntLLROutputS2xD(278)(1);
  CNStageIntLLRInputS3xD(141)(4) <= VNStageIntLLROutputS2xD(278)(2);
  CNStageIntLLRInputS3xD(229)(4) <= VNStageIntLLROutputS2xD(278)(3);
  CNStageIntLLRInputS3xD(328)(4) <= VNStageIntLLROutputS2xD(278)(4);
  CNStageIntLLRInputS3xD(31)(4) <= VNStageIntLLROutputS2xD(279)(0);
  CNStageIntLLRInputS3xD(58)(4) <= VNStageIntLLROutputS2xD(279)(1);
  CNStageIntLLRInputS3xD(144)(4) <= VNStageIntLLROutputS2xD(279)(2);
  CNStageIntLLRInputS3xD(219)(4) <= VNStageIntLLROutputS2xD(279)(3);
  CNStageIntLLRInputS3xD(239)(4) <= VNStageIntLLROutputS2xD(279)(4);
  CNStageIntLLRInputS3xD(368)(4) <= VNStageIntLLROutputS2xD(279)(5);
  CNStageIntLLRInputS3xD(30)(4) <= VNStageIntLLROutputS2xD(280)(0);
  CNStageIntLLRInputS3xD(84)(4) <= VNStageIntLLROutputS2xD(280)(1);
  CNStageIntLLRInputS3xD(129)(4) <= VNStageIntLLROutputS2xD(280)(2);
  CNStageIntLLRInputS3xD(215)(4) <= VNStageIntLLROutputS2xD(280)(3);
  CNStageIntLLRInputS3xD(233)(4) <= VNStageIntLLROutputS2xD(280)(4);
  CNStageIntLLRInputS3xD(310)(4) <= VNStageIntLLROutputS2xD(280)(5);
  CNStageIntLLRInputS3xD(376)(4) <= VNStageIntLLROutputS2xD(280)(6);
  CNStageIntLLRInputS3xD(29)(4) <= VNStageIntLLROutputS2xD(281)(0);
  CNStageIntLLRInputS3xD(90)(4) <= VNStageIntLLROutputS2xD(281)(1);
  CNStageIntLLRInputS3xD(163)(4) <= VNStageIntLLROutputS2xD(281)(2);
  CNStageIntLLRInputS3xD(182)(4) <= VNStageIntLLROutputS2xD(281)(3);
  CNStageIntLLRInputS3xD(236)(4) <= VNStageIntLLROutputS2xD(281)(4);
  CNStageIntLLRInputS3xD(298)(4) <= VNStageIntLLROutputS2xD(281)(5);
  CNStageIntLLRInputS3xD(340)(4) <= VNStageIntLLROutputS2xD(281)(6);
  CNStageIntLLRInputS3xD(28)(4) <= VNStageIntLLROutputS2xD(282)(0);
  CNStageIntLLRInputS3xD(74)(4) <= VNStageIntLLROutputS2xD(282)(1);
  CNStageIntLLRInputS3xD(125)(4) <= VNStageIntLLROutputS2xD(282)(2);
  CNStageIntLLRInputS3xD(200)(4) <= VNStageIntLLROutputS2xD(282)(3);
  CNStageIntLLRInputS3xD(226)(4) <= VNStageIntLLROutputS2xD(282)(4);
  CNStageIntLLRInputS3xD(338)(4) <= VNStageIntLLROutputS2xD(282)(5);
  CNStageIntLLRInputS3xD(27)(4) <= VNStageIntLLROutputS2xD(283)(0);
  CNStageIntLLRInputS3xD(76)(4) <= VNStageIntLLROutputS2xD(283)(1);
  CNStageIntLLRInputS3xD(153)(4) <= VNStageIntLLROutputS2xD(283)(2);
  CNStageIntLLRInputS3xD(201)(4) <= VNStageIntLLROutputS2xD(283)(3);
  CNStageIntLLRInputS3xD(260)(4) <= VNStageIntLLROutputS2xD(283)(4);
  CNStageIntLLRInputS3xD(294)(4) <= VNStageIntLLROutputS2xD(283)(5);
  CNStageIntLLRInputS3xD(374)(4) <= VNStageIntLLROutputS2xD(283)(6);
  CNStageIntLLRInputS3xD(26)(4) <= VNStageIntLLROutputS2xD(284)(0);
  CNStageIntLLRInputS3xD(100)(4) <= VNStageIntLLROutputS2xD(284)(1);
  CNStageIntLLRInputS3xD(137)(4) <= VNStageIntLLROutputS2xD(284)(2);
  CNStageIntLLRInputS3xD(181)(4) <= VNStageIntLLROutputS2xD(284)(3);
  CNStageIntLLRInputS3xD(245)(4) <= VNStageIntLLROutputS2xD(284)(4);
  CNStageIntLLRInputS3xD(320)(4) <= VNStageIntLLROutputS2xD(284)(5);
  CNStageIntLLRInputS3xD(353)(4) <= VNStageIntLLROutputS2xD(284)(6);
  CNStageIntLLRInputS3xD(25)(4) <= VNStageIntLLROutputS2xD(285)(0);
  CNStageIntLLRInputS3xD(82)(4) <= VNStageIntLLROutputS2xD(285)(1);
  CNStageIntLLRInputS3xD(165)(4) <= VNStageIntLLROutputS2xD(285)(2);
  CNStageIntLLRInputS3xD(172)(4) <= VNStageIntLLROutputS2xD(285)(3);
  CNStageIntLLRInputS3xD(255)(4) <= VNStageIntLLROutputS2xD(285)(4);
  CNStageIntLLRInputS3xD(304)(4) <= VNStageIntLLROutputS2xD(285)(5);
  CNStageIntLLRInputS3xD(355)(4) <= VNStageIntLLROutputS2xD(285)(6);
  CNStageIntLLRInputS3xD(24)(4) <= VNStageIntLLROutputS2xD(286)(0);
  CNStageIntLLRInputS3xD(93)(4) <= VNStageIntLLROutputS2xD(286)(1);
  CNStageIntLLRInputS3xD(155)(4) <= VNStageIntLLROutputS2xD(286)(2);
  CNStageIntLLRInputS3xD(189)(4) <= VNStageIntLLROutputS2xD(286)(3);
  CNStageIntLLRInputS3xD(267)(4) <= VNStageIntLLROutputS2xD(286)(4);
  CNStageIntLLRInputS3xD(330)(4) <= VNStageIntLLROutputS2xD(286)(5);
  CNStageIntLLRInputS3xD(341)(4) <= VNStageIntLLROutputS2xD(286)(6);
  CNStageIntLLRInputS3xD(23)(4) <= VNStageIntLLROutputS2xD(287)(0);
  CNStageIntLLRInputS3xD(101)(4) <= VNStageIntLLROutputS2xD(287)(1);
  CNStageIntLLRInputS3xD(142)(4) <= VNStageIntLLROutputS2xD(287)(2);
  CNStageIntLLRInputS3xD(193)(4) <= VNStageIntLLROutputS2xD(287)(3);
  CNStageIntLLRInputS3xD(240)(4) <= VNStageIntLLROutputS2xD(287)(4);
  CNStageIntLLRInputS3xD(322)(4) <= VNStageIntLLROutputS2xD(287)(5);
  CNStageIntLLRInputS3xD(375)(4) <= VNStageIntLLROutputS2xD(287)(6);
  CNStageIntLLRInputS3xD(22)(4) <= VNStageIntLLROutputS2xD(288)(0);
  CNStageIntLLRInputS3xD(75)(4) <= VNStageIntLLROutputS2xD(288)(1);
  CNStageIntLLRInputS3xD(161)(4) <= VNStageIntLLROutputS2xD(288)(2);
  CNStageIntLLRInputS3xD(224)(4) <= VNStageIntLLROutputS2xD(288)(3);
  CNStageIntLLRInputS3xD(228)(4) <= VNStageIntLLROutputS2xD(288)(4);
  CNStageIntLLRInputS3xD(308)(4) <= VNStageIntLLROutputS2xD(288)(5);
  CNStageIntLLRInputS3xD(337)(4) <= VNStageIntLLROutputS2xD(288)(6);
  CNStageIntLLRInputS3xD(21)(4) <= VNStageIntLLROutputS2xD(289)(0);
  CNStageIntLLRInputS3xD(89)(4) <= VNStageIntLLROutputS2xD(289)(1);
  CNStageIntLLRInputS3xD(134)(4) <= VNStageIntLLROutputS2xD(289)(2);
  CNStageIntLLRInputS3xD(192)(4) <= VNStageIntLLROutputS2xD(289)(3);
  CNStageIntLLRInputS3xD(269)(4) <= VNStageIntLLROutputS2xD(289)(4);
  CNStageIntLLRInputS3xD(327)(4) <= VNStageIntLLROutputS2xD(289)(5);
  CNStageIntLLRInputS3xD(365)(4) <= VNStageIntLLROutputS2xD(289)(6);
  CNStageIntLLRInputS3xD(20)(4) <= VNStageIntLLROutputS2xD(290)(0);
  CNStageIntLLRInputS3xD(60)(4) <= VNStageIntLLROutputS2xD(290)(1);
  CNStageIntLLRInputS3xD(131)(4) <= VNStageIntLLROutputS2xD(290)(2);
  CNStageIntLLRInputS3xD(187)(4) <= VNStageIntLLROutputS2xD(290)(3);
  CNStageIntLLRInputS3xD(231)(4) <= VNStageIntLLROutputS2xD(290)(4);
  CNStageIntLLRInputS3xD(350)(4) <= VNStageIntLLROutputS2xD(290)(5);
  CNStageIntLLRInputS3xD(19)(4) <= VNStageIntLLROutputS2xD(291)(0);
  CNStageIntLLRInputS3xD(96)(4) <= VNStageIntLLROutputS2xD(291)(1);
  CNStageIntLLRInputS3xD(147)(4) <= VNStageIntLLROutputS2xD(291)(2);
  CNStageIntLLRInputS3xD(223)(4) <= VNStageIntLLROutputS2xD(291)(3);
  CNStageIntLLRInputS3xD(249)(4) <= VNStageIntLLROutputS2xD(291)(4);
  CNStageIntLLRInputS3xD(377)(4) <= VNStageIntLLROutputS2xD(291)(5);
  CNStageIntLLRInputS3xD(18)(4) <= VNStageIntLLROutputS2xD(292)(0);
  CNStageIntLLRInputS3xD(62)(4) <= VNStageIntLLROutputS2xD(292)(1);
  CNStageIntLLRInputS3xD(139)(4) <= VNStageIntLLROutputS2xD(292)(2);
  CNStageIntLLRInputS3xD(177)(4) <= VNStageIntLLROutputS2xD(292)(3);
  CNStageIntLLRInputS3xD(257)(4) <= VNStageIntLLROutputS2xD(292)(4);
  CNStageIntLLRInputS3xD(313)(4) <= VNStageIntLLROutputS2xD(292)(5);
  CNStageIntLLRInputS3xD(367)(4) <= VNStageIntLLROutputS2xD(292)(6);
  CNStageIntLLRInputS3xD(17)(4) <= VNStageIntLLROutputS2xD(293)(0);
  CNStageIntLLRInputS3xD(77)(4) <= VNStageIntLLROutputS2xD(293)(1);
  CNStageIntLLRInputS3xD(113)(4) <= VNStageIntLLROutputS2xD(293)(2);
  CNStageIntLLRInputS3xD(197)(4) <= VNStageIntLLROutputS2xD(293)(3);
  CNStageIntLLRInputS3xD(306)(4) <= VNStageIntLLROutputS2xD(293)(4);
  CNStageIntLLRInputS3xD(354)(4) <= VNStageIntLLROutputS2xD(293)(5);
  CNStageIntLLRInputS3xD(16)(4) <= VNStageIntLLROutputS2xD(294)(0);
  CNStageIntLLRInputS3xD(73)(4) <= VNStageIntLLROutputS2xD(294)(1);
  CNStageIntLLRInputS3xD(123)(4) <= VNStageIntLLROutputS2xD(294)(2);
  CNStageIntLLRInputS3xD(196)(4) <= VNStageIntLLROutputS2xD(294)(3);
  CNStageIntLLRInputS3xD(258)(4) <= VNStageIntLLROutputS2xD(294)(4);
  CNStageIntLLRInputS3xD(284)(4) <= VNStageIntLLROutputS2xD(294)(5);
  CNStageIntLLRInputS3xD(373)(4) <= VNStageIntLLROutputS2xD(294)(6);
  CNStageIntLLRInputS3xD(15)(4) <= VNStageIntLLROutputS2xD(295)(0);
  CNStageIntLLRInputS3xD(92)(4) <= VNStageIntLLROutputS2xD(295)(1);
  CNStageIntLLRInputS3xD(117)(4) <= VNStageIntLLROutputS2xD(295)(2);
  CNStageIntLLRInputS3xD(175)(4) <= VNStageIntLLROutputS2xD(295)(3);
  CNStageIntLLRInputS3xD(346)(4) <= VNStageIntLLROutputS2xD(295)(4);
  CNStageIntLLRInputS3xD(14)(4) <= VNStageIntLLROutputS2xD(296)(0);
  CNStageIntLLRInputS3xD(55)(4) <= VNStageIntLLROutputS2xD(296)(1);
  CNStageIntLLRInputS3xD(121)(4) <= VNStageIntLLROutputS2xD(296)(2);
  CNStageIntLLRInputS3xD(208)(4) <= VNStageIntLLROutputS2xD(296)(3);
  CNStageIntLLRInputS3xD(286)(4) <= VNStageIntLLROutputS2xD(296)(4);
  CNStageIntLLRInputS3xD(343)(4) <= VNStageIntLLROutputS2xD(296)(5);
  CNStageIntLLRInputS3xD(13)(4) <= VNStageIntLLROutputS2xD(297)(0);
  CNStageIntLLRInputS3xD(56)(4) <= VNStageIntLLROutputS2xD(297)(1);
  CNStageIntLLRInputS3xD(111)(4) <= VNStageIntLLROutputS2xD(297)(2);
  CNStageIntLLRInputS3xD(211)(4) <= VNStageIntLLROutputS2xD(297)(3);
  CNStageIntLLRInputS3xD(277)(4) <= VNStageIntLLROutputS2xD(297)(4);
  CNStageIntLLRInputS3xD(290)(4) <= VNStageIntLLROutputS2xD(297)(5);
  CNStageIntLLRInputS3xD(358)(4) <= VNStageIntLLROutputS2xD(297)(6);
  CNStageIntLLRInputS3xD(12)(4) <= VNStageIntLLROutputS2xD(298)(0);
  CNStageIntLLRInputS3xD(91)(4) <= VNStageIntLLROutputS2xD(298)(1);
  CNStageIntLLRInputS3xD(148)(4) <= VNStageIntLLROutputS2xD(298)(2);
  CNStageIntLLRInputS3xD(198)(4) <= VNStageIntLLROutputS2xD(298)(3);
  CNStageIntLLRInputS3xD(262)(4) <= VNStageIntLLROutputS2xD(298)(4);
  CNStageIntLLRInputS3xD(282)(4) <= VNStageIntLLROutputS2xD(298)(5);
  CNStageIntLLRInputS3xD(351)(4) <= VNStageIntLLROutputS2xD(298)(6);
  CNStageIntLLRInputS3xD(83)(4) <= VNStageIntLLROutputS2xD(299)(0);
  CNStageIntLLRInputS3xD(130)(4) <= VNStageIntLLROutputS2xD(299)(1);
  CNStageIntLLRInputS3xD(176)(4) <= VNStageIntLLROutputS2xD(299)(2);
  CNStageIntLLRInputS3xD(264)(4) <= VNStageIntLLROutputS2xD(299)(3);
  CNStageIntLLRInputS3xD(314)(4) <= VNStageIntLLROutputS2xD(299)(4);
  CNStageIntLLRInputS3xD(11)(4) <= VNStageIntLLROutputS2xD(300)(0);
  CNStageIntLLRInputS3xD(99)(4) <= VNStageIntLLROutputS2xD(300)(1);
  CNStageIntLLRInputS3xD(143)(4) <= VNStageIntLLROutputS2xD(300)(2);
  CNStageIntLLRInputS3xD(195)(4) <= VNStageIntLLROutputS2xD(300)(3);
  CNStageIntLLRInputS3xD(299)(4) <= VNStageIntLLROutputS2xD(300)(4);
  CNStageIntLLRInputS3xD(335)(4) <= VNStageIntLLROutputS2xD(300)(5);
  CNStageIntLLRInputS3xD(10)(4) <= VNStageIntLLROutputS2xD(301)(0);
  CNStageIntLLRInputS3xD(103)(4) <= VNStageIntLLROutputS2xD(301)(1);
  CNStageIntLLRInputS3xD(154)(4) <= VNStageIntLLROutputS2xD(301)(2);
  CNStageIntLLRInputS3xD(220)(4) <= VNStageIntLLROutputS2xD(301)(3);
  CNStageIntLLRInputS3xD(270)(4) <= VNStageIntLLROutputS2xD(301)(4);
  CNStageIntLLRInputS3xD(309)(4) <= VNStageIntLLROutputS2xD(301)(5);
  CNStageIntLLRInputS3xD(9)(4) <= VNStageIntLLROutputS2xD(302)(0);
  CNStageIntLLRInputS3xD(110)(4) <= VNStageIntLLROutputS2xD(302)(1);
  CNStageIntLLRInputS3xD(124)(4) <= VNStageIntLLROutputS2xD(302)(2);
  CNStageIntLLRInputS3xD(206)(4) <= VNStageIntLLROutputS2xD(302)(3);
  CNStageIntLLRInputS3xD(227)(4) <= VNStageIntLLROutputS2xD(302)(4);
  CNStageIntLLRInputS3xD(321)(4) <= VNStageIntLLROutputS2xD(302)(5);
  CNStageIntLLRInputS3xD(8)(4) <= VNStageIntLLROutputS2xD(303)(0);
  CNStageIntLLRInputS3xD(102)(4) <= VNStageIntLLROutputS2xD(303)(1);
  CNStageIntLLRInputS3xD(112)(4) <= VNStageIntLLROutputS2xD(303)(2);
  CNStageIntLLRInputS3xD(178)(4) <= VNStageIntLLROutputS2xD(303)(3);
  CNStageIntLLRInputS3xD(235)(4) <= VNStageIntLLROutputS2xD(303)(4);
  CNStageIntLLRInputS3xD(293)(4) <= VNStageIntLLROutputS2xD(303)(5);
  CNStageIntLLRInputS3xD(382)(4) <= VNStageIntLLROutputS2xD(303)(6);
  CNStageIntLLRInputS3xD(7)(4) <= VNStageIntLLROutputS2xD(304)(0);
  CNStageIntLLRInputS3xD(97)(4) <= VNStageIntLLROutputS2xD(304)(1);
  CNStageIntLLRInputS3xD(157)(4) <= VNStageIntLLROutputS2xD(304)(2);
  CNStageIntLLRInputS3xD(222)(4) <= VNStageIntLLROutputS2xD(304)(3);
  CNStageIntLLRInputS3xD(263)(4) <= VNStageIntLLROutputS2xD(304)(4);
  CNStageIntLLRInputS3xD(283)(4) <= VNStageIntLLROutputS2xD(304)(5);
  CNStageIntLLRInputS3xD(359)(4) <= VNStageIntLLROutputS2xD(304)(6);
  CNStageIntLLRInputS3xD(6)(4) <= VNStageIntLLROutputS2xD(305)(0);
  CNStageIntLLRInputS3xD(80)(4) <= VNStageIntLLROutputS2xD(305)(1);
  CNStageIntLLRInputS3xD(115)(4) <= VNStageIntLLROutputS2xD(305)(2);
  CNStageIntLLRInputS3xD(209)(4) <= VNStageIntLLROutputS2xD(305)(3);
  CNStageIntLLRInputS3xD(276)(4) <= VNStageIntLLROutputS2xD(305)(4);
  CNStageIntLLRInputS3xD(323)(4) <= VNStageIntLLROutputS2xD(305)(5);
  CNStageIntLLRInputS3xD(342)(4) <= VNStageIntLLROutputS2xD(305)(6);
  CNStageIntLLRInputS3xD(5)(4) <= VNStageIntLLROutputS2xD(306)(0);
  CNStageIntLLRInputS3xD(87)(4) <= VNStageIntLLROutputS2xD(306)(1);
  CNStageIntLLRInputS3xD(136)(4) <= VNStageIntLLROutputS2xD(306)(2);
  CNStageIntLLRInputS3xD(174)(4) <= VNStageIntLLROutputS2xD(306)(3);
  CNStageIntLLRInputS3xD(4)(4) <= VNStageIntLLROutputS2xD(307)(0);
  CNStageIntLLRInputS3xD(107)(4) <= VNStageIntLLROutputS2xD(307)(1);
  CNStageIntLLRInputS3xD(145)(4) <= VNStageIntLLROutputS2xD(307)(2);
  CNStageIntLLRInputS3xD(202)(4) <= VNStageIntLLROutputS2xD(307)(3);
  CNStageIntLLRInputS3xD(230)(4) <= VNStageIntLLROutputS2xD(307)(4);
  CNStageIntLLRInputS3xD(302)(4) <= VNStageIntLLROutputS2xD(307)(5);
  CNStageIntLLRInputS3xD(366)(4) <= VNStageIntLLROutputS2xD(307)(6);
  CNStageIntLLRInputS3xD(140)(4) <= VNStageIntLLROutputS2xD(308)(0);
  CNStageIntLLRInputS3xD(199)(4) <= VNStageIntLLROutputS2xD(308)(1);
  CNStageIntLLRInputS3xD(251)(4) <= VNStageIntLLROutputS2xD(308)(2);
  CNStageIntLLRInputS3xD(311)(4) <= VNStageIntLLROutputS2xD(308)(3);
  CNStageIntLLRInputS3xD(336)(4) <= VNStageIntLLROutputS2xD(308)(4);
  CNStageIntLLRInputS3xD(3)(4) <= VNStageIntLLROutputS2xD(309)(0);
  CNStageIntLLRInputS3xD(86)(4) <= VNStageIntLLROutputS2xD(309)(1);
  CNStageIntLLRInputS3xD(146)(4) <= VNStageIntLLROutputS2xD(309)(2);
  CNStageIntLLRInputS3xD(214)(4) <= VNStageIntLLROutputS2xD(309)(3);
  CNStageIntLLRInputS3xD(265)(4) <= VNStageIntLLROutputS2xD(309)(4);
  CNStageIntLLRInputS3xD(307)(4) <= VNStageIntLLROutputS2xD(309)(5);
  CNStageIntLLRInputS3xD(2)(4) <= VNStageIntLLROutputS2xD(310)(0);
  CNStageIntLLRInputS3xD(65)(4) <= VNStageIntLLROutputS2xD(310)(1);
  CNStageIntLLRInputS3xD(135)(4) <= VNStageIntLLROutputS2xD(310)(2);
  CNStageIntLLRInputS3xD(261)(4) <= VNStageIntLLROutputS2xD(310)(3);
  CNStageIntLLRInputS3xD(312)(4) <= VNStageIntLLROutputS2xD(310)(4);
  CNStageIntLLRInputS3xD(369)(4) <= VNStageIntLLROutputS2xD(310)(5);
  CNStageIntLLRInputS3xD(1)(4) <= VNStageIntLLROutputS2xD(311)(0);
  CNStageIntLLRInputS3xD(68)(4) <= VNStageIntLLROutputS2xD(311)(1);
  CNStageIntLLRInputS3xD(160)(4) <= VNStageIntLLROutputS2xD(311)(2);
  CNStageIntLLRInputS3xD(225)(4) <= VNStageIntLLROutputS2xD(311)(3);
  CNStageIntLLRInputS3xD(301)(4) <= VNStageIntLLROutputS2xD(311)(4);
  CNStageIntLLRInputS3xD(0)(4) <= VNStageIntLLROutputS2xD(312)(0);
  CNStageIntLLRInputS3xD(108)(4) <= VNStageIntLLROutputS2xD(312)(1);
  CNStageIntLLRInputS3xD(167)(4) <= VNStageIntLLROutputS2xD(312)(2);
  CNStageIntLLRInputS3xD(246)(4) <= VNStageIntLLROutputS2xD(312)(3);
  CNStageIntLLRInputS3xD(326)(4) <= VNStageIntLLROutputS2xD(312)(4);
  CNStageIntLLRInputS3xD(348)(4) <= VNStageIntLLROutputS2xD(312)(5);
  CNStageIntLLRInputS3xD(150)(4) <= VNStageIntLLROutputS2xD(313)(0);
  CNStageIntLLRInputS3xD(188)(4) <= VNStageIntLLROutputS2xD(313)(1);
  CNStageIntLLRInputS3xD(247)(4) <= VNStageIntLLROutputS2xD(313)(2);
  CNStageIntLLRInputS3xD(356)(4) <= VNStageIntLLROutputS2xD(313)(3);
  CNStageIntLLRInputS3xD(191)(4) <= VNStageIntLLROutputS2xD(314)(0);
  CNStageIntLLRInputS3xD(278)(4) <= VNStageIntLLROutputS2xD(314)(1);
  CNStageIntLLRInputS3xD(316)(4) <= VNStageIntLLROutputS2xD(314)(2);
  CNStageIntLLRInputS3xD(352)(4) <= VNStageIntLLROutputS2xD(314)(3);
  CNStageIntLLRInputS3xD(78)(4) <= VNStageIntLLROutputS2xD(315)(0);
  CNStageIntLLRInputS3xD(119)(4) <= VNStageIntLLROutputS2xD(315)(1);
  CNStageIntLLRInputS3xD(183)(4) <= VNStageIntLLROutputS2xD(315)(2);
  CNStageIntLLRInputS3xD(271)(4) <= VNStageIntLLROutputS2xD(315)(3);
  CNStageIntLLRInputS3xD(318)(4) <= VNStageIntLLROutputS2xD(315)(4);
  CNStageIntLLRInputS3xD(357)(4) <= VNStageIntLLROutputS2xD(315)(5);
  CNStageIntLLRInputS3xD(61)(4) <= VNStageIntLLROutputS2xD(316)(0);
  CNStageIntLLRInputS3xD(158)(4) <= VNStageIntLLROutputS2xD(316)(1);
  CNStageIntLLRInputS3xD(234)(4) <= VNStageIntLLROutputS2xD(316)(2);
  CNStageIntLLRInputS3xD(288)(4) <= VNStageIntLLROutputS2xD(316)(3);
  CNStageIntLLRInputS3xD(347)(4) <= VNStageIntLLROutputS2xD(316)(4);
  CNStageIntLLRInputS3xD(88)(4) <= VNStageIntLLROutputS2xD(317)(0);
  CNStageIntLLRInputS3xD(238)(4) <= VNStageIntLLROutputS2xD(317)(1);
  CNStageIntLLRInputS3xD(324)(4) <= VNStageIntLLROutputS2xD(317)(2);
  CNStageIntLLRInputS3xD(372)(4) <= VNStageIntLLROutputS2xD(317)(3);
  CNStageIntLLRInputS3xD(120)(4) <= VNStageIntLLROutputS2xD(318)(0);
  CNStageIntLLRInputS3xD(210)(4) <= VNStageIntLLROutputS2xD(318)(1);
  CNStageIntLLRInputS3xD(279)(4) <= VNStageIntLLROutputS2xD(318)(2);
  CNStageIntLLRInputS3xD(379)(4) <= VNStageIntLLROutputS2xD(318)(3);
  CNStageIntLLRInputS3xD(52)(4) <= VNStageIntLLROutputS2xD(319)(0);
  CNStageIntLLRInputS3xD(66)(4) <= VNStageIntLLROutputS2xD(319)(1);
  CNStageIntLLRInputS3xD(151)(4) <= VNStageIntLLROutputS2xD(319)(2);
  CNStageIntLLRInputS3xD(221)(4) <= VNStageIntLLROutputS2xD(319)(3);
  CNStageIntLLRInputS3xD(237)(4) <= VNStageIntLLROutputS2xD(319)(4);
  CNStageIntLLRInputS3xD(289)(4) <= VNStageIntLLROutputS2xD(319)(5);
  CNStageIntLLRInputS3xD(361)(4) <= VNStageIntLLROutputS2xD(319)(6);
  CNStageIntLLRInputS3xD(53)(5) <= VNStageIntLLROutputS2xD(320)(0);
  CNStageIntLLRInputS3xD(126)(5) <= VNStageIntLLROutputS2xD(320)(1);
  CNStageIntLLRInputS3xD(196)(5) <= VNStageIntLLROutputS2xD(320)(2);
  CNStageIntLLRInputS3xD(295)(5) <= VNStageIntLLROutputS2xD(320)(3);
  CNStageIntLLRInputS3xD(338)(5) <= VNStageIntLLROutputS2xD(320)(4);
  CNStageIntLLRInputS3xD(51)(5) <= VNStageIntLLROutputS2xD(321)(0);
  CNStageIntLLRInputS3xD(65)(5) <= VNStageIntLLROutputS2xD(321)(1);
  CNStageIntLLRInputS3xD(150)(5) <= VNStageIntLLROutputS2xD(321)(2);
  CNStageIntLLRInputS3xD(220)(5) <= VNStageIntLLROutputS2xD(321)(3);
  CNStageIntLLRInputS3xD(236)(5) <= VNStageIntLLROutputS2xD(321)(4);
  CNStageIntLLRInputS3xD(288)(5) <= VNStageIntLLROutputS2xD(321)(5);
  CNStageIntLLRInputS3xD(360)(5) <= VNStageIntLLROutputS2xD(321)(6);
  CNStageIntLLRInputS3xD(50)(5) <= VNStageIntLLROutputS2xD(322)(0);
  CNStageIntLLRInputS3xD(84)(5) <= VNStageIntLLROutputS2xD(322)(1);
  CNStageIntLLRInputS3xD(165)(5) <= VNStageIntLLROutputS2xD(322)(2);
  CNStageIntLLRInputS3xD(231)(5) <= VNStageIntLLROutputS2xD(322)(3);
  CNStageIntLLRInputS3xD(316)(5) <= VNStageIntLLROutputS2xD(322)(4);
  CNStageIntLLRInputS3xD(362)(5) <= VNStageIntLLROutputS2xD(322)(5);
  CNStageIntLLRInputS3xD(56)(5) <= VNStageIntLLROutputS2xD(323)(0);
  CNStageIntLLRInputS3xD(136)(5) <= VNStageIntLLROutputS2xD(323)(1);
  CNStageIntLLRInputS3xD(184)(5) <= VNStageIntLLROutputS2xD(323)(2);
  CNStageIntLLRInputS3xD(268)(5) <= VNStageIntLLROutputS2xD(323)(3);
  CNStageIntLLRInputS3xD(330)(5) <= VNStageIntLLROutputS2xD(323)(4);
  CNStageIntLLRInputS3xD(49)(5) <= VNStageIntLLROutputS2xD(324)(0);
  CNStageIntLLRInputS3xD(109)(5) <= VNStageIntLLROutputS2xD(324)(1);
  CNStageIntLLRInputS3xD(113)(5) <= VNStageIntLLROutputS2xD(324)(2);
  CNStageIntLLRInputS3xD(223)(5) <= VNStageIntLLROutputS2xD(324)(3);
  CNStageIntLLRInputS3xD(273)(5) <= VNStageIntLLROutputS2xD(324)(4);
  CNStageIntLLRInputS3xD(302)(5) <= VNStageIntLLROutputS2xD(324)(5);
  CNStageIntLLRInputS3xD(369)(5) <= VNStageIntLLROutputS2xD(324)(6);
  CNStageIntLLRInputS3xD(48)(5) <= VNStageIntLLROutputS2xD(325)(0);
  CNStageIntLLRInputS3xD(70)(5) <= VNStageIntLLROutputS2xD(325)(1);
  CNStageIntLLRInputS3xD(137)(5) <= VNStageIntLLROutputS2xD(325)(2);
  CNStageIntLLRInputS3xD(185)(5) <= VNStageIntLLROutputS2xD(325)(3);
  CNStageIntLLRInputS3xD(242)(5) <= VNStageIntLLROutputS2xD(325)(4);
  CNStageIntLLRInputS3xD(284)(5) <= VNStageIntLLROutputS2xD(325)(5);
  CNStageIntLLRInputS3xD(382)(5) <= VNStageIntLLROutputS2xD(325)(6);
  CNStageIntLLRInputS3xD(47)(5) <= VNStageIntLLROutputS2xD(326)(0);
  CNStageIntLLRInputS3xD(62)(5) <= VNStageIntLLROutputS2xD(326)(1);
  CNStageIntLLRInputS3xD(203)(5) <= VNStageIntLLROutputS2xD(326)(2);
  CNStageIntLLRInputS3xD(241)(5) <= VNStageIntLLROutputS2xD(326)(3);
  CNStageIntLLRInputS3xD(304)(5) <= VNStageIntLLROutputS2xD(326)(4);
  CNStageIntLLRInputS3xD(46)(5) <= VNStageIntLLROutputS2xD(327)(0);
  CNStageIntLLRInputS3xD(94)(5) <= VNStageIntLLROutputS2xD(327)(1);
  CNStageIntLLRInputS3xD(148)(5) <= VNStageIntLLROutputS2xD(327)(2);
  CNStageIntLLRInputS3xD(211)(5) <= VNStageIntLLROutputS2xD(327)(3);
  CNStageIntLLRInputS3xD(272)(5) <= VNStageIntLLROutputS2xD(327)(4);
  CNStageIntLLRInputS3xD(318)(5) <= VNStageIntLLROutputS2xD(327)(5);
  CNStageIntLLRInputS3xD(361)(5) <= VNStageIntLLROutputS2xD(327)(6);
  CNStageIntLLRInputS3xD(45)(5) <= VNStageIntLLROutputS2xD(328)(0);
  CNStageIntLLRInputS3xD(103)(5) <= VNStageIntLLROutputS2xD(328)(1);
  CNStageIntLLRInputS3xD(168)(5) <= VNStageIntLLROutputS2xD(328)(2);
  CNStageIntLLRInputS3xD(314)(5) <= VNStageIntLLROutputS2xD(328)(3);
  CNStageIntLLRInputS3xD(377)(5) <= VNStageIntLLROutputS2xD(328)(4);
  CNStageIntLLRInputS3xD(44)(5) <= VNStageIntLLROutputS2xD(329)(0);
  CNStageIntLLRInputS3xD(97)(5) <= VNStageIntLLROutputS2xD(329)(1);
  CNStageIntLLRInputS3xD(131)(5) <= VNStageIntLLROutputS2xD(329)(2);
  CNStageIntLLRInputS3xD(212)(5) <= VNStageIntLLROutputS2xD(329)(3);
  CNStageIntLLRInputS3xD(255)(5) <= VNStageIntLLROutputS2xD(329)(4);
  CNStageIntLLRInputS3xD(280)(5) <= VNStageIntLLROutputS2xD(329)(5);
  CNStageIntLLRInputS3xD(348)(5) <= VNStageIntLLROutputS2xD(329)(6);
  CNStageIntLLRInputS3xD(43)(5) <= VNStageIntLLROutputS2xD(330)(0);
  CNStageIntLLRInputS3xD(101)(5) <= VNStageIntLLROutputS2xD(330)(1);
  CNStageIntLLRInputS3xD(132)(5) <= VNStageIntLLROutputS2xD(330)(2);
  CNStageIntLLRInputS3xD(202)(5) <= VNStageIntLLROutputS2xD(330)(3);
  CNStageIntLLRInputS3xD(243)(5) <= VNStageIntLLROutputS2xD(330)(4);
  CNStageIntLLRInputS3xD(42)(5) <= VNStageIntLLROutputS2xD(331)(0);
  CNStageIntLLRInputS3xD(92)(5) <= VNStageIntLLROutputS2xD(331)(1);
  CNStageIntLLRInputS3xD(167)(5) <= VNStageIntLLROutputS2xD(331)(2);
  CNStageIntLLRInputS3xD(172)(5) <= VNStageIntLLROutputS2xD(331)(3);
  CNStageIntLLRInputS3xD(350)(5) <= VNStageIntLLROutputS2xD(331)(4);
  CNStageIntLLRInputS3xD(41)(5) <= VNStageIntLLROutputS2xD(332)(0);
  CNStageIntLLRInputS3xD(71)(5) <= VNStageIntLLROutputS2xD(332)(1);
  CNStageIntLLRInputS3xD(158)(5) <= VNStageIntLLROutputS2xD(332)(2);
  CNStageIntLLRInputS3xD(179)(5) <= VNStageIntLLROutputS2xD(332)(3);
  CNStageIntLLRInputS3xD(240)(5) <= VNStageIntLLROutputS2xD(332)(4);
  CNStageIntLLRInputS3xD(363)(5) <= VNStageIntLLROutputS2xD(332)(5);
  CNStageIntLLRInputS3xD(108)(5) <= VNStageIntLLROutputS2xD(333)(0);
  CNStageIntLLRInputS3xD(117)(5) <= VNStageIntLLROutputS2xD(333)(1);
  CNStageIntLLRInputS3xD(215)(5) <= VNStageIntLLROutputS2xD(333)(2);
  CNStageIntLLRInputS3xD(265)(5) <= VNStageIntLLROutputS2xD(333)(3);
  CNStageIntLLRInputS3xD(324)(5) <= VNStageIntLLROutputS2xD(333)(4);
  CNStageIntLLRInputS3xD(359)(5) <= VNStageIntLLROutputS2xD(333)(5);
  CNStageIntLLRInputS3xD(40)(5) <= VNStageIntLLROutputS2xD(334)(0);
  CNStageIntLLRInputS3xD(66)(5) <= VNStageIntLLROutputS2xD(334)(1);
  CNStageIntLLRInputS3xD(217)(5) <= VNStageIntLLROutputS2xD(334)(2);
  CNStageIntLLRInputS3xD(286)(5) <= VNStageIntLLROutputS2xD(334)(3);
  CNStageIntLLRInputS3xD(380)(5) <= VNStageIntLLROutputS2xD(334)(4);
  CNStageIntLLRInputS3xD(39)(5) <= VNStageIntLLROutputS2xD(335)(0);
  CNStageIntLLRInputS3xD(78)(5) <= VNStageIntLLROutputS2xD(335)(1);
  CNStageIntLLRInputS3xD(170)(5) <= VNStageIntLLROutputS2xD(335)(2);
  CNStageIntLLRInputS3xD(189)(5) <= VNStageIntLLROutputS2xD(335)(3);
  CNStageIntLLRInputS3xD(274)(5) <= VNStageIntLLROutputS2xD(335)(4);
  CNStageIntLLRInputS3xD(291)(5) <= VNStageIntLLROutputS2xD(335)(5);
  CNStageIntLLRInputS3xD(343)(5) <= VNStageIntLLROutputS2xD(335)(6);
  CNStageIntLLRInputS3xD(38)(5) <= VNStageIntLLROutputS2xD(336)(0);
  CNStageIntLLRInputS3xD(104)(5) <= VNStageIntLLROutputS2xD(336)(1);
  CNStageIntLLRInputS3xD(121)(5) <= VNStageIntLLROutputS2xD(336)(2);
  CNStageIntLLRInputS3xD(267)(5) <= VNStageIntLLROutputS2xD(336)(3);
  CNStageIntLLRInputS3xD(332)(5) <= VNStageIntLLROutputS2xD(336)(4);
  CNStageIntLLRInputS3xD(344)(5) <= VNStageIntLLROutputS2xD(336)(5);
  CNStageIntLLRInputS3xD(37)(5) <= VNStageIntLLROutputS2xD(337)(0);
  CNStageIntLLRInputS3xD(93)(5) <= VNStageIntLLROutputS2xD(337)(1);
  CNStageIntLLRInputS3xD(115)(5) <= VNStageIntLLROutputS2xD(337)(2);
  CNStageIntLLRInputS3xD(183)(5) <= VNStageIntLLROutputS2xD(337)(3);
  CNStageIntLLRInputS3xD(253)(5) <= VNStageIntLLROutputS2xD(337)(4);
  CNStageIntLLRInputS3xD(290)(5) <= VNStageIntLLROutputS2xD(337)(5);
  CNStageIntLLRInputS3xD(379)(5) <= VNStageIntLLROutputS2xD(337)(6);
  CNStageIntLLRInputS3xD(36)(5) <= VNStageIntLLROutputS2xD(338)(0);
  CNStageIntLLRInputS3xD(80)(5) <= VNStageIntLLROutputS2xD(338)(1);
  CNStageIntLLRInputS3xD(155)(5) <= VNStageIntLLROutputS2xD(338)(2);
  CNStageIntLLRInputS3xD(190)(5) <= VNStageIntLLROutputS2xD(338)(3);
  CNStageIntLLRInputS3xD(370)(5) <= VNStageIntLLROutputS2xD(338)(4);
  CNStageIntLLRInputS3xD(35)(5) <= VNStageIntLLROutputS2xD(339)(0);
  CNStageIntLLRInputS3xD(96)(5) <= VNStageIntLLROutputS2xD(339)(1);
  CNStageIntLLRInputS3xD(163)(5) <= VNStageIntLLROutputS2xD(339)(2);
  CNStageIntLLRInputS3xD(216)(5) <= VNStageIntLLROutputS2xD(339)(3);
  CNStageIntLLRInputS3xD(247)(5) <= VNStageIntLLROutputS2xD(339)(4);
  CNStageIntLLRInputS3xD(322)(5) <= VNStageIntLLROutputS2xD(339)(5);
  CNStageIntLLRInputS3xD(34)(5) <= VNStageIntLLROutputS2xD(340)(0);
  CNStageIntLLRInputS3xD(58)(5) <= VNStageIntLLROutputS2xD(340)(1);
  CNStageIntLLRInputS3xD(127)(5) <= VNStageIntLLROutputS2xD(340)(2);
  CNStageIntLLRInputS3xD(178)(5) <= VNStageIntLLROutputS2xD(340)(3);
  CNStageIntLLRInputS3xD(245)(5) <= VNStageIntLLROutputS2xD(340)(4);
  CNStageIntLLRInputS3xD(334)(5) <= VNStageIntLLROutputS2xD(340)(5);
  CNStageIntLLRInputS3xD(33)(5) <= VNStageIntLLROutputS2xD(341)(0);
  CNStageIntLLRInputS3xD(68)(5) <= VNStageIntLLROutputS2xD(341)(1);
  CNStageIntLLRInputS3xD(125)(5) <= VNStageIntLLROutputS2xD(341)(2);
  CNStageIntLLRInputS3xD(204)(5) <= VNStageIntLLROutputS2xD(341)(3);
  CNStageIntLLRInputS3xD(258)(5) <= VNStageIntLLROutputS2xD(341)(4);
  CNStageIntLLRInputS3xD(296)(5) <= VNStageIntLLROutputS2xD(341)(5);
  CNStageIntLLRInputS3xD(32)(5) <= VNStageIntLLROutputS2xD(342)(0);
  CNStageIntLLRInputS3xD(63)(5) <= VNStageIntLLROutputS2xD(342)(1);
  CNStageIntLLRInputS3xD(161)(5) <= VNStageIntLLROutputS2xD(342)(2);
  CNStageIntLLRInputS3xD(251)(5) <= VNStageIntLLROutputS2xD(342)(3);
  CNStageIntLLRInputS3xD(294)(5) <= VNStageIntLLROutputS2xD(342)(4);
  CNStageIntLLRInputS3xD(31)(5) <= VNStageIntLLROutputS2xD(343)(0);
  CNStageIntLLRInputS3xD(69)(5) <= VNStageIntLLROutputS2xD(343)(1);
  CNStageIntLLRInputS3xD(140)(5) <= VNStageIntLLROutputS2xD(343)(2);
  CNStageIntLLRInputS3xD(206)(5) <= VNStageIntLLROutputS2xD(343)(3);
  CNStageIntLLRInputS3xD(228)(5) <= VNStageIntLLROutputS2xD(343)(4);
  CNStageIntLLRInputS3xD(327)(5) <= VNStageIntLLROutputS2xD(343)(5);
  CNStageIntLLRInputS3xD(30)(5) <= VNStageIntLLROutputS2xD(344)(0);
  CNStageIntLLRInputS3xD(57)(5) <= VNStageIntLLROutputS2xD(344)(1);
  CNStageIntLLRInputS3xD(143)(5) <= VNStageIntLLROutputS2xD(344)(2);
  CNStageIntLLRInputS3xD(218)(5) <= VNStageIntLLROutputS2xD(344)(3);
  CNStageIntLLRInputS3xD(238)(5) <= VNStageIntLLROutputS2xD(344)(4);
  CNStageIntLLRInputS3xD(307)(5) <= VNStageIntLLROutputS2xD(344)(5);
  CNStageIntLLRInputS3xD(367)(5) <= VNStageIntLLROutputS2xD(344)(6);
  CNStageIntLLRInputS3xD(29)(5) <= VNStageIntLLROutputS2xD(345)(0);
  CNStageIntLLRInputS3xD(83)(5) <= VNStageIntLLROutputS2xD(345)(1);
  CNStageIntLLRInputS3xD(128)(5) <= VNStageIntLLROutputS2xD(345)(2);
  CNStageIntLLRInputS3xD(232)(5) <= VNStageIntLLROutputS2xD(345)(3);
  CNStageIntLLRInputS3xD(309)(5) <= VNStageIntLLROutputS2xD(345)(4);
  CNStageIntLLRInputS3xD(375)(5) <= VNStageIntLLROutputS2xD(345)(5);
  CNStageIntLLRInputS3xD(28)(5) <= VNStageIntLLROutputS2xD(346)(0);
  CNStageIntLLRInputS3xD(89)(5) <= VNStageIntLLROutputS2xD(346)(1);
  CNStageIntLLRInputS3xD(162)(5) <= VNStageIntLLROutputS2xD(346)(2);
  CNStageIntLLRInputS3xD(181)(5) <= VNStageIntLLROutputS2xD(346)(3);
  CNStageIntLLRInputS3xD(235)(5) <= VNStageIntLLROutputS2xD(346)(4);
  CNStageIntLLRInputS3xD(297)(5) <= VNStageIntLLROutputS2xD(346)(5);
  CNStageIntLLRInputS3xD(339)(5) <= VNStageIntLLROutputS2xD(346)(6);
  CNStageIntLLRInputS3xD(27)(5) <= VNStageIntLLROutputS2xD(347)(0);
  CNStageIntLLRInputS3xD(73)(5) <= VNStageIntLLROutputS2xD(347)(1);
  CNStageIntLLRInputS3xD(124)(5) <= VNStageIntLLROutputS2xD(347)(2);
  CNStageIntLLRInputS3xD(199)(5) <= VNStageIntLLROutputS2xD(347)(3);
  CNStageIntLLRInputS3xD(225)(5) <= VNStageIntLLROutputS2xD(347)(4);
  CNStageIntLLRInputS3xD(328)(5) <= VNStageIntLLROutputS2xD(347)(5);
  CNStageIntLLRInputS3xD(337)(5) <= VNStageIntLLROutputS2xD(347)(6);
  CNStageIntLLRInputS3xD(26)(5) <= VNStageIntLLROutputS2xD(348)(0);
  CNStageIntLLRInputS3xD(75)(5) <= VNStageIntLLROutputS2xD(348)(1);
  CNStageIntLLRInputS3xD(152)(5) <= VNStageIntLLROutputS2xD(348)(2);
  CNStageIntLLRInputS3xD(200)(5) <= VNStageIntLLROutputS2xD(348)(3);
  CNStageIntLLRInputS3xD(259)(5) <= VNStageIntLLROutputS2xD(348)(4);
  CNStageIntLLRInputS3xD(293)(5) <= VNStageIntLLROutputS2xD(348)(5);
  CNStageIntLLRInputS3xD(373)(5) <= VNStageIntLLROutputS2xD(348)(6);
  CNStageIntLLRInputS3xD(25)(5) <= VNStageIntLLROutputS2xD(349)(0);
  CNStageIntLLRInputS3xD(99)(5) <= VNStageIntLLROutputS2xD(349)(1);
  CNStageIntLLRInputS3xD(180)(5) <= VNStageIntLLROutputS2xD(349)(2);
  CNStageIntLLRInputS3xD(244)(5) <= VNStageIntLLROutputS2xD(349)(3);
  CNStageIntLLRInputS3xD(319)(5) <= VNStageIntLLROutputS2xD(349)(4);
  CNStageIntLLRInputS3xD(352)(5) <= VNStageIntLLROutputS2xD(349)(5);
  CNStageIntLLRInputS3xD(24)(5) <= VNStageIntLLROutputS2xD(350)(0);
  CNStageIntLLRInputS3xD(81)(5) <= VNStageIntLLROutputS2xD(350)(1);
  CNStageIntLLRInputS3xD(164)(5) <= VNStageIntLLROutputS2xD(350)(2);
  CNStageIntLLRInputS3xD(171)(5) <= VNStageIntLLROutputS2xD(350)(3);
  CNStageIntLLRInputS3xD(254)(5) <= VNStageIntLLROutputS2xD(350)(4);
  CNStageIntLLRInputS3xD(303)(5) <= VNStageIntLLROutputS2xD(350)(5);
  CNStageIntLLRInputS3xD(23)(5) <= VNStageIntLLROutputS2xD(351)(0);
  CNStageIntLLRInputS3xD(154)(5) <= VNStageIntLLROutputS2xD(351)(1);
  CNStageIntLLRInputS3xD(188)(5) <= VNStageIntLLROutputS2xD(351)(2);
  CNStageIntLLRInputS3xD(266)(5) <= VNStageIntLLROutputS2xD(351)(3);
  CNStageIntLLRInputS3xD(329)(5) <= VNStageIntLLROutputS2xD(351)(4);
  CNStageIntLLRInputS3xD(340)(5) <= VNStageIntLLROutputS2xD(351)(5);
  CNStageIntLLRInputS3xD(22)(5) <= VNStageIntLLROutputS2xD(352)(0);
  CNStageIntLLRInputS3xD(100)(5) <= VNStageIntLLROutputS2xD(352)(1);
  CNStageIntLLRInputS3xD(141)(5) <= VNStageIntLLROutputS2xD(352)(2);
  CNStageIntLLRInputS3xD(192)(5) <= VNStageIntLLROutputS2xD(352)(3);
  CNStageIntLLRInputS3xD(239)(5) <= VNStageIntLLROutputS2xD(352)(4);
  CNStageIntLLRInputS3xD(321)(5) <= VNStageIntLLROutputS2xD(352)(5);
  CNStageIntLLRInputS3xD(374)(5) <= VNStageIntLLROutputS2xD(352)(6);
  CNStageIntLLRInputS3xD(21)(5) <= VNStageIntLLROutputS2xD(353)(0);
  CNStageIntLLRInputS3xD(74)(5) <= VNStageIntLLROutputS2xD(353)(1);
  CNStageIntLLRInputS3xD(160)(5) <= VNStageIntLLROutputS2xD(353)(2);
  CNStageIntLLRInputS3xD(224)(5) <= VNStageIntLLROutputS2xD(353)(3);
  CNStageIntLLRInputS3xD(227)(5) <= VNStageIntLLROutputS2xD(353)(4);
  CNStageIntLLRInputS3xD(336)(5) <= VNStageIntLLROutputS2xD(353)(5);
  CNStageIntLLRInputS3xD(20)(5) <= VNStageIntLLROutputS2xD(354)(0);
  CNStageIntLLRInputS3xD(88)(5) <= VNStageIntLLROutputS2xD(354)(1);
  CNStageIntLLRInputS3xD(133)(5) <= VNStageIntLLROutputS2xD(354)(2);
  CNStageIntLLRInputS3xD(191)(5) <= VNStageIntLLROutputS2xD(354)(3);
  CNStageIntLLRInputS3xD(326)(5) <= VNStageIntLLROutputS2xD(354)(4);
  CNStageIntLLRInputS3xD(364)(5) <= VNStageIntLLROutputS2xD(354)(5);
  CNStageIntLLRInputS3xD(19)(5) <= VNStageIntLLROutputS2xD(355)(0);
  CNStageIntLLRInputS3xD(59)(5) <= VNStageIntLLROutputS2xD(355)(1);
  CNStageIntLLRInputS3xD(130)(5) <= VNStageIntLLROutputS2xD(355)(2);
  CNStageIntLLRInputS3xD(186)(5) <= VNStageIntLLROutputS2xD(355)(3);
  CNStageIntLLRInputS3xD(230)(5) <= VNStageIntLLROutputS2xD(355)(4);
  CNStageIntLLRInputS3xD(300)(5) <= VNStageIntLLROutputS2xD(355)(5);
  CNStageIntLLRInputS3xD(349)(5) <= VNStageIntLLROutputS2xD(355)(6);
  CNStageIntLLRInputS3xD(18)(5) <= VNStageIntLLROutputS2xD(356)(0);
  CNStageIntLLRInputS3xD(95)(5) <= VNStageIntLLROutputS2xD(356)(1);
  CNStageIntLLRInputS3xD(146)(5) <= VNStageIntLLROutputS2xD(356)(2);
  CNStageIntLLRInputS3xD(222)(5) <= VNStageIntLLROutputS2xD(356)(3);
  CNStageIntLLRInputS3xD(299)(5) <= VNStageIntLLROutputS2xD(356)(4);
  CNStageIntLLRInputS3xD(376)(5) <= VNStageIntLLROutputS2xD(356)(5);
  CNStageIntLLRInputS3xD(17)(5) <= VNStageIntLLROutputS2xD(357)(0);
  CNStageIntLLRInputS3xD(61)(5) <= VNStageIntLLROutputS2xD(357)(1);
  CNStageIntLLRInputS3xD(138)(5) <= VNStageIntLLROutputS2xD(357)(2);
  CNStageIntLLRInputS3xD(176)(5) <= VNStageIntLLROutputS2xD(357)(3);
  CNStageIntLLRInputS3xD(256)(5) <= VNStageIntLLROutputS2xD(357)(4);
  CNStageIntLLRInputS3xD(312)(5) <= VNStageIntLLROutputS2xD(357)(5);
  CNStageIntLLRInputS3xD(366)(5) <= VNStageIntLLROutputS2xD(357)(6);
  CNStageIntLLRInputS3xD(16)(5) <= VNStageIntLLROutputS2xD(358)(0);
  CNStageIntLLRInputS3xD(76)(5) <= VNStageIntLLROutputS2xD(358)(1);
  CNStageIntLLRInputS3xD(112)(5) <= VNStageIntLLROutputS2xD(358)(2);
  CNStageIntLLRInputS3xD(252)(5) <= VNStageIntLLROutputS2xD(358)(3);
  CNStageIntLLRInputS3xD(305)(5) <= VNStageIntLLROutputS2xD(358)(4);
  CNStageIntLLRInputS3xD(353)(5) <= VNStageIntLLROutputS2xD(358)(5);
  CNStageIntLLRInputS3xD(15)(5) <= VNStageIntLLROutputS2xD(359)(0);
  CNStageIntLLRInputS3xD(72)(5) <= VNStageIntLLROutputS2xD(359)(1);
  CNStageIntLLRInputS3xD(122)(5) <= VNStageIntLLROutputS2xD(359)(2);
  CNStageIntLLRInputS3xD(195)(5) <= VNStageIntLLROutputS2xD(359)(3);
  CNStageIntLLRInputS3xD(257)(5) <= VNStageIntLLROutputS2xD(359)(4);
  CNStageIntLLRInputS3xD(283)(5) <= VNStageIntLLROutputS2xD(359)(5);
  CNStageIntLLRInputS3xD(372)(5) <= VNStageIntLLROutputS2xD(359)(6);
  CNStageIntLLRInputS3xD(14)(5) <= VNStageIntLLROutputS2xD(360)(0);
  CNStageIntLLRInputS3xD(91)(5) <= VNStageIntLLROutputS2xD(360)(1);
  CNStageIntLLRInputS3xD(116)(5) <= VNStageIntLLROutputS2xD(360)(2);
  CNStageIntLLRInputS3xD(174)(5) <= VNStageIntLLROutputS2xD(360)(3);
  CNStageIntLLRInputS3xD(248)(5) <= VNStageIntLLROutputS2xD(360)(4);
  CNStageIntLLRInputS3xD(292)(5) <= VNStageIntLLROutputS2xD(360)(5);
  CNStageIntLLRInputS3xD(345)(5) <= VNStageIntLLROutputS2xD(360)(6);
  CNStageIntLLRInputS3xD(13)(5) <= VNStageIntLLROutputS2xD(361)(0);
  CNStageIntLLRInputS3xD(54)(5) <= VNStageIntLLROutputS2xD(361)(1);
  CNStageIntLLRInputS3xD(120)(5) <= VNStageIntLLROutputS2xD(361)(2);
  CNStageIntLLRInputS3xD(207)(5) <= VNStageIntLLROutputS2xD(361)(3);
  CNStageIntLLRInputS3xD(271)(5) <= VNStageIntLLROutputS2xD(361)(4);
  CNStageIntLLRInputS3xD(285)(5) <= VNStageIntLLROutputS2xD(361)(5);
  CNStageIntLLRInputS3xD(342)(5) <= VNStageIntLLROutputS2xD(361)(6);
  CNStageIntLLRInputS3xD(12)(5) <= VNStageIntLLROutputS2xD(362)(0);
  CNStageIntLLRInputS3xD(55)(5) <= VNStageIntLLROutputS2xD(362)(1);
  CNStageIntLLRInputS3xD(169)(5) <= VNStageIntLLROutputS2xD(362)(2);
  CNStageIntLLRInputS3xD(210)(5) <= VNStageIntLLROutputS2xD(362)(3);
  CNStageIntLLRInputS3xD(276)(5) <= VNStageIntLLROutputS2xD(362)(4);
  CNStageIntLLRInputS3xD(289)(5) <= VNStageIntLLROutputS2xD(362)(5);
  CNStageIntLLRInputS3xD(357)(5) <= VNStageIntLLROutputS2xD(362)(6);
  CNStageIntLLRInputS3xD(90)(5) <= VNStageIntLLROutputS2xD(363)(0);
  CNStageIntLLRInputS3xD(147)(5) <= VNStageIntLLROutputS2xD(363)(1);
  CNStageIntLLRInputS3xD(197)(5) <= VNStageIntLLROutputS2xD(363)(2);
  CNStageIntLLRInputS3xD(261)(5) <= VNStageIntLLROutputS2xD(363)(3);
  CNStageIntLLRInputS3xD(281)(5) <= VNStageIntLLROutputS2xD(363)(4);
  CNStageIntLLRInputS3xD(11)(5) <= VNStageIntLLROutputS2xD(364)(0);
  CNStageIntLLRInputS3xD(82)(5) <= VNStageIntLLROutputS2xD(364)(1);
  CNStageIntLLRInputS3xD(129)(5) <= VNStageIntLLROutputS2xD(364)(2);
  CNStageIntLLRInputS3xD(175)(5) <= VNStageIntLLROutputS2xD(364)(3);
  CNStageIntLLRInputS3xD(263)(5) <= VNStageIntLLROutputS2xD(364)(4);
  CNStageIntLLRInputS3xD(313)(5) <= VNStageIntLLROutputS2xD(364)(5);
  CNStageIntLLRInputS3xD(10)(5) <= VNStageIntLLROutputS2xD(365)(0);
  CNStageIntLLRInputS3xD(98)(5) <= VNStageIntLLROutputS2xD(365)(1);
  CNStageIntLLRInputS3xD(142)(5) <= VNStageIntLLROutputS2xD(365)(2);
  CNStageIntLLRInputS3xD(194)(5) <= VNStageIntLLROutputS2xD(365)(3);
  CNStageIntLLRInputS3xD(234)(5) <= VNStageIntLLROutputS2xD(365)(4);
  CNStageIntLLRInputS3xD(298)(5) <= VNStageIntLLROutputS2xD(365)(5);
  CNStageIntLLRInputS3xD(9)(5) <= VNStageIntLLROutputS2xD(366)(0);
  CNStageIntLLRInputS3xD(102)(5) <= VNStageIntLLROutputS2xD(366)(1);
  CNStageIntLLRInputS3xD(153)(5) <= VNStageIntLLROutputS2xD(366)(2);
  CNStageIntLLRInputS3xD(219)(5) <= VNStageIntLLROutputS2xD(366)(3);
  CNStageIntLLRInputS3xD(269)(5) <= VNStageIntLLROutputS2xD(366)(4);
  CNStageIntLLRInputS3xD(308)(5) <= VNStageIntLLROutputS2xD(366)(5);
  CNStageIntLLRInputS3xD(8)(5) <= VNStageIntLLROutputS2xD(367)(0);
  CNStageIntLLRInputS3xD(110)(5) <= VNStageIntLLROutputS2xD(367)(1);
  CNStageIntLLRInputS3xD(123)(5) <= VNStageIntLLROutputS2xD(367)(2);
  CNStageIntLLRInputS3xD(205)(5) <= VNStageIntLLROutputS2xD(367)(3);
  CNStageIntLLRInputS3xD(226)(5) <= VNStageIntLLROutputS2xD(367)(4);
  CNStageIntLLRInputS3xD(320)(5) <= VNStageIntLLROutputS2xD(367)(5);
  CNStageIntLLRInputS3xD(333)(5) <= VNStageIntLLROutputS2xD(367)(6);
  CNStageIntLLRInputS3xD(7)(5) <= VNStageIntLLROutputS2xD(368)(0);
  CNStageIntLLRInputS3xD(177)(5) <= VNStageIntLLROutputS2xD(368)(1);
  CNStageIntLLRInputS3xD(381)(5) <= VNStageIntLLROutputS2xD(368)(2);
  CNStageIntLLRInputS3xD(6)(5) <= VNStageIntLLROutputS2xD(369)(0);
  CNStageIntLLRInputS3xD(156)(5) <= VNStageIntLLROutputS2xD(369)(1);
  CNStageIntLLRInputS3xD(221)(5) <= VNStageIntLLROutputS2xD(369)(2);
  CNStageIntLLRInputS3xD(262)(5) <= VNStageIntLLROutputS2xD(369)(3);
  CNStageIntLLRInputS3xD(358)(5) <= VNStageIntLLROutputS2xD(369)(4);
  CNStageIntLLRInputS3xD(5)(5) <= VNStageIntLLROutputS2xD(370)(0);
  CNStageIntLLRInputS3xD(114)(5) <= VNStageIntLLROutputS2xD(370)(1);
  CNStageIntLLRInputS3xD(208)(5) <= VNStageIntLLROutputS2xD(370)(2);
  CNStageIntLLRInputS3xD(275)(5) <= VNStageIntLLROutputS2xD(370)(3);
  CNStageIntLLRInputS3xD(341)(5) <= VNStageIntLLROutputS2xD(370)(4);
  CNStageIntLLRInputS3xD(4)(5) <= VNStageIntLLROutputS2xD(371)(0);
  CNStageIntLLRInputS3xD(135)(5) <= VNStageIntLLROutputS2xD(371)(1);
  CNStageIntLLRInputS3xD(173)(5) <= VNStageIntLLROutputS2xD(371)(2);
  CNStageIntLLRInputS3xD(249)(5) <= VNStageIntLLROutputS2xD(371)(3);
  CNStageIntLLRInputS3xD(354)(5) <= VNStageIntLLROutputS2xD(371)(4);
  CNStageIntLLRInputS3xD(106)(5) <= VNStageIntLLROutputS2xD(372)(0);
  CNStageIntLLRInputS3xD(144)(5) <= VNStageIntLLROutputS2xD(372)(1);
  CNStageIntLLRInputS3xD(201)(5) <= VNStageIntLLROutputS2xD(372)(2);
  CNStageIntLLRInputS3xD(229)(5) <= VNStageIntLLROutputS2xD(372)(3);
  CNStageIntLLRInputS3xD(301)(5) <= VNStageIntLLROutputS2xD(372)(4);
  CNStageIntLLRInputS3xD(365)(5) <= VNStageIntLLROutputS2xD(372)(5);
  CNStageIntLLRInputS3xD(3)(5) <= VNStageIntLLROutputS2xD(373)(0);
  CNStageIntLLRInputS3xD(139)(5) <= VNStageIntLLROutputS2xD(373)(1);
  CNStageIntLLRInputS3xD(250)(5) <= VNStageIntLLROutputS2xD(373)(2);
  CNStageIntLLRInputS3xD(310)(5) <= VNStageIntLLROutputS2xD(373)(3);
  CNStageIntLLRInputS3xD(335)(5) <= VNStageIntLLROutputS2xD(373)(4);
  CNStageIntLLRInputS3xD(2)(5) <= VNStageIntLLROutputS2xD(374)(0);
  CNStageIntLLRInputS3xD(85)(5) <= VNStageIntLLROutputS2xD(374)(1);
  CNStageIntLLRInputS3xD(145)(5) <= VNStageIntLLROutputS2xD(374)(2);
  CNStageIntLLRInputS3xD(213)(5) <= VNStageIntLLROutputS2xD(374)(3);
  CNStageIntLLRInputS3xD(264)(5) <= VNStageIntLLROutputS2xD(374)(4);
  CNStageIntLLRInputS3xD(306)(5) <= VNStageIntLLROutputS2xD(374)(5);
  CNStageIntLLRInputS3xD(383)(5) <= VNStageIntLLROutputS2xD(374)(6);
  CNStageIntLLRInputS3xD(1)(5) <= VNStageIntLLROutputS2xD(375)(0);
  CNStageIntLLRInputS3xD(64)(5) <= VNStageIntLLROutputS2xD(375)(1);
  CNStageIntLLRInputS3xD(134)(5) <= VNStageIntLLROutputS2xD(375)(2);
  CNStageIntLLRInputS3xD(260)(5) <= VNStageIntLLROutputS2xD(375)(3);
  CNStageIntLLRInputS3xD(311)(5) <= VNStageIntLLROutputS2xD(375)(4);
  CNStageIntLLRInputS3xD(368)(5) <= VNStageIntLLROutputS2xD(375)(5);
  CNStageIntLLRInputS3xD(0)(5) <= VNStageIntLLROutputS2xD(376)(0);
  CNStageIntLLRInputS3xD(67)(5) <= VNStageIntLLROutputS2xD(376)(1);
  CNStageIntLLRInputS3xD(159)(5) <= VNStageIntLLROutputS2xD(376)(2);
  CNStageIntLLRInputS3xD(278)(5) <= VNStageIntLLROutputS2xD(376)(3);
  CNStageIntLLRInputS3xD(107)(5) <= VNStageIntLLROutputS2xD(377)(0);
  CNStageIntLLRInputS3xD(166)(5) <= VNStageIntLLROutputS2xD(377)(1);
  CNStageIntLLRInputS3xD(193)(5) <= VNStageIntLLROutputS2xD(377)(2);
  CNStageIntLLRInputS3xD(325)(5) <= VNStageIntLLROutputS2xD(377)(3);
  CNStageIntLLRInputS3xD(347)(5) <= VNStageIntLLROutputS2xD(377)(4);
  CNStageIntLLRInputS3xD(86)(5) <= VNStageIntLLROutputS2xD(378)(0);
  CNStageIntLLRInputS3xD(149)(5) <= VNStageIntLLROutputS2xD(378)(1);
  CNStageIntLLRInputS3xD(187)(5) <= VNStageIntLLROutputS2xD(378)(2);
  CNStageIntLLRInputS3xD(246)(5) <= VNStageIntLLROutputS2xD(378)(3);
  CNStageIntLLRInputS3xD(331)(5) <= VNStageIntLLROutputS2xD(378)(4);
  CNStageIntLLRInputS3xD(355)(5) <= VNStageIntLLROutputS2xD(378)(5);
  CNStageIntLLRInputS3xD(105)(5) <= VNStageIntLLROutputS2xD(379)(0);
  CNStageIntLLRInputS3xD(151)(5) <= VNStageIntLLROutputS2xD(379)(1);
  CNStageIntLLRInputS3xD(277)(5) <= VNStageIntLLROutputS2xD(379)(2);
  CNStageIntLLRInputS3xD(315)(5) <= VNStageIntLLROutputS2xD(379)(3);
  CNStageIntLLRInputS3xD(351)(5) <= VNStageIntLLROutputS2xD(379)(4);
  CNStageIntLLRInputS3xD(77)(5) <= VNStageIntLLROutputS2xD(380)(0);
  CNStageIntLLRInputS3xD(118)(5) <= VNStageIntLLROutputS2xD(380)(1);
  CNStageIntLLRInputS3xD(182)(5) <= VNStageIntLLROutputS2xD(380)(2);
  CNStageIntLLRInputS3xD(270)(5) <= VNStageIntLLROutputS2xD(380)(3);
  CNStageIntLLRInputS3xD(317)(5) <= VNStageIntLLROutputS2xD(380)(4);
  CNStageIntLLRInputS3xD(356)(5) <= VNStageIntLLROutputS2xD(380)(5);
  CNStageIntLLRInputS3xD(60)(5) <= VNStageIntLLROutputS2xD(381)(0);
  CNStageIntLLRInputS3xD(157)(5) <= VNStageIntLLROutputS2xD(381)(1);
  CNStageIntLLRInputS3xD(214)(5) <= VNStageIntLLROutputS2xD(381)(2);
  CNStageIntLLRInputS3xD(233)(5) <= VNStageIntLLROutputS2xD(381)(3);
  CNStageIntLLRInputS3xD(287)(5) <= VNStageIntLLROutputS2xD(381)(4);
  CNStageIntLLRInputS3xD(346)(5) <= VNStageIntLLROutputS2xD(381)(5);
  CNStageIntLLRInputS3xD(87)(5) <= VNStageIntLLROutputS2xD(382)(0);
  CNStageIntLLRInputS3xD(111)(5) <= VNStageIntLLROutputS2xD(382)(1);
  CNStageIntLLRInputS3xD(198)(5) <= VNStageIntLLROutputS2xD(382)(2);
  CNStageIntLLRInputS3xD(237)(5) <= VNStageIntLLROutputS2xD(382)(3);
  CNStageIntLLRInputS3xD(323)(5) <= VNStageIntLLROutputS2xD(382)(4);
  CNStageIntLLRInputS3xD(371)(5) <= VNStageIntLLROutputS2xD(382)(5);
  CNStageIntLLRInputS3xD(52)(5) <= VNStageIntLLROutputS2xD(383)(0);
  CNStageIntLLRInputS3xD(79)(5) <= VNStageIntLLROutputS2xD(383)(1);
  CNStageIntLLRInputS3xD(119)(5) <= VNStageIntLLROutputS2xD(383)(2);
  CNStageIntLLRInputS3xD(209)(5) <= VNStageIntLLROutputS2xD(383)(3);
  CNStageIntLLRInputS3xD(279)(5) <= VNStageIntLLROutputS2xD(383)(4);
  CNStageIntLLRInputS3xD(282)(5) <= VNStageIntLLROutputS2xD(383)(5);
  CNStageIntLLRInputS3xD(378)(5) <= VNStageIntLLROutputS2xD(383)(6);

  -- Variable Nodes (Iteration 3)
  VNStageIntLLRInputS3xD(56)(0) <= CNStageIntLLROutputS3xD(0)(0);
  VNStageIntLLRInputS3xD(120)(0) <= CNStageIntLLROutputS3xD(0)(1);
  VNStageIntLLRInputS3xD(184)(0) <= CNStageIntLLROutputS3xD(0)(2);
  VNStageIntLLRInputS3xD(248)(0) <= CNStageIntLLROutputS3xD(0)(3);
  VNStageIntLLRInputS3xD(312)(0) <= CNStageIntLLROutputS3xD(0)(4);
  VNStageIntLLRInputS3xD(376)(0) <= CNStageIntLLROutputS3xD(0)(5);
  VNStageIntLLRInputS3xD(55)(0) <= CNStageIntLLROutputS3xD(1)(0);
  VNStageIntLLRInputS3xD(119)(0) <= CNStageIntLLROutputS3xD(1)(1);
  VNStageIntLLRInputS3xD(183)(0) <= CNStageIntLLROutputS3xD(1)(2);
  VNStageIntLLRInputS3xD(247)(0) <= CNStageIntLLROutputS3xD(1)(3);
  VNStageIntLLRInputS3xD(311)(0) <= CNStageIntLLROutputS3xD(1)(4);
  VNStageIntLLRInputS3xD(375)(0) <= CNStageIntLLROutputS3xD(1)(5);
  VNStageIntLLRInputS3xD(54)(0) <= CNStageIntLLROutputS3xD(2)(0);
  VNStageIntLLRInputS3xD(118)(0) <= CNStageIntLLROutputS3xD(2)(1);
  VNStageIntLLRInputS3xD(182)(0) <= CNStageIntLLROutputS3xD(2)(2);
  VNStageIntLLRInputS3xD(246)(0) <= CNStageIntLLROutputS3xD(2)(3);
  VNStageIntLLRInputS3xD(310)(0) <= CNStageIntLLROutputS3xD(2)(4);
  VNStageIntLLRInputS3xD(374)(0) <= CNStageIntLLROutputS3xD(2)(5);
  VNStageIntLLRInputS3xD(53)(0) <= CNStageIntLLROutputS3xD(3)(0);
  VNStageIntLLRInputS3xD(117)(0) <= CNStageIntLLROutputS3xD(3)(1);
  VNStageIntLLRInputS3xD(181)(0) <= CNStageIntLLROutputS3xD(3)(2);
  VNStageIntLLRInputS3xD(245)(0) <= CNStageIntLLROutputS3xD(3)(3);
  VNStageIntLLRInputS3xD(309)(0) <= CNStageIntLLROutputS3xD(3)(4);
  VNStageIntLLRInputS3xD(373)(0) <= CNStageIntLLROutputS3xD(3)(5);
  VNStageIntLLRInputS3xD(51)(0) <= CNStageIntLLROutputS3xD(4)(0);
  VNStageIntLLRInputS3xD(115)(0) <= CNStageIntLLROutputS3xD(4)(1);
  VNStageIntLLRInputS3xD(179)(0) <= CNStageIntLLROutputS3xD(4)(2);
  VNStageIntLLRInputS3xD(243)(0) <= CNStageIntLLROutputS3xD(4)(3);
  VNStageIntLLRInputS3xD(307)(0) <= CNStageIntLLROutputS3xD(4)(4);
  VNStageIntLLRInputS3xD(371)(0) <= CNStageIntLLROutputS3xD(4)(5);
  VNStageIntLLRInputS3xD(50)(0) <= CNStageIntLLROutputS3xD(5)(0);
  VNStageIntLLRInputS3xD(114)(0) <= CNStageIntLLROutputS3xD(5)(1);
  VNStageIntLLRInputS3xD(178)(0) <= CNStageIntLLROutputS3xD(5)(2);
  VNStageIntLLRInputS3xD(242)(0) <= CNStageIntLLROutputS3xD(5)(3);
  VNStageIntLLRInputS3xD(306)(0) <= CNStageIntLLROutputS3xD(5)(4);
  VNStageIntLLRInputS3xD(370)(0) <= CNStageIntLLROutputS3xD(5)(5);
  VNStageIntLLRInputS3xD(49)(0) <= CNStageIntLLROutputS3xD(6)(0);
  VNStageIntLLRInputS3xD(113)(0) <= CNStageIntLLROutputS3xD(6)(1);
  VNStageIntLLRInputS3xD(177)(0) <= CNStageIntLLROutputS3xD(6)(2);
  VNStageIntLLRInputS3xD(241)(0) <= CNStageIntLLROutputS3xD(6)(3);
  VNStageIntLLRInputS3xD(305)(0) <= CNStageIntLLROutputS3xD(6)(4);
  VNStageIntLLRInputS3xD(369)(0) <= CNStageIntLLROutputS3xD(6)(5);
  VNStageIntLLRInputS3xD(48)(0) <= CNStageIntLLROutputS3xD(7)(0);
  VNStageIntLLRInputS3xD(112)(0) <= CNStageIntLLROutputS3xD(7)(1);
  VNStageIntLLRInputS3xD(176)(0) <= CNStageIntLLROutputS3xD(7)(2);
  VNStageIntLLRInputS3xD(240)(0) <= CNStageIntLLROutputS3xD(7)(3);
  VNStageIntLLRInputS3xD(304)(0) <= CNStageIntLLROutputS3xD(7)(4);
  VNStageIntLLRInputS3xD(368)(0) <= CNStageIntLLROutputS3xD(7)(5);
  VNStageIntLLRInputS3xD(47)(0) <= CNStageIntLLROutputS3xD(8)(0);
  VNStageIntLLRInputS3xD(111)(0) <= CNStageIntLLROutputS3xD(8)(1);
  VNStageIntLLRInputS3xD(175)(0) <= CNStageIntLLROutputS3xD(8)(2);
  VNStageIntLLRInputS3xD(239)(0) <= CNStageIntLLROutputS3xD(8)(3);
  VNStageIntLLRInputS3xD(303)(0) <= CNStageIntLLROutputS3xD(8)(4);
  VNStageIntLLRInputS3xD(367)(0) <= CNStageIntLLROutputS3xD(8)(5);
  VNStageIntLLRInputS3xD(46)(0) <= CNStageIntLLROutputS3xD(9)(0);
  VNStageIntLLRInputS3xD(110)(0) <= CNStageIntLLROutputS3xD(9)(1);
  VNStageIntLLRInputS3xD(174)(0) <= CNStageIntLLROutputS3xD(9)(2);
  VNStageIntLLRInputS3xD(238)(0) <= CNStageIntLLROutputS3xD(9)(3);
  VNStageIntLLRInputS3xD(302)(0) <= CNStageIntLLROutputS3xD(9)(4);
  VNStageIntLLRInputS3xD(366)(0) <= CNStageIntLLROutputS3xD(9)(5);
  VNStageIntLLRInputS3xD(45)(0) <= CNStageIntLLROutputS3xD(10)(0);
  VNStageIntLLRInputS3xD(109)(0) <= CNStageIntLLROutputS3xD(10)(1);
  VNStageIntLLRInputS3xD(173)(0) <= CNStageIntLLROutputS3xD(10)(2);
  VNStageIntLLRInputS3xD(237)(0) <= CNStageIntLLROutputS3xD(10)(3);
  VNStageIntLLRInputS3xD(301)(0) <= CNStageIntLLROutputS3xD(10)(4);
  VNStageIntLLRInputS3xD(365)(0) <= CNStageIntLLROutputS3xD(10)(5);
  VNStageIntLLRInputS3xD(44)(0) <= CNStageIntLLROutputS3xD(11)(0);
  VNStageIntLLRInputS3xD(108)(0) <= CNStageIntLLROutputS3xD(11)(1);
  VNStageIntLLRInputS3xD(172)(0) <= CNStageIntLLROutputS3xD(11)(2);
  VNStageIntLLRInputS3xD(236)(0) <= CNStageIntLLROutputS3xD(11)(3);
  VNStageIntLLRInputS3xD(300)(0) <= CNStageIntLLROutputS3xD(11)(4);
  VNStageIntLLRInputS3xD(364)(0) <= CNStageIntLLROutputS3xD(11)(5);
  VNStageIntLLRInputS3xD(42)(0) <= CNStageIntLLROutputS3xD(12)(0);
  VNStageIntLLRInputS3xD(106)(0) <= CNStageIntLLROutputS3xD(12)(1);
  VNStageIntLLRInputS3xD(170)(0) <= CNStageIntLLROutputS3xD(12)(2);
  VNStageIntLLRInputS3xD(234)(0) <= CNStageIntLLROutputS3xD(12)(3);
  VNStageIntLLRInputS3xD(298)(0) <= CNStageIntLLROutputS3xD(12)(4);
  VNStageIntLLRInputS3xD(362)(0) <= CNStageIntLLROutputS3xD(12)(5);
  VNStageIntLLRInputS3xD(41)(0) <= CNStageIntLLROutputS3xD(13)(0);
  VNStageIntLLRInputS3xD(105)(0) <= CNStageIntLLROutputS3xD(13)(1);
  VNStageIntLLRInputS3xD(169)(0) <= CNStageIntLLROutputS3xD(13)(2);
  VNStageIntLLRInputS3xD(233)(0) <= CNStageIntLLROutputS3xD(13)(3);
  VNStageIntLLRInputS3xD(297)(0) <= CNStageIntLLROutputS3xD(13)(4);
  VNStageIntLLRInputS3xD(361)(0) <= CNStageIntLLROutputS3xD(13)(5);
  VNStageIntLLRInputS3xD(40)(0) <= CNStageIntLLROutputS3xD(14)(0);
  VNStageIntLLRInputS3xD(104)(0) <= CNStageIntLLROutputS3xD(14)(1);
  VNStageIntLLRInputS3xD(168)(0) <= CNStageIntLLROutputS3xD(14)(2);
  VNStageIntLLRInputS3xD(232)(0) <= CNStageIntLLROutputS3xD(14)(3);
  VNStageIntLLRInputS3xD(296)(0) <= CNStageIntLLROutputS3xD(14)(4);
  VNStageIntLLRInputS3xD(360)(0) <= CNStageIntLLROutputS3xD(14)(5);
  VNStageIntLLRInputS3xD(39)(0) <= CNStageIntLLROutputS3xD(15)(0);
  VNStageIntLLRInputS3xD(103)(0) <= CNStageIntLLROutputS3xD(15)(1);
  VNStageIntLLRInputS3xD(167)(0) <= CNStageIntLLROutputS3xD(15)(2);
  VNStageIntLLRInputS3xD(231)(0) <= CNStageIntLLROutputS3xD(15)(3);
  VNStageIntLLRInputS3xD(295)(0) <= CNStageIntLLROutputS3xD(15)(4);
  VNStageIntLLRInputS3xD(359)(0) <= CNStageIntLLROutputS3xD(15)(5);
  VNStageIntLLRInputS3xD(38)(0) <= CNStageIntLLROutputS3xD(16)(0);
  VNStageIntLLRInputS3xD(102)(0) <= CNStageIntLLROutputS3xD(16)(1);
  VNStageIntLLRInputS3xD(166)(0) <= CNStageIntLLROutputS3xD(16)(2);
  VNStageIntLLRInputS3xD(230)(0) <= CNStageIntLLROutputS3xD(16)(3);
  VNStageIntLLRInputS3xD(294)(0) <= CNStageIntLLROutputS3xD(16)(4);
  VNStageIntLLRInputS3xD(358)(0) <= CNStageIntLLROutputS3xD(16)(5);
  VNStageIntLLRInputS3xD(37)(0) <= CNStageIntLLROutputS3xD(17)(0);
  VNStageIntLLRInputS3xD(101)(0) <= CNStageIntLLROutputS3xD(17)(1);
  VNStageIntLLRInputS3xD(165)(0) <= CNStageIntLLROutputS3xD(17)(2);
  VNStageIntLLRInputS3xD(229)(0) <= CNStageIntLLROutputS3xD(17)(3);
  VNStageIntLLRInputS3xD(293)(0) <= CNStageIntLLROutputS3xD(17)(4);
  VNStageIntLLRInputS3xD(357)(0) <= CNStageIntLLROutputS3xD(17)(5);
  VNStageIntLLRInputS3xD(36)(0) <= CNStageIntLLROutputS3xD(18)(0);
  VNStageIntLLRInputS3xD(100)(0) <= CNStageIntLLROutputS3xD(18)(1);
  VNStageIntLLRInputS3xD(164)(0) <= CNStageIntLLROutputS3xD(18)(2);
  VNStageIntLLRInputS3xD(228)(0) <= CNStageIntLLROutputS3xD(18)(3);
  VNStageIntLLRInputS3xD(292)(0) <= CNStageIntLLROutputS3xD(18)(4);
  VNStageIntLLRInputS3xD(356)(0) <= CNStageIntLLROutputS3xD(18)(5);
  VNStageIntLLRInputS3xD(35)(0) <= CNStageIntLLROutputS3xD(19)(0);
  VNStageIntLLRInputS3xD(99)(0) <= CNStageIntLLROutputS3xD(19)(1);
  VNStageIntLLRInputS3xD(163)(0) <= CNStageIntLLROutputS3xD(19)(2);
  VNStageIntLLRInputS3xD(227)(0) <= CNStageIntLLROutputS3xD(19)(3);
  VNStageIntLLRInputS3xD(291)(0) <= CNStageIntLLROutputS3xD(19)(4);
  VNStageIntLLRInputS3xD(355)(0) <= CNStageIntLLROutputS3xD(19)(5);
  VNStageIntLLRInputS3xD(34)(0) <= CNStageIntLLROutputS3xD(20)(0);
  VNStageIntLLRInputS3xD(98)(0) <= CNStageIntLLROutputS3xD(20)(1);
  VNStageIntLLRInputS3xD(162)(0) <= CNStageIntLLROutputS3xD(20)(2);
  VNStageIntLLRInputS3xD(226)(0) <= CNStageIntLLROutputS3xD(20)(3);
  VNStageIntLLRInputS3xD(290)(0) <= CNStageIntLLROutputS3xD(20)(4);
  VNStageIntLLRInputS3xD(354)(0) <= CNStageIntLLROutputS3xD(20)(5);
  VNStageIntLLRInputS3xD(33)(0) <= CNStageIntLLROutputS3xD(21)(0);
  VNStageIntLLRInputS3xD(97)(0) <= CNStageIntLLROutputS3xD(21)(1);
  VNStageIntLLRInputS3xD(161)(0) <= CNStageIntLLROutputS3xD(21)(2);
  VNStageIntLLRInputS3xD(225)(0) <= CNStageIntLLROutputS3xD(21)(3);
  VNStageIntLLRInputS3xD(289)(0) <= CNStageIntLLROutputS3xD(21)(4);
  VNStageIntLLRInputS3xD(353)(0) <= CNStageIntLLROutputS3xD(21)(5);
  VNStageIntLLRInputS3xD(32)(0) <= CNStageIntLLROutputS3xD(22)(0);
  VNStageIntLLRInputS3xD(96)(0) <= CNStageIntLLROutputS3xD(22)(1);
  VNStageIntLLRInputS3xD(160)(0) <= CNStageIntLLROutputS3xD(22)(2);
  VNStageIntLLRInputS3xD(224)(0) <= CNStageIntLLROutputS3xD(22)(3);
  VNStageIntLLRInputS3xD(288)(0) <= CNStageIntLLROutputS3xD(22)(4);
  VNStageIntLLRInputS3xD(352)(0) <= CNStageIntLLROutputS3xD(22)(5);
  VNStageIntLLRInputS3xD(31)(0) <= CNStageIntLLROutputS3xD(23)(0);
  VNStageIntLLRInputS3xD(95)(0) <= CNStageIntLLROutputS3xD(23)(1);
  VNStageIntLLRInputS3xD(159)(0) <= CNStageIntLLROutputS3xD(23)(2);
  VNStageIntLLRInputS3xD(223)(0) <= CNStageIntLLROutputS3xD(23)(3);
  VNStageIntLLRInputS3xD(287)(0) <= CNStageIntLLROutputS3xD(23)(4);
  VNStageIntLLRInputS3xD(351)(0) <= CNStageIntLLROutputS3xD(23)(5);
  VNStageIntLLRInputS3xD(30)(0) <= CNStageIntLLROutputS3xD(24)(0);
  VNStageIntLLRInputS3xD(94)(0) <= CNStageIntLLROutputS3xD(24)(1);
  VNStageIntLLRInputS3xD(158)(0) <= CNStageIntLLROutputS3xD(24)(2);
  VNStageIntLLRInputS3xD(222)(0) <= CNStageIntLLROutputS3xD(24)(3);
  VNStageIntLLRInputS3xD(286)(0) <= CNStageIntLLROutputS3xD(24)(4);
  VNStageIntLLRInputS3xD(350)(0) <= CNStageIntLLROutputS3xD(24)(5);
  VNStageIntLLRInputS3xD(29)(0) <= CNStageIntLLROutputS3xD(25)(0);
  VNStageIntLLRInputS3xD(93)(0) <= CNStageIntLLROutputS3xD(25)(1);
  VNStageIntLLRInputS3xD(157)(0) <= CNStageIntLLROutputS3xD(25)(2);
  VNStageIntLLRInputS3xD(221)(0) <= CNStageIntLLROutputS3xD(25)(3);
  VNStageIntLLRInputS3xD(285)(0) <= CNStageIntLLROutputS3xD(25)(4);
  VNStageIntLLRInputS3xD(349)(0) <= CNStageIntLLROutputS3xD(25)(5);
  VNStageIntLLRInputS3xD(28)(0) <= CNStageIntLLROutputS3xD(26)(0);
  VNStageIntLLRInputS3xD(92)(0) <= CNStageIntLLROutputS3xD(26)(1);
  VNStageIntLLRInputS3xD(156)(0) <= CNStageIntLLROutputS3xD(26)(2);
  VNStageIntLLRInputS3xD(220)(0) <= CNStageIntLLROutputS3xD(26)(3);
  VNStageIntLLRInputS3xD(284)(0) <= CNStageIntLLROutputS3xD(26)(4);
  VNStageIntLLRInputS3xD(348)(0) <= CNStageIntLLROutputS3xD(26)(5);
  VNStageIntLLRInputS3xD(27)(0) <= CNStageIntLLROutputS3xD(27)(0);
  VNStageIntLLRInputS3xD(91)(0) <= CNStageIntLLROutputS3xD(27)(1);
  VNStageIntLLRInputS3xD(155)(0) <= CNStageIntLLROutputS3xD(27)(2);
  VNStageIntLLRInputS3xD(219)(0) <= CNStageIntLLROutputS3xD(27)(3);
  VNStageIntLLRInputS3xD(283)(0) <= CNStageIntLLROutputS3xD(27)(4);
  VNStageIntLLRInputS3xD(347)(0) <= CNStageIntLLROutputS3xD(27)(5);
  VNStageIntLLRInputS3xD(26)(0) <= CNStageIntLLROutputS3xD(28)(0);
  VNStageIntLLRInputS3xD(90)(0) <= CNStageIntLLROutputS3xD(28)(1);
  VNStageIntLLRInputS3xD(154)(0) <= CNStageIntLLROutputS3xD(28)(2);
  VNStageIntLLRInputS3xD(218)(0) <= CNStageIntLLROutputS3xD(28)(3);
  VNStageIntLLRInputS3xD(282)(0) <= CNStageIntLLROutputS3xD(28)(4);
  VNStageIntLLRInputS3xD(346)(0) <= CNStageIntLLROutputS3xD(28)(5);
  VNStageIntLLRInputS3xD(25)(0) <= CNStageIntLLROutputS3xD(29)(0);
  VNStageIntLLRInputS3xD(89)(0) <= CNStageIntLLROutputS3xD(29)(1);
  VNStageIntLLRInputS3xD(153)(0) <= CNStageIntLLROutputS3xD(29)(2);
  VNStageIntLLRInputS3xD(217)(0) <= CNStageIntLLROutputS3xD(29)(3);
  VNStageIntLLRInputS3xD(281)(0) <= CNStageIntLLROutputS3xD(29)(4);
  VNStageIntLLRInputS3xD(345)(0) <= CNStageIntLLROutputS3xD(29)(5);
  VNStageIntLLRInputS3xD(24)(0) <= CNStageIntLLROutputS3xD(30)(0);
  VNStageIntLLRInputS3xD(88)(0) <= CNStageIntLLROutputS3xD(30)(1);
  VNStageIntLLRInputS3xD(152)(0) <= CNStageIntLLROutputS3xD(30)(2);
  VNStageIntLLRInputS3xD(216)(0) <= CNStageIntLLROutputS3xD(30)(3);
  VNStageIntLLRInputS3xD(280)(0) <= CNStageIntLLROutputS3xD(30)(4);
  VNStageIntLLRInputS3xD(344)(0) <= CNStageIntLLROutputS3xD(30)(5);
  VNStageIntLLRInputS3xD(23)(0) <= CNStageIntLLROutputS3xD(31)(0);
  VNStageIntLLRInputS3xD(87)(0) <= CNStageIntLLROutputS3xD(31)(1);
  VNStageIntLLRInputS3xD(151)(0) <= CNStageIntLLROutputS3xD(31)(2);
  VNStageIntLLRInputS3xD(215)(0) <= CNStageIntLLROutputS3xD(31)(3);
  VNStageIntLLRInputS3xD(279)(0) <= CNStageIntLLROutputS3xD(31)(4);
  VNStageIntLLRInputS3xD(343)(0) <= CNStageIntLLROutputS3xD(31)(5);
  VNStageIntLLRInputS3xD(22)(0) <= CNStageIntLLROutputS3xD(32)(0);
  VNStageIntLLRInputS3xD(86)(0) <= CNStageIntLLROutputS3xD(32)(1);
  VNStageIntLLRInputS3xD(150)(0) <= CNStageIntLLROutputS3xD(32)(2);
  VNStageIntLLRInputS3xD(214)(0) <= CNStageIntLLROutputS3xD(32)(3);
  VNStageIntLLRInputS3xD(278)(0) <= CNStageIntLLROutputS3xD(32)(4);
  VNStageIntLLRInputS3xD(342)(0) <= CNStageIntLLROutputS3xD(32)(5);
  VNStageIntLLRInputS3xD(21)(0) <= CNStageIntLLROutputS3xD(33)(0);
  VNStageIntLLRInputS3xD(85)(0) <= CNStageIntLLROutputS3xD(33)(1);
  VNStageIntLLRInputS3xD(149)(0) <= CNStageIntLLROutputS3xD(33)(2);
  VNStageIntLLRInputS3xD(213)(0) <= CNStageIntLLROutputS3xD(33)(3);
  VNStageIntLLRInputS3xD(277)(0) <= CNStageIntLLROutputS3xD(33)(4);
  VNStageIntLLRInputS3xD(341)(0) <= CNStageIntLLROutputS3xD(33)(5);
  VNStageIntLLRInputS3xD(20)(0) <= CNStageIntLLROutputS3xD(34)(0);
  VNStageIntLLRInputS3xD(84)(0) <= CNStageIntLLROutputS3xD(34)(1);
  VNStageIntLLRInputS3xD(148)(0) <= CNStageIntLLROutputS3xD(34)(2);
  VNStageIntLLRInputS3xD(212)(0) <= CNStageIntLLROutputS3xD(34)(3);
  VNStageIntLLRInputS3xD(276)(0) <= CNStageIntLLROutputS3xD(34)(4);
  VNStageIntLLRInputS3xD(340)(0) <= CNStageIntLLROutputS3xD(34)(5);
  VNStageIntLLRInputS3xD(19)(0) <= CNStageIntLLROutputS3xD(35)(0);
  VNStageIntLLRInputS3xD(83)(0) <= CNStageIntLLROutputS3xD(35)(1);
  VNStageIntLLRInputS3xD(147)(0) <= CNStageIntLLROutputS3xD(35)(2);
  VNStageIntLLRInputS3xD(211)(0) <= CNStageIntLLROutputS3xD(35)(3);
  VNStageIntLLRInputS3xD(275)(0) <= CNStageIntLLROutputS3xD(35)(4);
  VNStageIntLLRInputS3xD(339)(0) <= CNStageIntLLROutputS3xD(35)(5);
  VNStageIntLLRInputS3xD(18)(0) <= CNStageIntLLROutputS3xD(36)(0);
  VNStageIntLLRInputS3xD(82)(0) <= CNStageIntLLROutputS3xD(36)(1);
  VNStageIntLLRInputS3xD(146)(0) <= CNStageIntLLROutputS3xD(36)(2);
  VNStageIntLLRInputS3xD(210)(0) <= CNStageIntLLROutputS3xD(36)(3);
  VNStageIntLLRInputS3xD(274)(0) <= CNStageIntLLROutputS3xD(36)(4);
  VNStageIntLLRInputS3xD(338)(0) <= CNStageIntLLROutputS3xD(36)(5);
  VNStageIntLLRInputS3xD(17)(0) <= CNStageIntLLROutputS3xD(37)(0);
  VNStageIntLLRInputS3xD(81)(0) <= CNStageIntLLROutputS3xD(37)(1);
  VNStageIntLLRInputS3xD(145)(0) <= CNStageIntLLROutputS3xD(37)(2);
  VNStageIntLLRInputS3xD(209)(0) <= CNStageIntLLROutputS3xD(37)(3);
  VNStageIntLLRInputS3xD(273)(0) <= CNStageIntLLROutputS3xD(37)(4);
  VNStageIntLLRInputS3xD(337)(0) <= CNStageIntLLROutputS3xD(37)(5);
  VNStageIntLLRInputS3xD(16)(0) <= CNStageIntLLROutputS3xD(38)(0);
  VNStageIntLLRInputS3xD(80)(0) <= CNStageIntLLROutputS3xD(38)(1);
  VNStageIntLLRInputS3xD(144)(0) <= CNStageIntLLROutputS3xD(38)(2);
  VNStageIntLLRInputS3xD(208)(0) <= CNStageIntLLROutputS3xD(38)(3);
  VNStageIntLLRInputS3xD(272)(0) <= CNStageIntLLROutputS3xD(38)(4);
  VNStageIntLLRInputS3xD(336)(0) <= CNStageIntLLROutputS3xD(38)(5);
  VNStageIntLLRInputS3xD(15)(0) <= CNStageIntLLROutputS3xD(39)(0);
  VNStageIntLLRInputS3xD(79)(0) <= CNStageIntLLROutputS3xD(39)(1);
  VNStageIntLLRInputS3xD(143)(0) <= CNStageIntLLROutputS3xD(39)(2);
  VNStageIntLLRInputS3xD(207)(0) <= CNStageIntLLROutputS3xD(39)(3);
  VNStageIntLLRInputS3xD(271)(0) <= CNStageIntLLROutputS3xD(39)(4);
  VNStageIntLLRInputS3xD(335)(0) <= CNStageIntLLROutputS3xD(39)(5);
  VNStageIntLLRInputS3xD(14)(0) <= CNStageIntLLROutputS3xD(40)(0);
  VNStageIntLLRInputS3xD(78)(0) <= CNStageIntLLROutputS3xD(40)(1);
  VNStageIntLLRInputS3xD(142)(0) <= CNStageIntLLROutputS3xD(40)(2);
  VNStageIntLLRInputS3xD(206)(0) <= CNStageIntLLROutputS3xD(40)(3);
  VNStageIntLLRInputS3xD(270)(0) <= CNStageIntLLROutputS3xD(40)(4);
  VNStageIntLLRInputS3xD(334)(0) <= CNStageIntLLROutputS3xD(40)(5);
  VNStageIntLLRInputS3xD(12)(0) <= CNStageIntLLROutputS3xD(41)(0);
  VNStageIntLLRInputS3xD(76)(0) <= CNStageIntLLROutputS3xD(41)(1);
  VNStageIntLLRInputS3xD(140)(0) <= CNStageIntLLROutputS3xD(41)(2);
  VNStageIntLLRInputS3xD(204)(0) <= CNStageIntLLROutputS3xD(41)(3);
  VNStageIntLLRInputS3xD(268)(0) <= CNStageIntLLROutputS3xD(41)(4);
  VNStageIntLLRInputS3xD(332)(0) <= CNStageIntLLROutputS3xD(41)(5);
  VNStageIntLLRInputS3xD(11)(0) <= CNStageIntLLROutputS3xD(42)(0);
  VNStageIntLLRInputS3xD(75)(0) <= CNStageIntLLROutputS3xD(42)(1);
  VNStageIntLLRInputS3xD(139)(0) <= CNStageIntLLROutputS3xD(42)(2);
  VNStageIntLLRInputS3xD(203)(0) <= CNStageIntLLROutputS3xD(42)(3);
  VNStageIntLLRInputS3xD(267)(0) <= CNStageIntLLROutputS3xD(42)(4);
  VNStageIntLLRInputS3xD(331)(0) <= CNStageIntLLROutputS3xD(42)(5);
  VNStageIntLLRInputS3xD(10)(0) <= CNStageIntLLROutputS3xD(43)(0);
  VNStageIntLLRInputS3xD(74)(0) <= CNStageIntLLROutputS3xD(43)(1);
  VNStageIntLLRInputS3xD(138)(0) <= CNStageIntLLROutputS3xD(43)(2);
  VNStageIntLLRInputS3xD(202)(0) <= CNStageIntLLROutputS3xD(43)(3);
  VNStageIntLLRInputS3xD(266)(0) <= CNStageIntLLROutputS3xD(43)(4);
  VNStageIntLLRInputS3xD(330)(0) <= CNStageIntLLROutputS3xD(43)(5);
  VNStageIntLLRInputS3xD(9)(0) <= CNStageIntLLROutputS3xD(44)(0);
  VNStageIntLLRInputS3xD(73)(0) <= CNStageIntLLROutputS3xD(44)(1);
  VNStageIntLLRInputS3xD(137)(0) <= CNStageIntLLROutputS3xD(44)(2);
  VNStageIntLLRInputS3xD(201)(0) <= CNStageIntLLROutputS3xD(44)(3);
  VNStageIntLLRInputS3xD(265)(0) <= CNStageIntLLROutputS3xD(44)(4);
  VNStageIntLLRInputS3xD(329)(0) <= CNStageIntLLROutputS3xD(44)(5);
  VNStageIntLLRInputS3xD(8)(0) <= CNStageIntLLROutputS3xD(45)(0);
  VNStageIntLLRInputS3xD(72)(0) <= CNStageIntLLROutputS3xD(45)(1);
  VNStageIntLLRInputS3xD(136)(0) <= CNStageIntLLROutputS3xD(45)(2);
  VNStageIntLLRInputS3xD(200)(0) <= CNStageIntLLROutputS3xD(45)(3);
  VNStageIntLLRInputS3xD(264)(0) <= CNStageIntLLROutputS3xD(45)(4);
  VNStageIntLLRInputS3xD(328)(0) <= CNStageIntLLROutputS3xD(45)(5);
  VNStageIntLLRInputS3xD(7)(0) <= CNStageIntLLROutputS3xD(46)(0);
  VNStageIntLLRInputS3xD(71)(0) <= CNStageIntLLROutputS3xD(46)(1);
  VNStageIntLLRInputS3xD(135)(0) <= CNStageIntLLROutputS3xD(46)(2);
  VNStageIntLLRInputS3xD(199)(0) <= CNStageIntLLROutputS3xD(46)(3);
  VNStageIntLLRInputS3xD(263)(0) <= CNStageIntLLROutputS3xD(46)(4);
  VNStageIntLLRInputS3xD(327)(0) <= CNStageIntLLROutputS3xD(46)(5);
  VNStageIntLLRInputS3xD(6)(0) <= CNStageIntLLROutputS3xD(47)(0);
  VNStageIntLLRInputS3xD(70)(0) <= CNStageIntLLROutputS3xD(47)(1);
  VNStageIntLLRInputS3xD(134)(0) <= CNStageIntLLROutputS3xD(47)(2);
  VNStageIntLLRInputS3xD(198)(0) <= CNStageIntLLROutputS3xD(47)(3);
  VNStageIntLLRInputS3xD(262)(0) <= CNStageIntLLROutputS3xD(47)(4);
  VNStageIntLLRInputS3xD(326)(0) <= CNStageIntLLROutputS3xD(47)(5);
  VNStageIntLLRInputS3xD(5)(0) <= CNStageIntLLROutputS3xD(48)(0);
  VNStageIntLLRInputS3xD(69)(0) <= CNStageIntLLROutputS3xD(48)(1);
  VNStageIntLLRInputS3xD(133)(0) <= CNStageIntLLROutputS3xD(48)(2);
  VNStageIntLLRInputS3xD(197)(0) <= CNStageIntLLROutputS3xD(48)(3);
  VNStageIntLLRInputS3xD(261)(0) <= CNStageIntLLROutputS3xD(48)(4);
  VNStageIntLLRInputS3xD(325)(0) <= CNStageIntLLROutputS3xD(48)(5);
  VNStageIntLLRInputS3xD(4)(0) <= CNStageIntLLROutputS3xD(49)(0);
  VNStageIntLLRInputS3xD(68)(0) <= CNStageIntLLROutputS3xD(49)(1);
  VNStageIntLLRInputS3xD(132)(0) <= CNStageIntLLROutputS3xD(49)(2);
  VNStageIntLLRInputS3xD(196)(0) <= CNStageIntLLROutputS3xD(49)(3);
  VNStageIntLLRInputS3xD(260)(0) <= CNStageIntLLROutputS3xD(49)(4);
  VNStageIntLLRInputS3xD(324)(0) <= CNStageIntLLROutputS3xD(49)(5);
  VNStageIntLLRInputS3xD(2)(0) <= CNStageIntLLROutputS3xD(50)(0);
  VNStageIntLLRInputS3xD(66)(0) <= CNStageIntLLROutputS3xD(50)(1);
  VNStageIntLLRInputS3xD(130)(0) <= CNStageIntLLROutputS3xD(50)(2);
  VNStageIntLLRInputS3xD(194)(0) <= CNStageIntLLROutputS3xD(50)(3);
  VNStageIntLLRInputS3xD(258)(0) <= CNStageIntLLROutputS3xD(50)(4);
  VNStageIntLLRInputS3xD(322)(0) <= CNStageIntLLROutputS3xD(50)(5);
  VNStageIntLLRInputS3xD(1)(0) <= CNStageIntLLROutputS3xD(51)(0);
  VNStageIntLLRInputS3xD(65)(0) <= CNStageIntLLROutputS3xD(51)(1);
  VNStageIntLLRInputS3xD(129)(0) <= CNStageIntLLROutputS3xD(51)(2);
  VNStageIntLLRInputS3xD(193)(0) <= CNStageIntLLROutputS3xD(51)(3);
  VNStageIntLLRInputS3xD(257)(0) <= CNStageIntLLROutputS3xD(51)(4);
  VNStageIntLLRInputS3xD(321)(0) <= CNStageIntLLROutputS3xD(51)(5);
  VNStageIntLLRInputS3xD(63)(0) <= CNStageIntLLROutputS3xD(52)(0);
  VNStageIntLLRInputS3xD(127)(0) <= CNStageIntLLROutputS3xD(52)(1);
  VNStageIntLLRInputS3xD(191)(0) <= CNStageIntLLROutputS3xD(52)(2);
  VNStageIntLLRInputS3xD(255)(0) <= CNStageIntLLROutputS3xD(52)(3);
  VNStageIntLLRInputS3xD(319)(0) <= CNStageIntLLROutputS3xD(52)(4);
  VNStageIntLLRInputS3xD(383)(0) <= CNStageIntLLROutputS3xD(52)(5);
  VNStageIntLLRInputS3xD(0)(0) <= CNStageIntLLROutputS3xD(53)(0);
  VNStageIntLLRInputS3xD(64)(0) <= CNStageIntLLROutputS3xD(53)(1);
  VNStageIntLLRInputS3xD(128)(0) <= CNStageIntLLROutputS3xD(53)(2);
  VNStageIntLLRInputS3xD(192)(0) <= CNStageIntLLROutputS3xD(53)(3);
  VNStageIntLLRInputS3xD(256)(0) <= CNStageIntLLROutputS3xD(53)(4);
  VNStageIntLLRInputS3xD(320)(0) <= CNStageIntLLROutputS3xD(53)(5);
  VNStageIntLLRInputS3xD(42)(1) <= CNStageIntLLROutputS3xD(54)(0);
  VNStageIntLLRInputS3xD(112)(1) <= CNStageIntLLROutputS3xD(54)(1);
  VNStageIntLLRInputS3xD(182)(1) <= CNStageIntLLROutputS3xD(54)(2);
  VNStageIntLLRInputS3xD(203)(1) <= CNStageIntLLROutputS3xD(54)(3);
  VNStageIntLLRInputS3xD(259)(0) <= CNStageIntLLROutputS3xD(54)(4);
  VNStageIntLLRInputS3xD(361)(1) <= CNStageIntLLROutputS3xD(54)(5);
  VNStageIntLLRInputS3xD(41)(1) <= CNStageIntLLROutputS3xD(55)(0);
  VNStageIntLLRInputS3xD(117)(1) <= CNStageIntLLROutputS3xD(55)(1);
  VNStageIntLLRInputS3xD(138)(1) <= CNStageIntLLROutputS3xD(55)(2);
  VNStageIntLLRInputS3xD(194)(1) <= CNStageIntLLROutputS3xD(55)(3);
  VNStageIntLLRInputS3xD(296)(1) <= CNStageIntLLROutputS3xD(55)(4);
  VNStageIntLLRInputS3xD(362)(1) <= CNStageIntLLROutputS3xD(55)(5);
  VNStageIntLLRInputS3xD(40)(1) <= CNStageIntLLROutputS3xD(56)(0);
  VNStageIntLLRInputS3xD(73)(1) <= CNStageIntLLROutputS3xD(56)(1);
  VNStageIntLLRInputS3xD(129)(1) <= CNStageIntLLROutputS3xD(56)(2);
  VNStageIntLLRInputS3xD(231)(1) <= CNStageIntLLROutputS3xD(56)(3);
  VNStageIntLLRInputS3xD(297)(1) <= CNStageIntLLROutputS3xD(56)(4);
  VNStageIntLLRInputS3xD(323)(0) <= CNStageIntLLROutputS3xD(56)(5);
  VNStageIntLLRInputS3xD(39)(1) <= CNStageIntLLROutputS3xD(57)(0);
  VNStageIntLLRInputS3xD(127)(1) <= CNStageIntLLROutputS3xD(57)(1);
  VNStageIntLLRInputS3xD(166)(1) <= CNStageIntLLROutputS3xD(57)(2);
  VNStageIntLLRInputS3xD(232)(1) <= CNStageIntLLROutputS3xD(57)(3);
  VNStageIntLLRInputS3xD(258)(1) <= CNStageIntLLROutputS3xD(57)(4);
  VNStageIntLLRInputS3xD(344)(1) <= CNStageIntLLROutputS3xD(57)(5);
  VNStageIntLLRInputS3xD(38)(1) <= CNStageIntLLROutputS3xD(58)(0);
  VNStageIntLLRInputS3xD(101)(1) <= CNStageIntLLROutputS3xD(58)(1);
  VNStageIntLLRInputS3xD(167)(1) <= CNStageIntLLROutputS3xD(58)(2);
  VNStageIntLLRInputS3xD(193)(1) <= CNStageIntLLROutputS3xD(58)(3);
  VNStageIntLLRInputS3xD(279)(1) <= CNStageIntLLROutputS3xD(58)(4);
  VNStageIntLLRInputS3xD(340)(1) <= CNStageIntLLROutputS3xD(58)(5);
  VNStageIntLLRInputS3xD(37)(1) <= CNStageIntLLROutputS3xD(59)(0);
  VNStageIntLLRInputS3xD(102)(1) <= CNStageIntLLROutputS3xD(59)(1);
  VNStageIntLLRInputS3xD(191)(1) <= CNStageIntLLROutputS3xD(59)(2);
  VNStageIntLLRInputS3xD(214)(1) <= CNStageIntLLROutputS3xD(59)(3);
  VNStageIntLLRInputS3xD(275)(1) <= CNStageIntLLROutputS3xD(59)(4);
  VNStageIntLLRInputS3xD(355)(1) <= CNStageIntLLROutputS3xD(59)(5);
  VNStageIntLLRInputS3xD(36)(1) <= CNStageIntLLROutputS3xD(60)(0);
  VNStageIntLLRInputS3xD(126)(0) <= CNStageIntLLROutputS3xD(60)(1);
  VNStageIntLLRInputS3xD(149)(1) <= CNStageIntLLROutputS3xD(60)(2);
  VNStageIntLLRInputS3xD(210)(1) <= CNStageIntLLROutputS3xD(60)(3);
  VNStageIntLLRInputS3xD(290)(1) <= CNStageIntLLROutputS3xD(60)(4);
  VNStageIntLLRInputS3xD(381)(0) <= CNStageIntLLROutputS3xD(60)(5);
  VNStageIntLLRInputS3xD(35)(1) <= CNStageIntLLROutputS3xD(61)(0);
  VNStageIntLLRInputS3xD(84)(1) <= CNStageIntLLROutputS3xD(61)(1);
  VNStageIntLLRInputS3xD(145)(1) <= CNStageIntLLROutputS3xD(61)(2);
  VNStageIntLLRInputS3xD(225)(1) <= CNStageIntLLROutputS3xD(61)(3);
  VNStageIntLLRInputS3xD(316)(0) <= CNStageIntLLROutputS3xD(61)(4);
  VNStageIntLLRInputS3xD(357)(1) <= CNStageIntLLROutputS3xD(61)(5);
  VNStageIntLLRInputS3xD(34)(1) <= CNStageIntLLROutputS3xD(62)(0);
  VNStageIntLLRInputS3xD(80)(1) <= CNStageIntLLROutputS3xD(62)(1);
  VNStageIntLLRInputS3xD(160)(1) <= CNStageIntLLROutputS3xD(62)(2);
  VNStageIntLLRInputS3xD(251)(0) <= CNStageIntLLROutputS3xD(62)(3);
  VNStageIntLLRInputS3xD(292)(1) <= CNStageIntLLROutputS3xD(62)(4);
  VNStageIntLLRInputS3xD(326)(1) <= CNStageIntLLROutputS3xD(62)(5);
  VNStageIntLLRInputS3xD(33)(1) <= CNStageIntLLROutputS3xD(63)(0);
  VNStageIntLLRInputS3xD(95)(1) <= CNStageIntLLROutputS3xD(63)(1);
  VNStageIntLLRInputS3xD(186)(0) <= CNStageIntLLROutputS3xD(63)(2);
  VNStageIntLLRInputS3xD(227)(1) <= CNStageIntLLROutputS3xD(63)(3);
  VNStageIntLLRInputS3xD(261)(1) <= CNStageIntLLROutputS3xD(63)(4);
  VNStageIntLLRInputS3xD(342)(1) <= CNStageIntLLROutputS3xD(63)(5);
  VNStageIntLLRInputS3xD(32)(1) <= CNStageIntLLROutputS3xD(64)(0);
  VNStageIntLLRInputS3xD(121)(0) <= CNStageIntLLROutputS3xD(64)(1);
  VNStageIntLLRInputS3xD(162)(1) <= CNStageIntLLROutputS3xD(64)(2);
  VNStageIntLLRInputS3xD(196)(1) <= CNStageIntLLROutputS3xD(64)(3);
  VNStageIntLLRInputS3xD(277)(1) <= CNStageIntLLROutputS3xD(64)(4);
  VNStageIntLLRInputS3xD(375)(1) <= CNStageIntLLROutputS3xD(64)(5);
  VNStageIntLLRInputS3xD(31)(1) <= CNStageIntLLROutputS3xD(65)(0);
  VNStageIntLLRInputS3xD(97)(1) <= CNStageIntLLROutputS3xD(65)(1);
  VNStageIntLLRInputS3xD(131)(0) <= CNStageIntLLROutputS3xD(65)(2);
  VNStageIntLLRInputS3xD(212)(1) <= CNStageIntLLROutputS3xD(65)(3);
  VNStageIntLLRInputS3xD(310)(1) <= CNStageIntLLROutputS3xD(65)(4);
  VNStageIntLLRInputS3xD(321)(1) <= CNStageIntLLROutputS3xD(65)(5);
  VNStageIntLLRInputS3xD(30)(1) <= CNStageIntLLROutputS3xD(66)(0);
  VNStageIntLLRInputS3xD(66)(1) <= CNStageIntLLROutputS3xD(66)(1);
  VNStageIntLLRInputS3xD(147)(1) <= CNStageIntLLROutputS3xD(66)(2);
  VNStageIntLLRInputS3xD(245)(1) <= CNStageIntLLROutputS3xD(66)(3);
  VNStageIntLLRInputS3xD(319)(1) <= CNStageIntLLROutputS3xD(66)(4);
  VNStageIntLLRInputS3xD(334)(1) <= CNStageIntLLROutputS3xD(66)(5);
  VNStageIntLLRInputS3xD(29)(1) <= CNStageIntLLROutputS3xD(67)(0);
  VNStageIntLLRInputS3xD(82)(1) <= CNStageIntLLROutputS3xD(67)(1);
  VNStageIntLLRInputS3xD(180)(0) <= CNStageIntLLROutputS3xD(67)(2);
  VNStageIntLLRInputS3xD(254)(0) <= CNStageIntLLROutputS3xD(67)(3);
  VNStageIntLLRInputS3xD(269)(0) <= CNStageIntLLROutputS3xD(67)(4);
  VNStageIntLLRInputS3xD(376)(1) <= CNStageIntLLROutputS3xD(67)(5);
  VNStageIntLLRInputS3xD(28)(1) <= CNStageIntLLROutputS3xD(68)(0);
  VNStageIntLLRInputS3xD(115)(1) <= CNStageIntLLROutputS3xD(68)(1);
  VNStageIntLLRInputS3xD(189)(0) <= CNStageIntLLROutputS3xD(68)(2);
  VNStageIntLLRInputS3xD(204)(1) <= CNStageIntLLROutputS3xD(68)(3);
  VNStageIntLLRInputS3xD(311)(1) <= CNStageIntLLROutputS3xD(68)(4);
  VNStageIntLLRInputS3xD(341)(1) <= CNStageIntLLROutputS3xD(68)(5);
  VNStageIntLLRInputS3xD(27)(1) <= CNStageIntLLROutputS3xD(69)(0);
  VNStageIntLLRInputS3xD(124)(0) <= CNStageIntLLROutputS3xD(69)(1);
  VNStageIntLLRInputS3xD(139)(1) <= CNStageIntLLROutputS3xD(69)(2);
  VNStageIntLLRInputS3xD(246)(1) <= CNStageIntLLROutputS3xD(69)(3);
  VNStageIntLLRInputS3xD(276)(1) <= CNStageIntLLROutputS3xD(69)(4);
  VNStageIntLLRInputS3xD(343)(1) <= CNStageIntLLROutputS3xD(69)(5);
  VNStageIntLLRInputS3xD(26)(1) <= CNStageIntLLROutputS3xD(70)(0);
  VNStageIntLLRInputS3xD(74)(1) <= CNStageIntLLROutputS3xD(70)(1);
  VNStageIntLLRInputS3xD(181)(1) <= CNStageIntLLROutputS3xD(70)(2);
  VNStageIntLLRInputS3xD(211)(1) <= CNStageIntLLROutputS3xD(70)(3);
  VNStageIntLLRInputS3xD(278)(1) <= CNStageIntLLROutputS3xD(70)(4);
  VNStageIntLLRInputS3xD(325)(1) <= CNStageIntLLROutputS3xD(70)(5);
  VNStageIntLLRInputS3xD(25)(1) <= CNStageIntLLROutputS3xD(71)(0);
  VNStageIntLLRInputS3xD(116)(0) <= CNStageIntLLROutputS3xD(71)(1);
  VNStageIntLLRInputS3xD(146)(1) <= CNStageIntLLROutputS3xD(71)(2);
  VNStageIntLLRInputS3xD(213)(1) <= CNStageIntLLROutputS3xD(71)(3);
  VNStageIntLLRInputS3xD(260)(1) <= CNStageIntLLROutputS3xD(71)(4);
  VNStageIntLLRInputS3xD(332)(1) <= CNStageIntLLROutputS3xD(71)(5);
  VNStageIntLLRInputS3xD(24)(1) <= CNStageIntLLROutputS3xD(72)(0);
  VNStageIntLLRInputS3xD(81)(1) <= CNStageIntLLROutputS3xD(72)(1);
  VNStageIntLLRInputS3xD(148)(1) <= CNStageIntLLROutputS3xD(72)(2);
  VNStageIntLLRInputS3xD(195)(0) <= CNStageIntLLROutputS3xD(72)(3);
  VNStageIntLLRInputS3xD(267)(1) <= CNStageIntLLROutputS3xD(72)(4);
  VNStageIntLLRInputS3xD(359)(1) <= CNStageIntLLROutputS3xD(72)(5);
  VNStageIntLLRInputS3xD(23)(1) <= CNStageIntLLROutputS3xD(73)(0);
  VNStageIntLLRInputS3xD(83)(1) <= CNStageIntLLROutputS3xD(73)(1);
  VNStageIntLLRInputS3xD(130)(1) <= CNStageIntLLROutputS3xD(73)(2);
  VNStageIntLLRInputS3xD(202)(1) <= CNStageIntLLROutputS3xD(73)(3);
  VNStageIntLLRInputS3xD(294)(1) <= CNStageIntLLROutputS3xD(73)(4);
  VNStageIntLLRInputS3xD(347)(1) <= CNStageIntLLROutputS3xD(73)(5);
  VNStageIntLLRInputS3xD(22)(1) <= CNStageIntLLROutputS3xD(74)(0);
  VNStageIntLLRInputS3xD(65)(1) <= CNStageIntLLROutputS3xD(74)(1);
  VNStageIntLLRInputS3xD(137)(1) <= CNStageIntLLROutputS3xD(74)(2);
  VNStageIntLLRInputS3xD(229)(1) <= CNStageIntLLROutputS3xD(74)(3);
  VNStageIntLLRInputS3xD(282)(1) <= CNStageIntLLROutputS3xD(74)(4);
  VNStageIntLLRInputS3xD(353)(1) <= CNStageIntLLROutputS3xD(74)(5);
  VNStageIntLLRInputS3xD(21)(1) <= CNStageIntLLROutputS3xD(75)(0);
  VNStageIntLLRInputS3xD(72)(1) <= CNStageIntLLROutputS3xD(75)(1);
  VNStageIntLLRInputS3xD(164)(1) <= CNStageIntLLROutputS3xD(75)(2);
  VNStageIntLLRInputS3xD(217)(1) <= CNStageIntLLROutputS3xD(75)(3);
  VNStageIntLLRInputS3xD(288)(1) <= CNStageIntLLROutputS3xD(75)(4);
  VNStageIntLLRInputS3xD(348)(1) <= CNStageIntLLROutputS3xD(75)(5);
  VNStageIntLLRInputS3xD(20)(1) <= CNStageIntLLROutputS3xD(76)(0);
  VNStageIntLLRInputS3xD(99)(1) <= CNStageIntLLROutputS3xD(76)(1);
  VNStageIntLLRInputS3xD(152)(1) <= CNStageIntLLROutputS3xD(76)(2);
  VNStageIntLLRInputS3xD(223)(1) <= CNStageIntLLROutputS3xD(76)(3);
  VNStageIntLLRInputS3xD(283)(1) <= CNStageIntLLROutputS3xD(76)(4);
  VNStageIntLLRInputS3xD(358)(1) <= CNStageIntLLROutputS3xD(76)(5);
  VNStageIntLLRInputS3xD(19)(1) <= CNStageIntLLROutputS3xD(77)(0);
  VNStageIntLLRInputS3xD(87)(1) <= CNStageIntLLROutputS3xD(77)(1);
  VNStageIntLLRInputS3xD(158)(1) <= CNStageIntLLROutputS3xD(77)(2);
  VNStageIntLLRInputS3xD(218)(1) <= CNStageIntLLROutputS3xD(77)(3);
  VNStageIntLLRInputS3xD(293)(1) <= CNStageIntLLROutputS3xD(77)(4);
  VNStageIntLLRInputS3xD(380)(0) <= CNStageIntLLROutputS3xD(77)(5);
  VNStageIntLLRInputS3xD(18)(1) <= CNStageIntLLROutputS3xD(78)(0);
  VNStageIntLLRInputS3xD(93)(1) <= CNStageIntLLROutputS3xD(78)(1);
  VNStageIntLLRInputS3xD(153)(1) <= CNStageIntLLROutputS3xD(78)(2);
  VNStageIntLLRInputS3xD(228)(1) <= CNStageIntLLROutputS3xD(78)(3);
  VNStageIntLLRInputS3xD(315)(0) <= CNStageIntLLROutputS3xD(78)(4);
  VNStageIntLLRInputS3xD(335)(1) <= CNStageIntLLROutputS3xD(78)(5);
  VNStageIntLLRInputS3xD(17)(1) <= CNStageIntLLROutputS3xD(79)(0);
  VNStageIntLLRInputS3xD(88)(1) <= CNStageIntLLROutputS3xD(79)(1);
  VNStageIntLLRInputS3xD(163)(1) <= CNStageIntLLROutputS3xD(79)(2);
  VNStageIntLLRInputS3xD(250)(0) <= CNStageIntLLROutputS3xD(79)(3);
  VNStageIntLLRInputS3xD(270)(1) <= CNStageIntLLROutputS3xD(79)(4);
  VNStageIntLLRInputS3xD(383)(1) <= CNStageIntLLROutputS3xD(79)(5);
  VNStageIntLLRInputS3xD(15)(1) <= CNStageIntLLROutputS3xD(80)(0);
  VNStageIntLLRInputS3xD(120)(1) <= CNStageIntLLROutputS3xD(80)(1);
  VNStageIntLLRInputS3xD(140)(1) <= CNStageIntLLROutputS3xD(80)(2);
  VNStageIntLLRInputS3xD(253)(0) <= CNStageIntLLROutputS3xD(80)(3);
  VNStageIntLLRInputS3xD(305)(1) <= CNStageIntLLROutputS3xD(80)(4);
  VNStageIntLLRInputS3xD(338)(1) <= CNStageIntLLROutputS3xD(80)(5);
  VNStageIntLLRInputS3xD(14)(1) <= CNStageIntLLROutputS3xD(81)(0);
  VNStageIntLLRInputS3xD(75)(1) <= CNStageIntLLROutputS3xD(81)(1);
  VNStageIntLLRInputS3xD(188)(0) <= CNStageIntLLROutputS3xD(81)(2);
  VNStageIntLLRInputS3xD(240)(1) <= CNStageIntLLROutputS3xD(81)(3);
  VNStageIntLLRInputS3xD(273)(1) <= CNStageIntLLROutputS3xD(81)(4);
  VNStageIntLLRInputS3xD(350)(1) <= CNStageIntLLROutputS3xD(81)(5);
  VNStageIntLLRInputS3xD(13)(0) <= CNStageIntLLROutputS3xD(82)(0);
  VNStageIntLLRInputS3xD(123)(0) <= CNStageIntLLROutputS3xD(82)(1);
  VNStageIntLLRInputS3xD(175)(1) <= CNStageIntLLROutputS3xD(82)(2);
  VNStageIntLLRInputS3xD(208)(1) <= CNStageIntLLROutputS3xD(82)(3);
  VNStageIntLLRInputS3xD(285)(1) <= CNStageIntLLROutputS3xD(82)(4);
  VNStageIntLLRInputS3xD(364)(1) <= CNStageIntLLROutputS3xD(82)(5);
  VNStageIntLLRInputS3xD(12)(1) <= CNStageIntLLROutputS3xD(83)(0);
  VNStageIntLLRInputS3xD(110)(1) <= CNStageIntLLROutputS3xD(83)(1);
  VNStageIntLLRInputS3xD(143)(1) <= CNStageIntLLROutputS3xD(83)(2);
  VNStageIntLLRInputS3xD(220)(1) <= CNStageIntLLROutputS3xD(83)(3);
  VNStageIntLLRInputS3xD(299)(0) <= CNStageIntLLROutputS3xD(83)(4);
  VNStageIntLLRInputS3xD(345)(1) <= CNStageIntLLROutputS3xD(83)(5);
  VNStageIntLLRInputS3xD(11)(1) <= CNStageIntLLROutputS3xD(84)(0);
  VNStageIntLLRInputS3xD(78)(1) <= CNStageIntLLROutputS3xD(84)(1);
  VNStageIntLLRInputS3xD(155)(1) <= CNStageIntLLROutputS3xD(84)(2);
  VNStageIntLLRInputS3xD(234)(1) <= CNStageIntLLROutputS3xD(84)(3);
  VNStageIntLLRInputS3xD(280)(1) <= CNStageIntLLROutputS3xD(84)(4);
  VNStageIntLLRInputS3xD(322)(1) <= CNStageIntLLROutputS3xD(84)(5);
  VNStageIntLLRInputS3xD(10)(1) <= CNStageIntLLROutputS3xD(85)(0);
  VNStageIntLLRInputS3xD(90)(1) <= CNStageIntLLROutputS3xD(85)(1);
  VNStageIntLLRInputS3xD(169)(1) <= CNStageIntLLROutputS3xD(85)(2);
  VNStageIntLLRInputS3xD(215)(1) <= CNStageIntLLROutputS3xD(85)(3);
  VNStageIntLLRInputS3xD(257)(1) <= CNStageIntLLROutputS3xD(85)(4);
  VNStageIntLLRInputS3xD(374)(1) <= CNStageIntLLROutputS3xD(85)(5);
  VNStageIntLLRInputS3xD(9)(1) <= CNStageIntLLROutputS3xD(86)(0);
  VNStageIntLLRInputS3xD(104)(1) <= CNStageIntLLROutputS3xD(86)(1);
  VNStageIntLLRInputS3xD(150)(1) <= CNStageIntLLROutputS3xD(86)(2);
  VNStageIntLLRInputS3xD(255)(1) <= CNStageIntLLROutputS3xD(86)(3);
  VNStageIntLLRInputS3xD(309)(1) <= CNStageIntLLROutputS3xD(86)(4);
  VNStageIntLLRInputS3xD(378)(0) <= CNStageIntLLROutputS3xD(86)(5);
  VNStageIntLLRInputS3xD(7)(1) <= CNStageIntLLROutputS3xD(87)(0);
  VNStageIntLLRInputS3xD(125)(0) <= CNStageIntLLROutputS3xD(87)(1);
  VNStageIntLLRInputS3xD(179)(1) <= CNStageIntLLROutputS3xD(87)(2);
  VNStageIntLLRInputS3xD(248)(1) <= CNStageIntLLROutputS3xD(87)(3);
  VNStageIntLLRInputS3xD(306)(1) <= CNStageIntLLROutputS3xD(87)(4);
  VNStageIntLLRInputS3xD(382)(0) <= CNStageIntLLROutputS3xD(87)(5);
  VNStageIntLLRInputS3xD(6)(1) <= CNStageIntLLROutputS3xD(88)(0);
  VNStageIntLLRInputS3xD(114)(1) <= CNStageIntLLROutputS3xD(88)(1);
  VNStageIntLLRInputS3xD(183)(1) <= CNStageIntLLROutputS3xD(88)(2);
  VNStageIntLLRInputS3xD(241)(1) <= CNStageIntLLROutputS3xD(88)(3);
  VNStageIntLLRInputS3xD(317)(0) <= CNStageIntLLROutputS3xD(88)(4);
  VNStageIntLLRInputS3xD(354)(1) <= CNStageIntLLROutputS3xD(88)(5);
  VNStageIntLLRInputS3xD(5)(1) <= CNStageIntLLROutputS3xD(89)(0);
  VNStageIntLLRInputS3xD(118)(1) <= CNStageIntLLROutputS3xD(89)(1);
  VNStageIntLLRInputS3xD(176)(1) <= CNStageIntLLROutputS3xD(89)(2);
  VNStageIntLLRInputS3xD(252)(0) <= CNStageIntLLROutputS3xD(89)(3);
  VNStageIntLLRInputS3xD(289)(1) <= CNStageIntLLROutputS3xD(89)(4);
  VNStageIntLLRInputS3xD(346)(1) <= CNStageIntLLROutputS3xD(89)(5);
  VNStageIntLLRInputS3xD(4)(1) <= CNStageIntLLROutputS3xD(90)(0);
  VNStageIntLLRInputS3xD(111)(1) <= CNStageIntLLROutputS3xD(90)(1);
  VNStageIntLLRInputS3xD(187)(0) <= CNStageIntLLROutputS3xD(90)(2);
  VNStageIntLLRInputS3xD(224)(1) <= CNStageIntLLROutputS3xD(90)(3);
  VNStageIntLLRInputS3xD(281)(1) <= CNStageIntLLROutputS3xD(90)(4);
  VNStageIntLLRInputS3xD(363)(0) <= CNStageIntLLROutputS3xD(90)(5);
  VNStageIntLLRInputS3xD(3)(0) <= CNStageIntLLROutputS3xD(91)(0);
  VNStageIntLLRInputS3xD(122)(0) <= CNStageIntLLROutputS3xD(91)(1);
  VNStageIntLLRInputS3xD(159)(1) <= CNStageIntLLROutputS3xD(91)(2);
  VNStageIntLLRInputS3xD(216)(1) <= CNStageIntLLROutputS3xD(91)(3);
  VNStageIntLLRInputS3xD(298)(1) <= CNStageIntLLROutputS3xD(91)(4);
  VNStageIntLLRInputS3xD(360)(1) <= CNStageIntLLROutputS3xD(91)(5);
  VNStageIntLLRInputS3xD(2)(1) <= CNStageIntLLROutputS3xD(92)(0);
  VNStageIntLLRInputS3xD(94)(1) <= CNStageIntLLROutputS3xD(92)(1);
  VNStageIntLLRInputS3xD(151)(1) <= CNStageIntLLROutputS3xD(92)(2);
  VNStageIntLLRInputS3xD(233)(1) <= CNStageIntLLROutputS3xD(92)(3);
  VNStageIntLLRInputS3xD(295)(1) <= CNStageIntLLROutputS3xD(92)(4);
  VNStageIntLLRInputS3xD(331)(1) <= CNStageIntLLROutputS3xD(92)(5);
  VNStageIntLLRInputS3xD(63)(1) <= CNStageIntLLROutputS3xD(93)(0);
  VNStageIntLLRInputS3xD(103)(1) <= CNStageIntLLROutputS3xD(93)(1);
  VNStageIntLLRInputS3xD(165)(1) <= CNStageIntLLROutputS3xD(93)(2);
  VNStageIntLLRInputS3xD(201)(1) <= CNStageIntLLROutputS3xD(93)(3);
  VNStageIntLLRInputS3xD(286)(1) <= CNStageIntLLROutputS3xD(93)(4);
  VNStageIntLLRInputS3xD(337)(1) <= CNStageIntLLROutputS3xD(93)(5);
  VNStageIntLLRInputS3xD(62)(0) <= CNStageIntLLROutputS3xD(94)(0);
  VNStageIntLLRInputS3xD(100)(1) <= CNStageIntLLROutputS3xD(94)(1);
  VNStageIntLLRInputS3xD(136)(1) <= CNStageIntLLROutputS3xD(94)(2);
  VNStageIntLLRInputS3xD(221)(1) <= CNStageIntLLROutputS3xD(94)(3);
  VNStageIntLLRInputS3xD(272)(1) <= CNStageIntLLROutputS3xD(94)(4);
  VNStageIntLLRInputS3xD(327)(1) <= CNStageIntLLROutputS3xD(94)(5);
  VNStageIntLLRInputS3xD(61)(0) <= CNStageIntLLROutputS3xD(95)(0);
  VNStageIntLLRInputS3xD(71)(1) <= CNStageIntLLROutputS3xD(95)(1);
  VNStageIntLLRInputS3xD(156)(1) <= CNStageIntLLROutputS3xD(95)(2);
  VNStageIntLLRInputS3xD(207)(1) <= CNStageIntLLROutputS3xD(95)(3);
  VNStageIntLLRInputS3xD(262)(1) <= CNStageIntLLROutputS3xD(95)(4);
  VNStageIntLLRInputS3xD(356)(1) <= CNStageIntLLROutputS3xD(95)(5);
  VNStageIntLLRInputS3xD(60)(0) <= CNStageIntLLROutputS3xD(96)(0);
  VNStageIntLLRInputS3xD(91)(1) <= CNStageIntLLROutputS3xD(96)(1);
  VNStageIntLLRInputS3xD(142)(1) <= CNStageIntLLROutputS3xD(96)(2);
  VNStageIntLLRInputS3xD(197)(1) <= CNStageIntLLROutputS3xD(96)(3);
  VNStageIntLLRInputS3xD(291)(1) <= CNStageIntLLROutputS3xD(96)(4);
  VNStageIntLLRInputS3xD(339)(1) <= CNStageIntLLROutputS3xD(96)(5);
  VNStageIntLLRInputS3xD(58)(0) <= CNStageIntLLROutputS3xD(97)(0);
  VNStageIntLLRInputS3xD(67)(0) <= CNStageIntLLROutputS3xD(97)(1);
  VNStageIntLLRInputS3xD(161)(1) <= CNStageIntLLROutputS3xD(97)(2);
  VNStageIntLLRInputS3xD(209)(1) <= CNStageIntLLROutputS3xD(97)(3);
  VNStageIntLLRInputS3xD(304)(1) <= CNStageIntLLROutputS3xD(97)(4);
  VNStageIntLLRInputS3xD(329)(1) <= CNStageIntLLROutputS3xD(97)(5);
  VNStageIntLLRInputS3xD(57)(0) <= CNStageIntLLROutputS3xD(98)(0);
  VNStageIntLLRInputS3xD(96)(1) <= CNStageIntLLROutputS3xD(98)(1);
  VNStageIntLLRInputS3xD(144)(1) <= CNStageIntLLROutputS3xD(98)(2);
  VNStageIntLLRInputS3xD(239)(1) <= CNStageIntLLROutputS3xD(98)(3);
  VNStageIntLLRInputS3xD(264)(1) <= CNStageIntLLROutputS3xD(98)(4);
  VNStageIntLLRInputS3xD(365)(1) <= CNStageIntLLROutputS3xD(98)(5);
  VNStageIntLLRInputS3xD(56)(1) <= CNStageIntLLROutputS3xD(99)(0);
  VNStageIntLLRInputS3xD(79)(1) <= CNStageIntLLROutputS3xD(99)(1);
  VNStageIntLLRInputS3xD(174)(1) <= CNStageIntLLROutputS3xD(99)(2);
  VNStageIntLLRInputS3xD(199)(1) <= CNStageIntLLROutputS3xD(99)(3);
  VNStageIntLLRInputS3xD(300)(1) <= CNStageIntLLROutputS3xD(99)(4);
  VNStageIntLLRInputS3xD(349)(1) <= CNStageIntLLROutputS3xD(99)(5);
  VNStageIntLLRInputS3xD(55)(1) <= CNStageIntLLROutputS3xD(100)(0);
  VNStageIntLLRInputS3xD(109)(1) <= CNStageIntLLROutputS3xD(100)(1);
  VNStageIntLLRInputS3xD(134)(1) <= CNStageIntLLROutputS3xD(100)(2);
  VNStageIntLLRInputS3xD(235)(0) <= CNStageIntLLROutputS3xD(100)(3);
  VNStageIntLLRInputS3xD(284)(1) <= CNStageIntLLROutputS3xD(100)(4);
  VNStageIntLLRInputS3xD(352)(1) <= CNStageIntLLROutputS3xD(100)(5);
  VNStageIntLLRInputS3xD(54)(1) <= CNStageIntLLROutputS3xD(101)(0);
  VNStageIntLLRInputS3xD(69)(1) <= CNStageIntLLROutputS3xD(101)(1);
  VNStageIntLLRInputS3xD(170)(1) <= CNStageIntLLROutputS3xD(101)(2);
  VNStageIntLLRInputS3xD(219)(1) <= CNStageIntLLROutputS3xD(101)(3);
  VNStageIntLLRInputS3xD(287)(1) <= CNStageIntLLROutputS3xD(101)(4);
  VNStageIntLLRInputS3xD(330)(1) <= CNStageIntLLROutputS3xD(101)(5);
  VNStageIntLLRInputS3xD(52)(0) <= CNStageIntLLROutputS3xD(102)(0);
  VNStageIntLLRInputS3xD(89)(1) <= CNStageIntLLROutputS3xD(102)(1);
  VNStageIntLLRInputS3xD(157)(1) <= CNStageIntLLROutputS3xD(102)(2);
  VNStageIntLLRInputS3xD(200)(1) <= CNStageIntLLROutputS3xD(102)(3);
  VNStageIntLLRInputS3xD(303)(1) <= CNStageIntLLROutputS3xD(102)(4);
  VNStageIntLLRInputS3xD(366)(1) <= CNStageIntLLROutputS3xD(102)(5);
  VNStageIntLLRInputS3xD(51)(1) <= CNStageIntLLROutputS3xD(103)(0);
  VNStageIntLLRInputS3xD(92)(1) <= CNStageIntLLROutputS3xD(103)(1);
  VNStageIntLLRInputS3xD(135)(1) <= CNStageIntLLROutputS3xD(103)(2);
  VNStageIntLLRInputS3xD(238)(1) <= CNStageIntLLROutputS3xD(103)(3);
  VNStageIntLLRInputS3xD(301)(1) <= CNStageIntLLROutputS3xD(103)(4);
  VNStageIntLLRInputS3xD(328)(1) <= CNStageIntLLROutputS3xD(103)(5);
  VNStageIntLLRInputS3xD(50)(1) <= CNStageIntLLROutputS3xD(104)(0);
  VNStageIntLLRInputS3xD(70)(1) <= CNStageIntLLROutputS3xD(104)(1);
  VNStageIntLLRInputS3xD(173)(1) <= CNStageIntLLROutputS3xD(104)(2);
  VNStageIntLLRInputS3xD(236)(1) <= CNStageIntLLROutputS3xD(104)(3);
  VNStageIntLLRInputS3xD(263)(1) <= CNStageIntLLROutputS3xD(104)(4);
  VNStageIntLLRInputS3xD(336)(1) <= CNStageIntLLROutputS3xD(104)(5);
  VNStageIntLLRInputS3xD(49)(1) <= CNStageIntLLROutputS3xD(105)(0);
  VNStageIntLLRInputS3xD(108)(1) <= CNStageIntLLROutputS3xD(105)(1);
  VNStageIntLLRInputS3xD(171)(0) <= CNStageIntLLROutputS3xD(105)(2);
  VNStageIntLLRInputS3xD(198)(1) <= CNStageIntLLROutputS3xD(105)(3);
  VNStageIntLLRInputS3xD(271)(1) <= CNStageIntLLROutputS3xD(105)(4);
  VNStageIntLLRInputS3xD(379)(0) <= CNStageIntLLROutputS3xD(105)(5);
  VNStageIntLLRInputS3xD(46)(1) <= CNStageIntLLROutputS3xD(106)(0);
  VNStageIntLLRInputS3xD(76)(1) <= CNStageIntLLROutputS3xD(106)(1);
  VNStageIntLLRInputS3xD(184)(1) <= CNStageIntLLROutputS3xD(106)(2);
  VNStageIntLLRInputS3xD(243)(1) <= CNStageIntLLROutputS3xD(106)(3);
  VNStageIntLLRInputS3xD(256)(1) <= CNStageIntLLROutputS3xD(106)(4);
  VNStageIntLLRInputS3xD(372)(0) <= CNStageIntLLROutputS3xD(106)(5);
  VNStageIntLLRInputS3xD(45)(1) <= CNStageIntLLROutputS3xD(107)(0);
  VNStageIntLLRInputS3xD(119)(1) <= CNStageIntLLROutputS3xD(107)(1);
  VNStageIntLLRInputS3xD(178)(1) <= CNStageIntLLROutputS3xD(107)(2);
  VNStageIntLLRInputS3xD(192)(1) <= CNStageIntLLROutputS3xD(107)(3);
  VNStageIntLLRInputS3xD(307)(1) <= CNStageIntLLROutputS3xD(107)(4);
  VNStageIntLLRInputS3xD(377)(0) <= CNStageIntLLROutputS3xD(107)(5);
  VNStageIntLLRInputS3xD(44)(1) <= CNStageIntLLROutputS3xD(108)(0);
  VNStageIntLLRInputS3xD(113)(1) <= CNStageIntLLROutputS3xD(108)(1);
  VNStageIntLLRInputS3xD(128)(1) <= CNStageIntLLROutputS3xD(108)(2);
  VNStageIntLLRInputS3xD(242)(1) <= CNStageIntLLROutputS3xD(108)(3);
  VNStageIntLLRInputS3xD(312)(1) <= CNStageIntLLROutputS3xD(108)(4);
  VNStageIntLLRInputS3xD(333)(0) <= CNStageIntLLROutputS3xD(108)(5);
  VNStageIntLLRInputS3xD(43)(0) <= CNStageIntLLROutputS3xD(109)(0);
  VNStageIntLLRInputS3xD(64)(1) <= CNStageIntLLROutputS3xD(109)(1);
  VNStageIntLLRInputS3xD(177)(1) <= CNStageIntLLROutputS3xD(109)(2);
  VNStageIntLLRInputS3xD(247)(1) <= CNStageIntLLROutputS3xD(109)(3);
  VNStageIntLLRInputS3xD(268)(1) <= CNStageIntLLROutputS3xD(109)(4);
  VNStageIntLLRInputS3xD(324)(1) <= CNStageIntLLROutputS3xD(109)(5);
  VNStageIntLLRInputS3xD(0)(1) <= CNStageIntLLROutputS3xD(110)(0);
  VNStageIntLLRInputS3xD(107)(0) <= CNStageIntLLROutputS3xD(110)(1);
  VNStageIntLLRInputS3xD(172)(1) <= CNStageIntLLROutputS3xD(110)(2);
  VNStageIntLLRInputS3xD(237)(1) <= CNStageIntLLROutputS3xD(110)(3);
  VNStageIntLLRInputS3xD(302)(1) <= CNStageIntLLROutputS3xD(110)(4);
  VNStageIntLLRInputS3xD(367)(1) <= CNStageIntLLROutputS3xD(110)(5);
  VNStageIntLLRInputS3xD(32)(2) <= CNStageIntLLROutputS3xD(111)(0);
  VNStageIntLLRInputS3xD(117)(2) <= CNStageIntLLROutputS3xD(111)(1);
  VNStageIntLLRInputS3xD(136)(2) <= CNStageIntLLROutputS3xD(111)(2);
  VNStageIntLLRInputS3xD(198)(2) <= CNStageIntLLROutputS3xD(111)(3);
  VNStageIntLLRInputS3xD(297)(2) <= CNStageIntLLROutputS3xD(111)(4);
  VNStageIntLLRInputS3xD(382)(1) <= CNStageIntLLROutputS3xD(111)(5);
  VNStageIntLLRInputS3xD(30)(2) <= CNStageIntLLROutputS3xD(112)(0);
  VNStageIntLLRInputS3xD(68)(1) <= CNStageIntLLROutputS3xD(112)(1);
  VNStageIntLLRInputS3xD(167)(2) <= CNStageIntLLROutputS3xD(112)(2);
  VNStageIntLLRInputS3xD(252)(1) <= CNStageIntLLROutputS3xD(112)(3);
  VNStageIntLLRInputS3xD(303)(2) <= CNStageIntLLROutputS3xD(112)(4);
  VNStageIntLLRInputS3xD(358)(2) <= CNStageIntLLROutputS3xD(112)(5);
  VNStageIntLLRInputS3xD(29)(2) <= CNStageIntLLROutputS3xD(113)(0);
  VNStageIntLLRInputS3xD(102)(2) <= CNStageIntLLROutputS3xD(113)(1);
  VNStageIntLLRInputS3xD(187)(1) <= CNStageIntLLROutputS3xD(113)(2);
  VNStageIntLLRInputS3xD(238)(2) <= CNStageIntLLROutputS3xD(113)(3);
  VNStageIntLLRInputS3xD(293)(2) <= CNStageIntLLROutputS3xD(113)(4);
  VNStageIntLLRInputS3xD(324)(2) <= CNStageIntLLROutputS3xD(113)(5);
  VNStageIntLLRInputS3xD(28)(2) <= CNStageIntLLROutputS3xD(114)(0);
  VNStageIntLLRInputS3xD(122)(1) <= CNStageIntLLROutputS3xD(114)(1);
  VNStageIntLLRInputS3xD(173)(2) <= CNStageIntLLROutputS3xD(114)(2);
  VNStageIntLLRInputS3xD(228)(2) <= CNStageIntLLROutputS3xD(114)(3);
  VNStageIntLLRInputS3xD(259)(1) <= CNStageIntLLROutputS3xD(114)(4);
  VNStageIntLLRInputS3xD(370)(1) <= CNStageIntLLROutputS3xD(114)(5);
  VNStageIntLLRInputS3xD(27)(2) <= CNStageIntLLROutputS3xD(115)(0);
  VNStageIntLLRInputS3xD(108)(2) <= CNStageIntLLROutputS3xD(115)(1);
  VNStageIntLLRInputS3xD(163)(2) <= CNStageIntLLROutputS3xD(115)(2);
  VNStageIntLLRInputS3xD(194)(2) <= CNStageIntLLROutputS3xD(115)(3);
  VNStageIntLLRInputS3xD(305)(2) <= CNStageIntLLROutputS3xD(115)(4);
  VNStageIntLLRInputS3xD(337)(2) <= CNStageIntLLROutputS3xD(115)(5);
  VNStageIntLLRInputS3xD(26)(2) <= CNStageIntLLROutputS3xD(116)(0);
  VNStageIntLLRInputS3xD(98)(1) <= CNStageIntLLROutputS3xD(116)(1);
  VNStageIntLLRInputS3xD(129)(2) <= CNStageIntLLROutputS3xD(116)(2);
  VNStageIntLLRInputS3xD(240)(2) <= CNStageIntLLROutputS3xD(116)(3);
  VNStageIntLLRInputS3xD(272)(2) <= CNStageIntLLROutputS3xD(116)(4);
  VNStageIntLLRInputS3xD(360)(2) <= CNStageIntLLROutputS3xD(116)(5);
  VNStageIntLLRInputS3xD(25)(2) <= CNStageIntLLROutputS3xD(117)(0);
  VNStageIntLLRInputS3xD(127)(2) <= CNStageIntLLROutputS3xD(117)(1);
  VNStageIntLLRInputS3xD(175)(2) <= CNStageIntLLROutputS3xD(117)(2);
  VNStageIntLLRInputS3xD(207)(2) <= CNStageIntLLROutputS3xD(117)(3);
  VNStageIntLLRInputS3xD(295)(2) <= CNStageIntLLROutputS3xD(117)(4);
  VNStageIntLLRInputS3xD(333)(1) <= CNStageIntLLROutputS3xD(117)(5);
  VNStageIntLLRInputS3xD(24)(2) <= CNStageIntLLROutputS3xD(118)(0);
  VNStageIntLLRInputS3xD(110)(2) <= CNStageIntLLROutputS3xD(118)(1);
  VNStageIntLLRInputS3xD(142)(2) <= CNStageIntLLROutputS3xD(118)(2);
  VNStageIntLLRInputS3xD(230)(1) <= CNStageIntLLROutputS3xD(118)(3);
  VNStageIntLLRInputS3xD(268)(2) <= CNStageIntLLROutputS3xD(118)(4);
  VNStageIntLLRInputS3xD(380)(1) <= CNStageIntLLROutputS3xD(118)(5);
  VNStageIntLLRInputS3xD(23)(2) <= CNStageIntLLROutputS3xD(119)(0);
  VNStageIntLLRInputS3xD(77)(0) <= CNStageIntLLROutputS3xD(119)(1);
  VNStageIntLLRInputS3xD(165)(2) <= CNStageIntLLROutputS3xD(119)(2);
  VNStageIntLLRInputS3xD(203)(2) <= CNStageIntLLROutputS3xD(119)(3);
  VNStageIntLLRInputS3xD(315)(1) <= CNStageIntLLROutputS3xD(119)(4);
  VNStageIntLLRInputS3xD(383)(2) <= CNStageIntLLROutputS3xD(119)(5);
  VNStageIntLLRInputS3xD(22)(2) <= CNStageIntLLROutputS3xD(120)(0);
  VNStageIntLLRInputS3xD(100)(2) <= CNStageIntLLROutputS3xD(120)(1);
  VNStageIntLLRInputS3xD(138)(2) <= CNStageIntLLROutputS3xD(120)(2);
  VNStageIntLLRInputS3xD(250)(1) <= CNStageIntLLROutputS3xD(120)(3);
  VNStageIntLLRInputS3xD(318)(0) <= CNStageIntLLROutputS3xD(120)(4);
  VNStageIntLLRInputS3xD(361)(2) <= CNStageIntLLROutputS3xD(120)(5);
  VNStageIntLLRInputS3xD(21)(2) <= CNStageIntLLROutputS3xD(121)(0);
  VNStageIntLLRInputS3xD(73)(2) <= CNStageIntLLROutputS3xD(121)(1);
  VNStageIntLLRInputS3xD(185)(0) <= CNStageIntLLROutputS3xD(121)(2);
  VNStageIntLLRInputS3xD(253)(1) <= CNStageIntLLROutputS3xD(121)(3);
  VNStageIntLLRInputS3xD(296)(2) <= CNStageIntLLROutputS3xD(121)(4);
  VNStageIntLLRInputS3xD(336)(2) <= CNStageIntLLROutputS3xD(121)(5);
  VNStageIntLLRInputS3xD(19)(2) <= CNStageIntLLROutputS3xD(122)(0);
  VNStageIntLLRInputS3xD(123)(1) <= CNStageIntLLROutputS3xD(122)(1);
  VNStageIntLLRInputS3xD(166)(2) <= CNStageIntLLROutputS3xD(122)(2);
  VNStageIntLLRInputS3xD(206)(1) <= CNStageIntLLROutputS3xD(122)(3);
  VNStageIntLLRInputS3xD(269)(1) <= CNStageIntLLROutputS3xD(122)(4);
  VNStageIntLLRInputS3xD(359)(2) <= CNStageIntLLROutputS3xD(122)(5);
  VNStageIntLLRInputS3xD(18)(2) <= CNStageIntLLROutputS3xD(123)(0);
  VNStageIntLLRInputS3xD(101)(2) <= CNStageIntLLROutputS3xD(123)(1);
  VNStageIntLLRInputS3xD(141)(0) <= CNStageIntLLROutputS3xD(123)(2);
  VNStageIntLLRInputS3xD(204)(2) <= CNStageIntLLROutputS3xD(123)(3);
  VNStageIntLLRInputS3xD(294)(2) <= CNStageIntLLROutputS3xD(123)(4);
  VNStageIntLLRInputS3xD(367)(2) <= CNStageIntLLROutputS3xD(123)(5);
  VNStageIntLLRInputS3xD(17)(2) <= CNStageIntLLROutputS3xD(124)(0);
  VNStageIntLLRInputS3xD(76)(2) <= CNStageIntLLROutputS3xD(124)(1);
  VNStageIntLLRInputS3xD(139)(2) <= CNStageIntLLROutputS3xD(124)(2);
  VNStageIntLLRInputS3xD(229)(2) <= CNStageIntLLROutputS3xD(124)(3);
  VNStageIntLLRInputS3xD(302)(2) <= CNStageIntLLROutputS3xD(124)(4);
  VNStageIntLLRInputS3xD(347)(2) <= CNStageIntLLROutputS3xD(124)(5);
  VNStageIntLLRInputS3xD(16)(1) <= CNStageIntLLROutputS3xD(125)(0);
  VNStageIntLLRInputS3xD(74)(2) <= CNStageIntLLROutputS3xD(125)(1);
  VNStageIntLLRInputS3xD(164)(2) <= CNStageIntLLROutputS3xD(125)(2);
  VNStageIntLLRInputS3xD(237)(2) <= CNStageIntLLROutputS3xD(125)(3);
  VNStageIntLLRInputS3xD(282)(2) <= CNStageIntLLROutputS3xD(125)(4);
  VNStageIntLLRInputS3xD(341)(2) <= CNStageIntLLROutputS3xD(125)(5);
  VNStageIntLLRInputS3xD(15)(2) <= CNStageIntLLROutputS3xD(126)(0);
  VNStageIntLLRInputS3xD(99)(2) <= CNStageIntLLROutputS3xD(126)(1);
  VNStageIntLLRInputS3xD(172)(2) <= CNStageIntLLROutputS3xD(126)(2);
  VNStageIntLLRInputS3xD(217)(2) <= CNStageIntLLROutputS3xD(126)(3);
  VNStageIntLLRInputS3xD(276)(2) <= CNStageIntLLROutputS3xD(126)(4);
  VNStageIntLLRInputS3xD(320)(1) <= CNStageIntLLROutputS3xD(126)(5);
  VNStageIntLLRInputS3xD(14)(2) <= CNStageIntLLROutputS3xD(127)(0);
  VNStageIntLLRInputS3xD(107)(1) <= CNStageIntLLROutputS3xD(127)(1);
  VNStageIntLLRInputS3xD(152)(2) <= CNStageIntLLROutputS3xD(127)(2);
  VNStageIntLLRInputS3xD(211)(2) <= CNStageIntLLROutputS3xD(127)(3);
  VNStageIntLLRInputS3xD(256)(2) <= CNStageIntLLROutputS3xD(127)(4);
  VNStageIntLLRInputS3xD(340)(2) <= CNStageIntLLROutputS3xD(127)(5);
  VNStageIntLLRInputS3xD(13)(1) <= CNStageIntLLROutputS3xD(128)(0);
  VNStageIntLLRInputS3xD(87)(2) <= CNStageIntLLROutputS3xD(128)(1);
  VNStageIntLLRInputS3xD(146)(2) <= CNStageIntLLROutputS3xD(128)(2);
  VNStageIntLLRInputS3xD(192)(2) <= CNStageIntLLROutputS3xD(128)(3);
  VNStageIntLLRInputS3xD(275)(2) <= CNStageIntLLROutputS3xD(128)(4);
  VNStageIntLLRInputS3xD(345)(2) <= CNStageIntLLROutputS3xD(128)(5);
  VNStageIntLLRInputS3xD(12)(2) <= CNStageIntLLROutputS3xD(129)(0);
  VNStageIntLLRInputS3xD(81)(2) <= CNStageIntLLROutputS3xD(129)(1);
  VNStageIntLLRInputS3xD(128)(2) <= CNStageIntLLROutputS3xD(129)(2);
  VNStageIntLLRInputS3xD(210)(2) <= CNStageIntLLROutputS3xD(129)(3);
  VNStageIntLLRInputS3xD(280)(2) <= CNStageIntLLROutputS3xD(129)(4);
  VNStageIntLLRInputS3xD(364)(2) <= CNStageIntLLROutputS3xD(129)(5);
  VNStageIntLLRInputS3xD(11)(2) <= CNStageIntLLROutputS3xD(130)(0);
  VNStageIntLLRInputS3xD(64)(2) <= CNStageIntLLROutputS3xD(130)(1);
  VNStageIntLLRInputS3xD(145)(2) <= CNStageIntLLROutputS3xD(130)(2);
  VNStageIntLLRInputS3xD(215)(2) <= CNStageIntLLROutputS3xD(130)(3);
  VNStageIntLLRInputS3xD(299)(1) <= CNStageIntLLROutputS3xD(130)(4);
  VNStageIntLLRInputS3xD(355)(2) <= CNStageIntLLROutputS3xD(130)(5);
  VNStageIntLLRInputS3xD(10)(2) <= CNStageIntLLROutputS3xD(131)(0);
  VNStageIntLLRInputS3xD(80)(2) <= CNStageIntLLROutputS3xD(131)(1);
  VNStageIntLLRInputS3xD(150)(2) <= CNStageIntLLROutputS3xD(131)(2);
  VNStageIntLLRInputS3xD(234)(2) <= CNStageIntLLROutputS3xD(131)(3);
  VNStageIntLLRInputS3xD(290)(2) <= CNStageIntLLROutputS3xD(131)(4);
  VNStageIntLLRInputS3xD(329)(2) <= CNStageIntLLROutputS3xD(131)(5);
  VNStageIntLLRInputS3xD(9)(2) <= CNStageIntLLROutputS3xD(132)(0);
  VNStageIntLLRInputS3xD(85)(1) <= CNStageIntLLROutputS3xD(132)(1);
  VNStageIntLLRInputS3xD(169)(2) <= CNStageIntLLROutputS3xD(132)(2);
  VNStageIntLLRInputS3xD(225)(2) <= CNStageIntLLROutputS3xD(132)(3);
  VNStageIntLLRInputS3xD(264)(2) <= CNStageIntLLROutputS3xD(132)(4);
  VNStageIntLLRInputS3xD(330)(2) <= CNStageIntLLROutputS3xD(132)(5);
  VNStageIntLLRInputS3xD(8)(1) <= CNStageIntLLROutputS3xD(133)(0);
  VNStageIntLLRInputS3xD(104)(2) <= CNStageIntLLROutputS3xD(133)(1);
  VNStageIntLLRInputS3xD(160)(2) <= CNStageIntLLROutputS3xD(133)(2);
  VNStageIntLLRInputS3xD(199)(2) <= CNStageIntLLROutputS3xD(133)(3);
  VNStageIntLLRInputS3xD(265)(1) <= CNStageIntLLROutputS3xD(133)(4);
  VNStageIntLLRInputS3xD(354)(2) <= CNStageIntLLROutputS3xD(133)(5);
  VNStageIntLLRInputS3xD(7)(2) <= CNStageIntLLROutputS3xD(134)(0);
  VNStageIntLLRInputS3xD(95)(2) <= CNStageIntLLROutputS3xD(134)(1);
  VNStageIntLLRInputS3xD(134)(2) <= CNStageIntLLROutputS3xD(134)(2);
  VNStageIntLLRInputS3xD(200)(2) <= CNStageIntLLROutputS3xD(134)(3);
  VNStageIntLLRInputS3xD(289)(2) <= CNStageIntLLROutputS3xD(134)(4);
  VNStageIntLLRInputS3xD(375)(2) <= CNStageIntLLROutputS3xD(134)(5);
  VNStageIntLLRInputS3xD(6)(2) <= CNStageIntLLROutputS3xD(135)(0);
  VNStageIntLLRInputS3xD(69)(2) <= CNStageIntLLROutputS3xD(135)(1);
  VNStageIntLLRInputS3xD(135)(2) <= CNStageIntLLROutputS3xD(135)(2);
  VNStageIntLLRInputS3xD(224)(2) <= CNStageIntLLROutputS3xD(135)(3);
  VNStageIntLLRInputS3xD(310)(2) <= CNStageIntLLROutputS3xD(135)(4);
  VNStageIntLLRInputS3xD(371)(1) <= CNStageIntLLROutputS3xD(135)(5);
  VNStageIntLLRInputS3xD(5)(2) <= CNStageIntLLROutputS3xD(136)(0);
  VNStageIntLLRInputS3xD(70)(2) <= CNStageIntLLROutputS3xD(136)(1);
  VNStageIntLLRInputS3xD(159)(2) <= CNStageIntLLROutputS3xD(136)(2);
  VNStageIntLLRInputS3xD(245)(2) <= CNStageIntLLROutputS3xD(136)(3);
  VNStageIntLLRInputS3xD(306)(2) <= CNStageIntLLROutputS3xD(136)(4);
  VNStageIntLLRInputS3xD(323)(1) <= CNStageIntLLROutputS3xD(136)(5);
  VNStageIntLLRInputS3xD(3)(1) <= CNStageIntLLROutputS3xD(137)(0);
  VNStageIntLLRInputS3xD(115)(2) <= CNStageIntLLROutputS3xD(137)(1);
  VNStageIntLLRInputS3xD(176)(2) <= CNStageIntLLROutputS3xD(137)(2);
  VNStageIntLLRInputS3xD(193)(2) <= CNStageIntLLROutputS3xD(137)(3);
  VNStageIntLLRInputS3xD(284)(2) <= CNStageIntLLROutputS3xD(137)(4);
  VNStageIntLLRInputS3xD(325)(2) <= CNStageIntLLROutputS3xD(137)(5);
  VNStageIntLLRInputS3xD(2)(2) <= CNStageIntLLROutputS3xD(138)(0);
  VNStageIntLLRInputS3xD(111)(2) <= CNStageIntLLROutputS3xD(138)(1);
  VNStageIntLLRInputS3xD(191)(2) <= CNStageIntLLROutputS3xD(138)(2);
  VNStageIntLLRInputS3xD(219)(2) <= CNStageIntLLROutputS3xD(138)(3);
  VNStageIntLLRInputS3xD(260)(2) <= CNStageIntLLROutputS3xD(138)(4);
  VNStageIntLLRInputS3xD(357)(2) <= CNStageIntLLROutputS3xD(138)(5);
  VNStageIntLLRInputS3xD(1)(1) <= CNStageIntLLROutputS3xD(139)(0);
  VNStageIntLLRInputS3xD(126)(1) <= CNStageIntLLROutputS3xD(139)(1);
  VNStageIntLLRInputS3xD(154)(1) <= CNStageIntLLROutputS3xD(139)(2);
  VNStageIntLLRInputS3xD(195)(1) <= CNStageIntLLROutputS3xD(139)(3);
  VNStageIntLLRInputS3xD(292)(2) <= CNStageIntLLROutputS3xD(139)(4);
  VNStageIntLLRInputS3xD(373)(1) <= CNStageIntLLROutputS3xD(139)(5);
  VNStageIntLLRInputS3xD(63)(2) <= CNStageIntLLROutputS3xD(140)(0);
  VNStageIntLLRInputS3xD(89)(2) <= CNStageIntLLROutputS3xD(140)(1);
  VNStageIntLLRInputS3xD(130)(2) <= CNStageIntLLROutputS3xD(140)(2);
  VNStageIntLLRInputS3xD(227)(2) <= CNStageIntLLROutputS3xD(140)(3);
  VNStageIntLLRInputS3xD(308)(0) <= CNStageIntLLROutputS3xD(140)(4);
  VNStageIntLLRInputS3xD(343)(2) <= CNStageIntLLROutputS3xD(140)(5);
  VNStageIntLLRInputS3xD(62)(1) <= CNStageIntLLROutputS3xD(141)(0);
  VNStageIntLLRInputS3xD(65)(2) <= CNStageIntLLROutputS3xD(141)(1);
  VNStageIntLLRInputS3xD(162)(2) <= CNStageIntLLROutputS3xD(141)(2);
  VNStageIntLLRInputS3xD(243)(2) <= CNStageIntLLROutputS3xD(141)(3);
  VNStageIntLLRInputS3xD(278)(2) <= CNStageIntLLROutputS3xD(141)(4);
  VNStageIntLLRInputS3xD(352)(2) <= CNStageIntLLROutputS3xD(141)(5);
  VNStageIntLLRInputS3xD(61)(1) <= CNStageIntLLROutputS3xD(142)(0);
  VNStageIntLLRInputS3xD(97)(2) <= CNStageIntLLROutputS3xD(142)(1);
  VNStageIntLLRInputS3xD(178)(2) <= CNStageIntLLROutputS3xD(142)(2);
  VNStageIntLLRInputS3xD(213)(2) <= CNStageIntLLROutputS3xD(142)(3);
  VNStageIntLLRInputS3xD(287)(2) <= CNStageIntLLROutputS3xD(142)(4);
  VNStageIntLLRInputS3xD(365)(2) <= CNStageIntLLROutputS3xD(142)(5);
  VNStageIntLLRInputS3xD(60)(1) <= CNStageIntLLROutputS3xD(143)(0);
  VNStageIntLLRInputS3xD(113)(2) <= CNStageIntLLROutputS3xD(143)(1);
  VNStageIntLLRInputS3xD(148)(2) <= CNStageIntLLROutputS3xD(143)(2);
  VNStageIntLLRInputS3xD(222)(1) <= CNStageIntLLROutputS3xD(143)(3);
  VNStageIntLLRInputS3xD(300)(2) <= CNStageIntLLROutputS3xD(143)(4);
  VNStageIntLLRInputS3xD(344)(2) <= CNStageIntLLROutputS3xD(143)(5);
  VNStageIntLLRInputS3xD(59)(0) <= CNStageIntLLROutputS3xD(144)(0);
  VNStageIntLLRInputS3xD(83)(2) <= CNStageIntLLROutputS3xD(144)(1);
  VNStageIntLLRInputS3xD(157)(2) <= CNStageIntLLROutputS3xD(144)(2);
  VNStageIntLLRInputS3xD(235)(1) <= CNStageIntLLROutputS3xD(144)(3);
  VNStageIntLLRInputS3xD(279)(2) <= CNStageIntLLROutputS3xD(144)(4);
  VNStageIntLLRInputS3xD(372)(1) <= CNStageIntLLROutputS3xD(144)(5);
  VNStageIntLLRInputS3xD(58)(1) <= CNStageIntLLROutputS3xD(145)(0);
  VNStageIntLLRInputS3xD(92)(2) <= CNStageIntLLROutputS3xD(145)(1);
  VNStageIntLLRInputS3xD(170)(2) <= CNStageIntLLROutputS3xD(145)(2);
  VNStageIntLLRInputS3xD(214)(2) <= CNStageIntLLROutputS3xD(145)(3);
  VNStageIntLLRInputS3xD(307)(2) <= CNStageIntLLROutputS3xD(145)(4);
  VNStageIntLLRInputS3xD(374)(2) <= CNStageIntLLROutputS3xD(145)(5);
  VNStageIntLLRInputS3xD(57)(1) <= CNStageIntLLROutputS3xD(146)(0);
  VNStageIntLLRInputS3xD(105)(1) <= CNStageIntLLROutputS3xD(146)(1);
  VNStageIntLLRInputS3xD(149)(2) <= CNStageIntLLROutputS3xD(146)(2);
  VNStageIntLLRInputS3xD(242)(2) <= CNStageIntLLROutputS3xD(146)(3);
  VNStageIntLLRInputS3xD(309)(2) <= CNStageIntLLROutputS3xD(146)(4);
  VNStageIntLLRInputS3xD(356)(2) <= CNStageIntLLROutputS3xD(146)(5);
  VNStageIntLLRInputS3xD(56)(2) <= CNStageIntLLROutputS3xD(147)(0);
  VNStageIntLLRInputS3xD(84)(2) <= CNStageIntLLROutputS3xD(147)(1);
  VNStageIntLLRInputS3xD(177)(2) <= CNStageIntLLROutputS3xD(147)(2);
  VNStageIntLLRInputS3xD(244)(0) <= CNStageIntLLROutputS3xD(147)(3);
  VNStageIntLLRInputS3xD(291)(2) <= CNStageIntLLROutputS3xD(147)(4);
  VNStageIntLLRInputS3xD(363)(1) <= CNStageIntLLROutputS3xD(147)(5);
  VNStageIntLLRInputS3xD(55)(2) <= CNStageIntLLROutputS3xD(148)(0);
  VNStageIntLLRInputS3xD(112)(2) <= CNStageIntLLROutputS3xD(148)(1);
  VNStageIntLLRInputS3xD(179)(2) <= CNStageIntLLROutputS3xD(148)(2);
  VNStageIntLLRInputS3xD(226)(1) <= CNStageIntLLROutputS3xD(148)(3);
  VNStageIntLLRInputS3xD(298)(2) <= CNStageIntLLROutputS3xD(148)(4);
  VNStageIntLLRInputS3xD(327)(2) <= CNStageIntLLROutputS3xD(148)(5);
  VNStageIntLLRInputS3xD(54)(2) <= CNStageIntLLROutputS3xD(149)(0);
  VNStageIntLLRInputS3xD(114)(2) <= CNStageIntLLROutputS3xD(149)(1);
  VNStageIntLLRInputS3xD(161)(2) <= CNStageIntLLROutputS3xD(149)(2);
  VNStageIntLLRInputS3xD(233)(2) <= CNStageIntLLROutputS3xD(149)(3);
  VNStageIntLLRInputS3xD(262)(2) <= CNStageIntLLROutputS3xD(149)(4);
  VNStageIntLLRInputS3xD(378)(1) <= CNStageIntLLROutputS3xD(149)(5);
  VNStageIntLLRInputS3xD(53)(1) <= CNStageIntLLROutputS3xD(150)(0);
  VNStageIntLLRInputS3xD(96)(2) <= CNStageIntLLROutputS3xD(150)(1);
  VNStageIntLLRInputS3xD(168)(1) <= CNStageIntLLROutputS3xD(150)(2);
  VNStageIntLLRInputS3xD(197)(2) <= CNStageIntLLROutputS3xD(150)(3);
  VNStageIntLLRInputS3xD(313)(0) <= CNStageIntLLROutputS3xD(150)(4);
  VNStageIntLLRInputS3xD(321)(2) <= CNStageIntLLROutputS3xD(150)(5);
  VNStageIntLLRInputS3xD(52)(1) <= CNStageIntLLROutputS3xD(151)(0);
  VNStageIntLLRInputS3xD(103)(2) <= CNStageIntLLROutputS3xD(151)(1);
  VNStageIntLLRInputS3xD(132)(1) <= CNStageIntLLROutputS3xD(151)(2);
  VNStageIntLLRInputS3xD(248)(2) <= CNStageIntLLROutputS3xD(151)(3);
  VNStageIntLLRInputS3xD(319)(2) <= CNStageIntLLROutputS3xD(151)(4);
  VNStageIntLLRInputS3xD(379)(1) <= CNStageIntLLROutputS3xD(151)(5);
  VNStageIntLLRInputS3xD(50)(2) <= CNStageIntLLROutputS3xD(152)(0);
  VNStageIntLLRInputS3xD(118)(2) <= CNStageIntLLROutputS3xD(152)(1);
  VNStageIntLLRInputS3xD(189)(1) <= CNStageIntLLROutputS3xD(152)(2);
  VNStageIntLLRInputS3xD(249)(0) <= CNStageIntLLROutputS3xD(152)(3);
  VNStageIntLLRInputS3xD(261)(2) <= CNStageIntLLROutputS3xD(152)(4);
  VNStageIntLLRInputS3xD(348)(2) <= CNStageIntLLROutputS3xD(152)(5);
  VNStageIntLLRInputS3xD(49)(2) <= CNStageIntLLROutputS3xD(153)(0);
  VNStageIntLLRInputS3xD(124)(1) <= CNStageIntLLROutputS3xD(153)(1);
  VNStageIntLLRInputS3xD(184)(2) <= CNStageIntLLROutputS3xD(153)(2);
  VNStageIntLLRInputS3xD(196)(2) <= CNStageIntLLROutputS3xD(153)(3);
  VNStageIntLLRInputS3xD(283)(2) <= CNStageIntLLROutputS3xD(153)(4);
  VNStageIntLLRInputS3xD(366)(2) <= CNStageIntLLROutputS3xD(153)(5);
  VNStageIntLLRInputS3xD(48)(1) <= CNStageIntLLROutputS3xD(154)(0);
  VNStageIntLLRInputS3xD(119)(2) <= CNStageIntLLROutputS3xD(154)(1);
  VNStageIntLLRInputS3xD(131)(1) <= CNStageIntLLROutputS3xD(154)(2);
  VNStageIntLLRInputS3xD(218)(2) <= CNStageIntLLROutputS3xD(154)(3);
  VNStageIntLLRInputS3xD(301)(2) <= CNStageIntLLROutputS3xD(154)(4);
  VNStageIntLLRInputS3xD(351)(1) <= CNStageIntLLROutputS3xD(154)(5);
  VNStageIntLLRInputS3xD(47)(1) <= CNStageIntLLROutputS3xD(155)(0);
  VNStageIntLLRInputS3xD(66)(2) <= CNStageIntLLROutputS3xD(155)(1);
  VNStageIntLLRInputS3xD(153)(2) <= CNStageIntLLROutputS3xD(155)(2);
  VNStageIntLLRInputS3xD(236)(2) <= CNStageIntLLROutputS3xD(155)(3);
  VNStageIntLLRInputS3xD(286)(2) <= CNStageIntLLROutputS3xD(155)(4);
  VNStageIntLLRInputS3xD(338)(2) <= CNStageIntLLROutputS3xD(155)(5);
  VNStageIntLLRInputS3xD(46)(2) <= CNStageIntLLROutputS3xD(156)(0);
  VNStageIntLLRInputS3xD(88)(2) <= CNStageIntLLROutputS3xD(156)(1);
  VNStageIntLLRInputS3xD(171)(1) <= CNStageIntLLROutputS3xD(156)(2);
  VNStageIntLLRInputS3xD(221)(2) <= CNStageIntLLROutputS3xD(156)(3);
  VNStageIntLLRInputS3xD(273)(2) <= CNStageIntLLROutputS3xD(156)(4);
  VNStageIntLLRInputS3xD(369)(1) <= CNStageIntLLROutputS3xD(156)(5);
  VNStageIntLLRInputS3xD(45)(2) <= CNStageIntLLROutputS3xD(157)(0);
  VNStageIntLLRInputS3xD(106)(1) <= CNStageIntLLROutputS3xD(157)(1);
  VNStageIntLLRInputS3xD(156)(2) <= CNStageIntLLROutputS3xD(157)(2);
  VNStageIntLLRInputS3xD(208)(2) <= CNStageIntLLROutputS3xD(157)(3);
  VNStageIntLLRInputS3xD(304)(2) <= CNStageIntLLROutputS3xD(157)(4);
  VNStageIntLLRInputS3xD(381)(1) <= CNStageIntLLROutputS3xD(157)(5);
  VNStageIntLLRInputS3xD(44)(2) <= CNStageIntLLROutputS3xD(158)(0);
  VNStageIntLLRInputS3xD(91)(2) <= CNStageIntLLROutputS3xD(158)(1);
  VNStageIntLLRInputS3xD(143)(2) <= CNStageIntLLROutputS3xD(158)(2);
  VNStageIntLLRInputS3xD(239)(2) <= CNStageIntLLROutputS3xD(158)(3);
  VNStageIntLLRInputS3xD(316)(1) <= CNStageIntLLROutputS3xD(158)(4);
  VNStageIntLLRInputS3xD(332)(2) <= CNStageIntLLROutputS3xD(158)(5);
  VNStageIntLLRInputS3xD(43)(1) <= CNStageIntLLROutputS3xD(159)(0);
  VNStageIntLLRInputS3xD(78)(2) <= CNStageIntLLROutputS3xD(159)(1);
  VNStageIntLLRInputS3xD(174)(2) <= CNStageIntLLROutputS3xD(159)(2);
  VNStageIntLLRInputS3xD(251)(1) <= CNStageIntLLROutputS3xD(159)(3);
  VNStageIntLLRInputS3xD(267)(2) <= CNStageIntLLROutputS3xD(159)(4);
  VNStageIntLLRInputS3xD(376)(2) <= CNStageIntLLROutputS3xD(159)(5);
  VNStageIntLLRInputS3xD(42)(2) <= CNStageIntLLROutputS3xD(160)(0);
  VNStageIntLLRInputS3xD(109)(2) <= CNStageIntLLROutputS3xD(160)(1);
  VNStageIntLLRInputS3xD(186)(1) <= CNStageIntLLROutputS3xD(160)(2);
  VNStageIntLLRInputS3xD(202)(2) <= CNStageIntLLROutputS3xD(160)(3);
  VNStageIntLLRInputS3xD(311)(2) <= CNStageIntLLROutputS3xD(160)(4);
  VNStageIntLLRInputS3xD(353)(2) <= CNStageIntLLROutputS3xD(160)(5);
  VNStageIntLLRInputS3xD(41)(2) <= CNStageIntLLROutputS3xD(161)(0);
  VNStageIntLLRInputS3xD(121)(1) <= CNStageIntLLROutputS3xD(161)(1);
  VNStageIntLLRInputS3xD(137)(2) <= CNStageIntLLROutputS3xD(161)(2);
  VNStageIntLLRInputS3xD(246)(2) <= CNStageIntLLROutputS3xD(161)(3);
  VNStageIntLLRInputS3xD(288)(2) <= CNStageIntLLROutputS3xD(161)(4);
  VNStageIntLLRInputS3xD(342)(2) <= CNStageIntLLROutputS3xD(161)(5);
  VNStageIntLLRInputS3xD(40)(2) <= CNStageIntLLROutputS3xD(162)(0);
  VNStageIntLLRInputS3xD(72)(2) <= CNStageIntLLROutputS3xD(162)(1);
  VNStageIntLLRInputS3xD(181)(2) <= CNStageIntLLROutputS3xD(162)(2);
  VNStageIntLLRInputS3xD(223)(2) <= CNStageIntLLROutputS3xD(162)(3);
  VNStageIntLLRInputS3xD(277)(2) <= CNStageIntLLROutputS3xD(162)(4);
  VNStageIntLLRInputS3xD(346)(2) <= CNStageIntLLROutputS3xD(162)(5);
  VNStageIntLLRInputS3xD(39)(2) <= CNStageIntLLROutputS3xD(163)(0);
  VNStageIntLLRInputS3xD(116)(1) <= CNStageIntLLROutputS3xD(163)(1);
  VNStageIntLLRInputS3xD(158)(2) <= CNStageIntLLROutputS3xD(163)(2);
  VNStageIntLLRInputS3xD(212)(2) <= CNStageIntLLROutputS3xD(163)(3);
  VNStageIntLLRInputS3xD(281)(2) <= CNStageIntLLROutputS3xD(163)(4);
  VNStageIntLLRInputS3xD(339)(2) <= CNStageIntLLROutputS3xD(163)(5);
  VNStageIntLLRInputS3xD(38)(2) <= CNStageIntLLROutputS3xD(164)(0);
  VNStageIntLLRInputS3xD(93)(2) <= CNStageIntLLROutputS3xD(164)(1);
  VNStageIntLLRInputS3xD(147)(2) <= CNStageIntLLROutputS3xD(164)(2);
  VNStageIntLLRInputS3xD(216)(2) <= CNStageIntLLROutputS3xD(164)(3);
  VNStageIntLLRInputS3xD(274)(1) <= CNStageIntLLROutputS3xD(164)(4);
  VNStageIntLLRInputS3xD(350)(2) <= CNStageIntLLROutputS3xD(164)(5);
  VNStageIntLLRInputS3xD(37)(2) <= CNStageIntLLROutputS3xD(165)(0);
  VNStageIntLLRInputS3xD(82)(2) <= CNStageIntLLROutputS3xD(165)(1);
  VNStageIntLLRInputS3xD(151)(2) <= CNStageIntLLROutputS3xD(165)(2);
  VNStageIntLLRInputS3xD(209)(2) <= CNStageIntLLROutputS3xD(165)(3);
  VNStageIntLLRInputS3xD(285)(2) <= CNStageIntLLROutputS3xD(165)(4);
  VNStageIntLLRInputS3xD(322)(2) <= CNStageIntLLROutputS3xD(165)(5);
  VNStageIntLLRInputS3xD(36)(2) <= CNStageIntLLROutputS3xD(166)(0);
  VNStageIntLLRInputS3xD(86)(1) <= CNStageIntLLROutputS3xD(166)(1);
  VNStageIntLLRInputS3xD(144)(2) <= CNStageIntLLROutputS3xD(166)(2);
  VNStageIntLLRInputS3xD(220)(2) <= CNStageIntLLROutputS3xD(166)(3);
  VNStageIntLLRInputS3xD(257)(2) <= CNStageIntLLROutputS3xD(166)(4);
  VNStageIntLLRInputS3xD(377)(1) <= CNStageIntLLROutputS3xD(166)(5);
  VNStageIntLLRInputS3xD(35)(2) <= CNStageIntLLROutputS3xD(167)(0);
  VNStageIntLLRInputS3xD(79)(2) <= CNStageIntLLROutputS3xD(167)(1);
  VNStageIntLLRInputS3xD(155)(2) <= CNStageIntLLROutputS3xD(167)(2);
  VNStageIntLLRInputS3xD(255)(2) <= CNStageIntLLROutputS3xD(167)(3);
  VNStageIntLLRInputS3xD(312)(2) <= CNStageIntLLROutputS3xD(167)(4);
  VNStageIntLLRInputS3xD(331)(2) <= CNStageIntLLROutputS3xD(167)(5);
  VNStageIntLLRInputS3xD(34)(2) <= CNStageIntLLROutputS3xD(168)(0);
  VNStageIntLLRInputS3xD(90)(2) <= CNStageIntLLROutputS3xD(168)(1);
  VNStageIntLLRInputS3xD(190)(0) <= CNStageIntLLROutputS3xD(168)(2);
  VNStageIntLLRInputS3xD(247)(2) <= CNStageIntLLROutputS3xD(168)(3);
  VNStageIntLLRInputS3xD(266)(1) <= CNStageIntLLROutputS3xD(168)(4);
  VNStageIntLLRInputS3xD(328)(2) <= CNStageIntLLROutputS3xD(168)(5);
  VNStageIntLLRInputS3xD(33)(2) <= CNStageIntLLROutputS3xD(169)(0);
  VNStageIntLLRInputS3xD(125)(1) <= CNStageIntLLROutputS3xD(169)(1);
  VNStageIntLLRInputS3xD(182)(2) <= CNStageIntLLROutputS3xD(169)(2);
  VNStageIntLLRInputS3xD(201)(2) <= CNStageIntLLROutputS3xD(169)(3);
  VNStageIntLLRInputS3xD(263)(2) <= CNStageIntLLROutputS3xD(169)(4);
  VNStageIntLLRInputS3xD(362)(2) <= CNStageIntLLROutputS3xD(169)(5);
  VNStageIntLLRInputS3xD(0)(2) <= CNStageIntLLROutputS3xD(170)(0);
  VNStageIntLLRInputS3xD(75)(2) <= CNStageIntLLROutputS3xD(170)(1);
  VNStageIntLLRInputS3xD(140)(2) <= CNStageIntLLROutputS3xD(170)(2);
  VNStageIntLLRInputS3xD(205)(0) <= CNStageIntLLROutputS3xD(170)(3);
  VNStageIntLLRInputS3xD(270)(2) <= CNStageIntLLROutputS3xD(170)(4);
  VNStageIntLLRInputS3xD(335)(2) <= CNStageIntLLROutputS3xD(170)(5);
  VNStageIntLLRInputS3xD(62)(2) <= CNStageIntLLROutputS3xD(171)(0);
  VNStageIntLLRInputS3xD(109)(3) <= CNStageIntLLROutputS3xD(171)(1);
  VNStageIntLLRInputS3xD(161)(3) <= CNStageIntLLROutputS3xD(171)(2);
  VNStageIntLLRInputS3xD(194)(3) <= CNStageIntLLROutputS3xD(171)(3);
  VNStageIntLLRInputS3xD(271)(2) <= CNStageIntLLROutputS3xD(171)(4);
  VNStageIntLLRInputS3xD(350)(3) <= CNStageIntLLROutputS3xD(171)(5);
  VNStageIntLLRInputS3xD(61)(2) <= CNStageIntLLROutputS3xD(172)(0);
  VNStageIntLLRInputS3xD(96)(3) <= CNStageIntLLROutputS3xD(172)(1);
  VNStageIntLLRInputS3xD(129)(3) <= CNStageIntLLROutputS3xD(172)(2);
  VNStageIntLLRInputS3xD(206)(2) <= CNStageIntLLROutputS3xD(172)(3);
  VNStageIntLLRInputS3xD(285)(3) <= CNStageIntLLROutputS3xD(172)(4);
  VNStageIntLLRInputS3xD(331)(3) <= CNStageIntLLROutputS3xD(172)(5);
  VNStageIntLLRInputS3xD(60)(2) <= CNStageIntLLROutputS3xD(173)(0);
  VNStageIntLLRInputS3xD(127)(3) <= CNStageIntLLROutputS3xD(173)(1);
  VNStageIntLLRInputS3xD(141)(1) <= CNStageIntLLROutputS3xD(173)(2);
  VNStageIntLLRInputS3xD(220)(3) <= CNStageIntLLROutputS3xD(173)(3);
  VNStageIntLLRInputS3xD(266)(2) <= CNStageIntLLROutputS3xD(173)(4);
  VNStageIntLLRInputS3xD(371)(2) <= CNStageIntLLROutputS3xD(173)(5);
  VNStageIntLLRInputS3xD(59)(1) <= CNStageIntLLROutputS3xD(174)(0);
  VNStageIntLLRInputS3xD(76)(3) <= CNStageIntLLROutputS3xD(174)(1);
  VNStageIntLLRInputS3xD(155)(3) <= CNStageIntLLROutputS3xD(174)(2);
  VNStageIntLLRInputS3xD(201)(3) <= CNStageIntLLROutputS3xD(174)(3);
  VNStageIntLLRInputS3xD(306)(3) <= CNStageIntLLROutputS3xD(174)(4);
  VNStageIntLLRInputS3xD(360)(3) <= CNStageIntLLROutputS3xD(174)(5);
  VNStageIntLLRInputS3xD(58)(2) <= CNStageIntLLROutputS3xD(175)(0);
  VNStageIntLLRInputS3xD(90)(3) <= CNStageIntLLROutputS3xD(175)(1);
  VNStageIntLLRInputS3xD(136)(3) <= CNStageIntLLROutputS3xD(175)(2);
  VNStageIntLLRInputS3xD(241)(2) <= CNStageIntLLROutputS3xD(175)(3);
  VNStageIntLLRInputS3xD(295)(3) <= CNStageIntLLROutputS3xD(175)(4);
  VNStageIntLLRInputS3xD(364)(3) <= CNStageIntLLROutputS3xD(175)(5);
  VNStageIntLLRInputS3xD(57)(2) <= CNStageIntLLROutputS3xD(176)(0);
  VNStageIntLLRInputS3xD(71)(2) <= CNStageIntLLROutputS3xD(176)(1);
  VNStageIntLLRInputS3xD(176)(3) <= CNStageIntLLROutputS3xD(176)(2);
  VNStageIntLLRInputS3xD(230)(2) <= CNStageIntLLROutputS3xD(176)(3);
  VNStageIntLLRInputS3xD(299)(2) <= CNStageIntLLROutputS3xD(176)(4);
  VNStageIntLLRInputS3xD(357)(3) <= CNStageIntLLROutputS3xD(176)(5);
  VNStageIntLLRInputS3xD(56)(3) <= CNStageIntLLROutputS3xD(177)(0);
  VNStageIntLLRInputS3xD(111)(3) <= CNStageIntLLROutputS3xD(177)(1);
  VNStageIntLLRInputS3xD(165)(3) <= CNStageIntLLROutputS3xD(177)(2);
  VNStageIntLLRInputS3xD(234)(3) <= CNStageIntLLROutputS3xD(177)(3);
  VNStageIntLLRInputS3xD(292)(3) <= CNStageIntLLROutputS3xD(177)(4);
  VNStageIntLLRInputS3xD(368)(1) <= CNStageIntLLROutputS3xD(177)(5);
  VNStageIntLLRInputS3xD(55)(3) <= CNStageIntLLROutputS3xD(178)(0);
  VNStageIntLLRInputS3xD(100)(3) <= CNStageIntLLROutputS3xD(178)(1);
  VNStageIntLLRInputS3xD(169)(3) <= CNStageIntLLROutputS3xD(178)(2);
  VNStageIntLLRInputS3xD(227)(3) <= CNStageIntLLROutputS3xD(178)(3);
  VNStageIntLLRInputS3xD(303)(3) <= CNStageIntLLROutputS3xD(178)(4);
  VNStageIntLLRInputS3xD(340)(3) <= CNStageIntLLROutputS3xD(178)(5);
  VNStageIntLLRInputS3xD(54)(3) <= CNStageIntLLROutputS3xD(179)(0);
  VNStageIntLLRInputS3xD(104)(3) <= CNStageIntLLROutputS3xD(179)(1);
  VNStageIntLLRInputS3xD(162)(3) <= CNStageIntLLROutputS3xD(179)(2);
  VNStageIntLLRInputS3xD(238)(3) <= CNStageIntLLROutputS3xD(179)(3);
  VNStageIntLLRInputS3xD(275)(3) <= CNStageIntLLROutputS3xD(179)(4);
  VNStageIntLLRInputS3xD(332)(3) <= CNStageIntLLROutputS3xD(179)(5);
  VNStageIntLLRInputS3xD(53)(2) <= CNStageIntLLROutputS3xD(180)(0);
  VNStageIntLLRInputS3xD(97)(3) <= CNStageIntLLROutputS3xD(180)(1);
  VNStageIntLLRInputS3xD(173)(3) <= CNStageIntLLROutputS3xD(180)(2);
  VNStageIntLLRInputS3xD(210)(3) <= CNStageIntLLROutputS3xD(180)(3);
  VNStageIntLLRInputS3xD(267)(3) <= CNStageIntLLROutputS3xD(180)(4);
  VNStageIntLLRInputS3xD(349)(2) <= CNStageIntLLROutputS3xD(180)(5);
  VNStageIntLLRInputS3xD(52)(2) <= CNStageIntLLROutputS3xD(181)(0);
  VNStageIntLLRInputS3xD(108)(3) <= CNStageIntLLROutputS3xD(181)(1);
  VNStageIntLLRInputS3xD(145)(3) <= CNStageIntLLROutputS3xD(181)(2);
  VNStageIntLLRInputS3xD(202)(3) <= CNStageIntLLROutputS3xD(181)(3);
  VNStageIntLLRInputS3xD(284)(3) <= CNStageIntLLROutputS3xD(181)(4);
  VNStageIntLLRInputS3xD(346)(3) <= CNStageIntLLROutputS3xD(181)(5);
  VNStageIntLLRInputS3xD(51)(2) <= CNStageIntLLROutputS3xD(182)(0);
  VNStageIntLLRInputS3xD(80)(3) <= CNStageIntLLROutputS3xD(182)(1);
  VNStageIntLLRInputS3xD(137)(3) <= CNStageIntLLROutputS3xD(182)(2);
  VNStageIntLLRInputS3xD(219)(3) <= CNStageIntLLROutputS3xD(182)(3);
  VNStageIntLLRInputS3xD(281)(3) <= CNStageIntLLROutputS3xD(182)(4);
  VNStageIntLLRInputS3xD(380)(2) <= CNStageIntLLROutputS3xD(182)(5);
  VNStageIntLLRInputS3xD(50)(3) <= CNStageIntLLROutputS3xD(183)(0);
  VNStageIntLLRInputS3xD(72)(3) <= CNStageIntLLROutputS3xD(183)(1);
  VNStageIntLLRInputS3xD(154)(2) <= CNStageIntLLROutputS3xD(183)(2);
  VNStageIntLLRInputS3xD(216)(3) <= CNStageIntLLROutputS3xD(183)(3);
  VNStageIntLLRInputS3xD(315)(2) <= CNStageIntLLROutputS3xD(183)(4);
  VNStageIntLLRInputS3xD(337)(3) <= CNStageIntLLROutputS3xD(183)(5);
  VNStageIntLLRInputS3xD(49)(3) <= CNStageIntLLROutputS3xD(184)(0);
  VNStageIntLLRInputS3xD(89)(3) <= CNStageIntLLROutputS3xD(184)(1);
  VNStageIntLLRInputS3xD(151)(3) <= CNStageIntLLROutputS3xD(184)(2);
  VNStageIntLLRInputS3xD(250)(2) <= CNStageIntLLROutputS3xD(184)(3);
  VNStageIntLLRInputS3xD(272)(3) <= CNStageIntLLROutputS3xD(184)(4);
  VNStageIntLLRInputS3xD(323)(2) <= CNStageIntLLROutputS3xD(184)(5);
  VNStageIntLLRInputS3xD(46)(3) <= CNStageIntLLROutputS3xD(185)(0);
  VNStageIntLLRInputS3xD(77)(1) <= CNStageIntLLROutputS3xD(185)(1);
  VNStageIntLLRInputS3xD(191)(3) <= CNStageIntLLROutputS3xD(185)(2);
  VNStageIntLLRInputS3xD(246)(3) <= CNStageIntLLROutputS3xD(185)(3);
  VNStageIntLLRInputS3xD(277)(3) <= CNStageIntLLROutputS3xD(185)(4);
  VNStageIntLLRInputS3xD(325)(3) <= CNStageIntLLROutputS3xD(185)(5);
  VNStageIntLLRInputS3xD(45)(3) <= CNStageIntLLROutputS3xD(186)(0);
  VNStageIntLLRInputS3xD(126)(2) <= CNStageIntLLROutputS3xD(186)(1);
  VNStageIntLLRInputS3xD(181)(3) <= CNStageIntLLROutputS3xD(186)(2);
  VNStageIntLLRInputS3xD(212)(3) <= CNStageIntLLROutputS3xD(186)(3);
  VNStageIntLLRInputS3xD(260)(3) <= CNStageIntLLROutputS3xD(186)(4);
  VNStageIntLLRInputS3xD(355)(3) <= CNStageIntLLROutputS3xD(186)(5);
  VNStageIntLLRInputS3xD(44)(3) <= CNStageIntLLROutputS3xD(187)(0);
  VNStageIntLLRInputS3xD(116)(2) <= CNStageIntLLROutputS3xD(187)(1);
  VNStageIntLLRInputS3xD(147)(3) <= CNStageIntLLROutputS3xD(187)(2);
  VNStageIntLLRInputS3xD(195)(2) <= CNStageIntLLROutputS3xD(187)(3);
  VNStageIntLLRInputS3xD(290)(3) <= CNStageIntLLROutputS3xD(187)(4);
  VNStageIntLLRInputS3xD(378)(2) <= CNStageIntLLROutputS3xD(187)(5);
  VNStageIntLLRInputS3xD(43)(2) <= CNStageIntLLROutputS3xD(188)(0);
  VNStageIntLLRInputS3xD(82)(3) <= CNStageIntLLROutputS3xD(188)(1);
  VNStageIntLLRInputS3xD(130)(3) <= CNStageIntLLROutputS3xD(188)(2);
  VNStageIntLLRInputS3xD(225)(3) <= CNStageIntLLROutputS3xD(188)(3);
  VNStageIntLLRInputS3xD(313)(1) <= CNStageIntLLROutputS3xD(188)(4);
  VNStageIntLLRInputS3xD(351)(2) <= CNStageIntLLROutputS3xD(188)(5);
  VNStageIntLLRInputS3xD(42)(3) <= CNStageIntLLROutputS3xD(189)(0);
  VNStageIntLLRInputS3xD(65)(3) <= CNStageIntLLROutputS3xD(189)(1);
  VNStageIntLLRInputS3xD(160)(3) <= CNStageIntLLROutputS3xD(189)(2);
  VNStageIntLLRInputS3xD(248)(3) <= CNStageIntLLROutputS3xD(189)(3);
  VNStageIntLLRInputS3xD(286)(3) <= CNStageIntLLROutputS3xD(189)(4);
  VNStageIntLLRInputS3xD(335)(3) <= CNStageIntLLROutputS3xD(189)(5);
  VNStageIntLLRInputS3xD(41)(3) <= CNStageIntLLROutputS3xD(190)(0);
  VNStageIntLLRInputS3xD(95)(3) <= CNStageIntLLROutputS3xD(190)(1);
  VNStageIntLLRInputS3xD(183)(2) <= CNStageIntLLROutputS3xD(190)(2);
  VNStageIntLLRInputS3xD(221)(3) <= CNStageIntLLROutputS3xD(190)(3);
  VNStageIntLLRInputS3xD(270)(3) <= CNStageIntLLROutputS3xD(190)(4);
  VNStageIntLLRInputS3xD(338)(3) <= CNStageIntLLROutputS3xD(190)(5);
  VNStageIntLLRInputS3xD(39)(3) <= CNStageIntLLROutputS3xD(191)(0);
  VNStageIntLLRInputS3xD(91)(3) <= CNStageIntLLROutputS3xD(191)(1);
  VNStageIntLLRInputS3xD(140)(3) <= CNStageIntLLROutputS3xD(191)(2);
  VNStageIntLLRInputS3xD(208)(3) <= CNStageIntLLROutputS3xD(191)(3);
  VNStageIntLLRInputS3xD(314)(0) <= CNStageIntLLROutputS3xD(191)(4);
  VNStageIntLLRInputS3xD(354)(3) <= CNStageIntLLROutputS3xD(191)(5);
  VNStageIntLLRInputS3xD(38)(3) <= CNStageIntLLROutputS3xD(192)(0);
  VNStageIntLLRInputS3xD(75)(3) <= CNStageIntLLROutputS3xD(192)(1);
  VNStageIntLLRInputS3xD(143)(3) <= CNStageIntLLROutputS3xD(192)(2);
  VNStageIntLLRInputS3xD(249)(1) <= CNStageIntLLROutputS3xD(192)(3);
  VNStageIntLLRInputS3xD(289)(3) <= CNStageIntLLROutputS3xD(192)(4);
  VNStageIntLLRInputS3xD(352)(3) <= CNStageIntLLROutputS3xD(192)(5);
  VNStageIntLLRInputS3xD(37)(3) <= CNStageIntLLROutputS3xD(193)(0);
  VNStageIntLLRInputS3xD(78)(3) <= CNStageIntLLROutputS3xD(193)(1);
  VNStageIntLLRInputS3xD(184)(3) <= CNStageIntLLROutputS3xD(193)(2);
  VNStageIntLLRInputS3xD(224)(3) <= CNStageIntLLROutputS3xD(193)(3);
  VNStageIntLLRInputS3xD(287)(3) <= CNStageIntLLROutputS3xD(193)(4);
  VNStageIntLLRInputS3xD(377)(2) <= CNStageIntLLROutputS3xD(193)(5);
  VNStageIntLLRInputS3xD(35)(3) <= CNStageIntLLROutputS3xD(194)(0);
  VNStageIntLLRInputS3xD(94)(2) <= CNStageIntLLROutputS3xD(194)(1);
  VNStageIntLLRInputS3xD(157)(3) <= CNStageIntLLROutputS3xD(194)(2);
  VNStageIntLLRInputS3xD(247)(3) <= CNStageIntLLROutputS3xD(194)(3);
  VNStageIntLLRInputS3xD(257)(3) <= CNStageIntLLROutputS3xD(194)(4);
  VNStageIntLLRInputS3xD(365)(3) <= CNStageIntLLROutputS3xD(194)(5);
  VNStageIntLLRInputS3xD(34)(3) <= CNStageIntLLROutputS3xD(195)(0);
  VNStageIntLLRInputS3xD(92)(3) <= CNStageIntLLROutputS3xD(195)(1);
  VNStageIntLLRInputS3xD(182)(3) <= CNStageIntLLROutputS3xD(195)(2);
  VNStageIntLLRInputS3xD(255)(3) <= CNStageIntLLROutputS3xD(195)(3);
  VNStageIntLLRInputS3xD(300)(3) <= CNStageIntLLROutputS3xD(195)(4);
  VNStageIntLLRInputS3xD(359)(3) <= CNStageIntLLROutputS3xD(195)(5);
  VNStageIntLLRInputS3xD(33)(3) <= CNStageIntLLROutputS3xD(196)(0);
  VNStageIntLLRInputS3xD(117)(3) <= CNStageIntLLROutputS3xD(196)(1);
  VNStageIntLLRInputS3xD(190)(1) <= CNStageIntLLROutputS3xD(196)(2);
  VNStageIntLLRInputS3xD(235)(2) <= CNStageIntLLROutputS3xD(196)(3);
  VNStageIntLLRInputS3xD(294)(3) <= CNStageIntLLROutputS3xD(196)(4);
  VNStageIntLLRInputS3xD(320)(2) <= CNStageIntLLROutputS3xD(196)(5);
  VNStageIntLLRInputS3xD(31)(2) <= CNStageIntLLROutputS3xD(197)(0);
  VNStageIntLLRInputS3xD(105)(2) <= CNStageIntLLROutputS3xD(197)(1);
  VNStageIntLLRInputS3xD(164)(3) <= CNStageIntLLROutputS3xD(197)(2);
  VNStageIntLLRInputS3xD(192)(3) <= CNStageIntLLROutputS3xD(197)(3);
  VNStageIntLLRInputS3xD(293)(3) <= CNStageIntLLROutputS3xD(197)(4);
  VNStageIntLLRInputS3xD(363)(2) <= CNStageIntLLROutputS3xD(197)(5);
  VNStageIntLLRInputS3xD(30)(3) <= CNStageIntLLROutputS3xD(198)(0);
  VNStageIntLLRInputS3xD(99)(3) <= CNStageIntLLROutputS3xD(198)(1);
  VNStageIntLLRInputS3xD(128)(3) <= CNStageIntLLROutputS3xD(198)(2);
  VNStageIntLLRInputS3xD(228)(3) <= CNStageIntLLROutputS3xD(198)(3);
  VNStageIntLLRInputS3xD(298)(3) <= CNStageIntLLROutputS3xD(198)(4);
  VNStageIntLLRInputS3xD(382)(2) <= CNStageIntLLROutputS3xD(198)(5);
  VNStageIntLLRInputS3xD(28)(3) <= CNStageIntLLROutputS3xD(199)(0);
  VNStageIntLLRInputS3xD(98)(2) <= CNStageIntLLROutputS3xD(199)(1);
  VNStageIntLLRInputS3xD(168)(2) <= CNStageIntLLROutputS3xD(199)(2);
  VNStageIntLLRInputS3xD(252)(2) <= CNStageIntLLROutputS3xD(199)(3);
  VNStageIntLLRInputS3xD(308)(1) <= CNStageIntLLROutputS3xD(199)(4);
  VNStageIntLLRInputS3xD(347)(3) <= CNStageIntLLROutputS3xD(199)(5);
  VNStageIntLLRInputS3xD(27)(3) <= CNStageIntLLROutputS3xD(200)(0);
  VNStageIntLLRInputS3xD(103)(3) <= CNStageIntLLROutputS3xD(200)(1);
  VNStageIntLLRInputS3xD(187)(2) <= CNStageIntLLROutputS3xD(200)(2);
  VNStageIntLLRInputS3xD(243)(3) <= CNStageIntLLROutputS3xD(200)(3);
  VNStageIntLLRInputS3xD(282)(3) <= CNStageIntLLROutputS3xD(200)(4);
  VNStageIntLLRInputS3xD(348)(3) <= CNStageIntLLROutputS3xD(200)(5);
  VNStageIntLLRInputS3xD(26)(3) <= CNStageIntLLROutputS3xD(201)(0);
  VNStageIntLLRInputS3xD(122)(2) <= CNStageIntLLROutputS3xD(201)(1);
  VNStageIntLLRInputS3xD(178)(3) <= CNStageIntLLROutputS3xD(201)(2);
  VNStageIntLLRInputS3xD(217)(3) <= CNStageIntLLROutputS3xD(201)(3);
  VNStageIntLLRInputS3xD(283)(3) <= CNStageIntLLROutputS3xD(201)(4);
  VNStageIntLLRInputS3xD(372)(2) <= CNStageIntLLROutputS3xD(201)(5);
  VNStageIntLLRInputS3xD(25)(3) <= CNStageIntLLROutputS3xD(202)(0);
  VNStageIntLLRInputS3xD(113)(3) <= CNStageIntLLROutputS3xD(202)(1);
  VNStageIntLLRInputS3xD(152)(3) <= CNStageIntLLROutputS3xD(202)(2);
  VNStageIntLLRInputS3xD(218)(3) <= CNStageIntLLROutputS3xD(202)(3);
  VNStageIntLLRInputS3xD(307)(3) <= CNStageIntLLROutputS3xD(202)(4);
  VNStageIntLLRInputS3xD(330)(3) <= CNStageIntLLROutputS3xD(202)(5);
  VNStageIntLLRInputS3xD(24)(3) <= CNStageIntLLROutputS3xD(203)(0);
  VNStageIntLLRInputS3xD(87)(3) <= CNStageIntLLROutputS3xD(203)(1);
  VNStageIntLLRInputS3xD(153)(3) <= CNStageIntLLROutputS3xD(203)(2);
  VNStageIntLLRInputS3xD(242)(3) <= CNStageIntLLROutputS3xD(203)(3);
  VNStageIntLLRInputS3xD(265)(2) <= CNStageIntLLROutputS3xD(203)(4);
  VNStageIntLLRInputS3xD(326)(2) <= CNStageIntLLROutputS3xD(203)(5);
  VNStageIntLLRInputS3xD(23)(3) <= CNStageIntLLROutputS3xD(204)(0);
  VNStageIntLLRInputS3xD(88)(3) <= CNStageIntLLROutputS3xD(204)(1);
  VNStageIntLLRInputS3xD(177)(3) <= CNStageIntLLROutputS3xD(204)(2);
  VNStageIntLLRInputS3xD(200)(3) <= CNStageIntLLROutputS3xD(204)(3);
  VNStageIntLLRInputS3xD(261)(3) <= CNStageIntLLROutputS3xD(204)(4);
  VNStageIntLLRInputS3xD(341)(3) <= CNStageIntLLROutputS3xD(204)(5);
  VNStageIntLLRInputS3xD(22)(3) <= CNStageIntLLROutputS3xD(205)(0);
  VNStageIntLLRInputS3xD(112)(3) <= CNStageIntLLROutputS3xD(205)(1);
  VNStageIntLLRInputS3xD(135)(3) <= CNStageIntLLROutputS3xD(205)(2);
  VNStageIntLLRInputS3xD(196)(3) <= CNStageIntLLROutputS3xD(205)(3);
  VNStageIntLLRInputS3xD(276)(3) <= CNStageIntLLROutputS3xD(205)(4);
  VNStageIntLLRInputS3xD(367)(3) <= CNStageIntLLROutputS3xD(205)(5);
  VNStageIntLLRInputS3xD(21)(3) <= CNStageIntLLROutputS3xD(206)(0);
  VNStageIntLLRInputS3xD(70)(3) <= CNStageIntLLROutputS3xD(206)(1);
  VNStageIntLLRInputS3xD(131)(2) <= CNStageIntLLROutputS3xD(206)(2);
  VNStageIntLLRInputS3xD(211)(3) <= CNStageIntLLROutputS3xD(206)(3);
  VNStageIntLLRInputS3xD(302)(3) <= CNStageIntLLROutputS3xD(206)(4);
  VNStageIntLLRInputS3xD(343)(3) <= CNStageIntLLROutputS3xD(206)(5);
  VNStageIntLLRInputS3xD(18)(3) <= CNStageIntLLROutputS3xD(207)(0);
  VNStageIntLLRInputS3xD(107)(2) <= CNStageIntLLROutputS3xD(207)(1);
  VNStageIntLLRInputS3xD(148)(3) <= CNStageIntLLROutputS3xD(207)(2);
  VNStageIntLLRInputS3xD(245)(3) <= CNStageIntLLROutputS3xD(207)(3);
  VNStageIntLLRInputS3xD(263)(3) <= CNStageIntLLROutputS3xD(207)(4);
  VNStageIntLLRInputS3xD(361)(3) <= CNStageIntLLROutputS3xD(207)(5);
  VNStageIntLLRInputS3xD(17)(3) <= CNStageIntLLROutputS3xD(208)(0);
  VNStageIntLLRInputS3xD(83)(3) <= CNStageIntLLROutputS3xD(208)(1);
  VNStageIntLLRInputS3xD(180)(1) <= CNStageIntLLROutputS3xD(208)(2);
  VNStageIntLLRInputS3xD(198)(3) <= CNStageIntLLROutputS3xD(208)(3);
  VNStageIntLLRInputS3xD(296)(3) <= CNStageIntLLROutputS3xD(208)(4);
  VNStageIntLLRInputS3xD(370)(2) <= CNStageIntLLROutputS3xD(208)(5);
  VNStageIntLLRInputS3xD(16)(2) <= CNStageIntLLROutputS3xD(209)(0);
  VNStageIntLLRInputS3xD(115)(3) <= CNStageIntLLROutputS3xD(209)(1);
  VNStageIntLLRInputS3xD(133)(1) <= CNStageIntLLROutputS3xD(209)(2);
  VNStageIntLLRInputS3xD(231)(2) <= CNStageIntLLROutputS3xD(209)(3);
  VNStageIntLLRInputS3xD(305)(3) <= CNStageIntLLROutputS3xD(209)(4);
  VNStageIntLLRInputS3xD(383)(3) <= CNStageIntLLROutputS3xD(209)(5);
  VNStageIntLLRInputS3xD(15)(3) <= CNStageIntLLROutputS3xD(210)(0);
  VNStageIntLLRInputS3xD(68)(2) <= CNStageIntLLROutputS3xD(210)(1);
  VNStageIntLLRInputS3xD(166)(3) <= CNStageIntLLROutputS3xD(210)(2);
  VNStageIntLLRInputS3xD(240)(3) <= CNStageIntLLROutputS3xD(210)(3);
  VNStageIntLLRInputS3xD(318)(1) <= CNStageIntLLROutputS3xD(210)(4);
  VNStageIntLLRInputS3xD(362)(3) <= CNStageIntLLROutputS3xD(210)(5);
  VNStageIntLLRInputS3xD(14)(3) <= CNStageIntLLROutputS3xD(211)(0);
  VNStageIntLLRInputS3xD(101)(3) <= CNStageIntLLROutputS3xD(211)(1);
  VNStageIntLLRInputS3xD(175)(3) <= CNStageIntLLROutputS3xD(211)(2);
  VNStageIntLLRInputS3xD(253)(2) <= CNStageIntLLROutputS3xD(211)(3);
  VNStageIntLLRInputS3xD(297)(3) <= CNStageIntLLROutputS3xD(211)(4);
  VNStageIntLLRInputS3xD(327)(3) <= CNStageIntLLROutputS3xD(211)(5);
  VNStageIntLLRInputS3xD(13)(2) <= CNStageIntLLROutputS3xD(212)(0);
  VNStageIntLLRInputS3xD(110)(3) <= CNStageIntLLROutputS3xD(212)(1);
  VNStageIntLLRInputS3xD(188)(1) <= CNStageIntLLROutputS3xD(212)(2);
  VNStageIntLLRInputS3xD(232)(2) <= CNStageIntLLROutputS3xD(212)(3);
  VNStageIntLLRInputS3xD(262)(3) <= CNStageIntLLROutputS3xD(212)(4);
  VNStageIntLLRInputS3xD(329)(3) <= CNStageIntLLROutputS3xD(212)(5);
  VNStageIntLLRInputS3xD(12)(3) <= CNStageIntLLROutputS3xD(213)(0);
  VNStageIntLLRInputS3xD(123)(2) <= CNStageIntLLROutputS3xD(213)(1);
  VNStageIntLLRInputS3xD(167)(3) <= CNStageIntLLROutputS3xD(213)(2);
  VNStageIntLLRInputS3xD(197)(3) <= CNStageIntLLROutputS3xD(213)(3);
  VNStageIntLLRInputS3xD(264)(3) <= CNStageIntLLROutputS3xD(213)(4);
  VNStageIntLLRInputS3xD(374)(3) <= CNStageIntLLROutputS3xD(213)(5);
  VNStageIntLLRInputS3xD(11)(3) <= CNStageIntLLROutputS3xD(214)(0);
  VNStageIntLLRInputS3xD(102)(3) <= CNStageIntLLROutputS3xD(214)(1);
  VNStageIntLLRInputS3xD(132)(2) <= CNStageIntLLROutputS3xD(214)(2);
  VNStageIntLLRInputS3xD(199)(3) <= CNStageIntLLROutputS3xD(214)(3);
  VNStageIntLLRInputS3xD(309)(3) <= CNStageIntLLROutputS3xD(214)(4);
  VNStageIntLLRInputS3xD(381)(2) <= CNStageIntLLROutputS3xD(214)(5);
  VNStageIntLLRInputS3xD(9)(3) <= CNStageIntLLROutputS3xD(215)(0);
  VNStageIntLLRInputS3xD(69)(3) <= CNStageIntLLROutputS3xD(215)(1);
  VNStageIntLLRInputS3xD(179)(3) <= CNStageIntLLROutputS3xD(215)(2);
  VNStageIntLLRInputS3xD(251)(2) <= CNStageIntLLROutputS3xD(215)(3);
  VNStageIntLLRInputS3xD(280)(3) <= CNStageIntLLROutputS3xD(215)(4);
  VNStageIntLLRInputS3xD(333)(2) <= CNStageIntLLROutputS3xD(215)(5);
  VNStageIntLLRInputS3xD(8)(2) <= CNStageIntLLROutputS3xD(216)(0);
  VNStageIntLLRInputS3xD(114)(3) <= CNStageIntLLROutputS3xD(216)(1);
  VNStageIntLLRInputS3xD(186)(2) <= CNStageIntLLROutputS3xD(216)(2);
  VNStageIntLLRInputS3xD(215)(3) <= CNStageIntLLROutputS3xD(216)(3);
  VNStageIntLLRInputS3xD(268)(3) <= CNStageIntLLROutputS3xD(216)(4);
  VNStageIntLLRInputS3xD(339)(3) <= CNStageIntLLROutputS3xD(216)(5);
  VNStageIntLLRInputS3xD(7)(3) <= CNStageIntLLROutputS3xD(217)(0);
  VNStageIntLLRInputS3xD(121)(2) <= CNStageIntLLROutputS3xD(217)(1);
  VNStageIntLLRInputS3xD(150)(3) <= CNStageIntLLROutputS3xD(217)(2);
  VNStageIntLLRInputS3xD(203)(3) <= CNStageIntLLROutputS3xD(217)(3);
  VNStageIntLLRInputS3xD(274)(2) <= CNStageIntLLROutputS3xD(217)(4);
  VNStageIntLLRInputS3xD(334)(2) <= CNStageIntLLROutputS3xD(217)(5);
  VNStageIntLLRInputS3xD(6)(3) <= CNStageIntLLROutputS3xD(218)(0);
  VNStageIntLLRInputS3xD(85)(2) <= CNStageIntLLROutputS3xD(218)(1);
  VNStageIntLLRInputS3xD(138)(3) <= CNStageIntLLROutputS3xD(218)(2);
  VNStageIntLLRInputS3xD(209)(3) <= CNStageIntLLROutputS3xD(218)(3);
  VNStageIntLLRInputS3xD(269)(2) <= CNStageIntLLROutputS3xD(218)(4);
  VNStageIntLLRInputS3xD(344)(3) <= CNStageIntLLROutputS3xD(218)(5);
  VNStageIntLLRInputS3xD(5)(3) <= CNStageIntLLROutputS3xD(219)(0);
  VNStageIntLLRInputS3xD(73)(3) <= CNStageIntLLROutputS3xD(219)(1);
  VNStageIntLLRInputS3xD(144)(3) <= CNStageIntLLROutputS3xD(219)(2);
  VNStageIntLLRInputS3xD(204)(3) <= CNStageIntLLROutputS3xD(219)(3);
  VNStageIntLLRInputS3xD(279)(3) <= CNStageIntLLROutputS3xD(219)(4);
  VNStageIntLLRInputS3xD(366)(3) <= CNStageIntLLROutputS3xD(219)(5);
  VNStageIntLLRInputS3xD(4)(2) <= CNStageIntLLROutputS3xD(220)(0);
  VNStageIntLLRInputS3xD(79)(3) <= CNStageIntLLROutputS3xD(220)(1);
  VNStageIntLLRInputS3xD(139)(3) <= CNStageIntLLROutputS3xD(220)(2);
  VNStageIntLLRInputS3xD(214)(3) <= CNStageIntLLROutputS3xD(220)(3);
  VNStageIntLLRInputS3xD(301)(3) <= CNStageIntLLROutputS3xD(220)(4);
  VNStageIntLLRInputS3xD(321)(3) <= CNStageIntLLROutputS3xD(220)(5);
  VNStageIntLLRInputS3xD(3)(2) <= CNStageIntLLROutputS3xD(221)(0);
  VNStageIntLLRInputS3xD(74)(3) <= CNStageIntLLROutputS3xD(221)(1);
  VNStageIntLLRInputS3xD(149)(3) <= CNStageIntLLROutputS3xD(221)(2);
  VNStageIntLLRInputS3xD(236)(3) <= CNStageIntLLROutputS3xD(221)(3);
  VNStageIntLLRInputS3xD(319)(3) <= CNStageIntLLROutputS3xD(221)(4);
  VNStageIntLLRInputS3xD(369)(2) <= CNStageIntLLROutputS3xD(221)(5);
  VNStageIntLLRInputS3xD(2)(3) <= CNStageIntLLROutputS3xD(222)(0);
  VNStageIntLLRInputS3xD(84)(3) <= CNStageIntLLROutputS3xD(222)(1);
  VNStageIntLLRInputS3xD(171)(2) <= CNStageIntLLROutputS3xD(222)(2);
  VNStageIntLLRInputS3xD(254)(1) <= CNStageIntLLROutputS3xD(222)(3);
  VNStageIntLLRInputS3xD(304)(3) <= CNStageIntLLROutputS3xD(222)(4);
  VNStageIntLLRInputS3xD(356)(3) <= CNStageIntLLROutputS3xD(222)(5);
  VNStageIntLLRInputS3xD(1)(2) <= CNStageIntLLROutputS3xD(223)(0);
  VNStageIntLLRInputS3xD(106)(2) <= CNStageIntLLROutputS3xD(223)(1);
  VNStageIntLLRInputS3xD(189)(2) <= CNStageIntLLROutputS3xD(223)(2);
  VNStageIntLLRInputS3xD(239)(3) <= CNStageIntLLROutputS3xD(223)(3);
  VNStageIntLLRInputS3xD(291)(3) <= CNStageIntLLROutputS3xD(223)(4);
  VNStageIntLLRInputS3xD(324)(3) <= CNStageIntLLROutputS3xD(223)(5);
  VNStageIntLLRInputS3xD(0)(3) <= CNStageIntLLROutputS3xD(224)(0);
  VNStageIntLLRInputS3xD(93)(3) <= CNStageIntLLROutputS3xD(224)(1);
  VNStageIntLLRInputS3xD(158)(3) <= CNStageIntLLROutputS3xD(224)(2);
  VNStageIntLLRInputS3xD(223)(3) <= CNStageIntLLROutputS3xD(224)(3);
  VNStageIntLLRInputS3xD(288)(3) <= CNStageIntLLROutputS3xD(224)(4);
  VNStageIntLLRInputS3xD(353)(3) <= CNStageIntLLROutputS3xD(224)(5);
  VNStageIntLLRInputS3xD(18)(4) <= CNStageIntLLROutputS3xD(225)(0);
  VNStageIntLLRInputS3xD(110)(4) <= CNStageIntLLROutputS3xD(225)(1);
  VNStageIntLLRInputS3xD(167)(4) <= CNStageIntLLROutputS3xD(225)(2);
  VNStageIntLLRInputS3xD(249)(2) <= CNStageIntLLROutputS3xD(225)(3);
  VNStageIntLLRInputS3xD(311)(3) <= CNStageIntLLROutputS3xD(225)(4);
  VNStageIntLLRInputS3xD(347)(4) <= CNStageIntLLROutputS3xD(225)(5);
  VNStageIntLLRInputS3xD(17)(4) <= CNStageIntLLROutputS3xD(226)(0);
  VNStageIntLLRInputS3xD(102)(4) <= CNStageIntLLROutputS3xD(226)(1);
  VNStageIntLLRInputS3xD(184)(4) <= CNStageIntLLROutputS3xD(226)(2);
  VNStageIntLLRInputS3xD(246)(4) <= CNStageIntLLROutputS3xD(226)(3);
  VNStageIntLLRInputS3xD(282)(4) <= CNStageIntLLROutputS3xD(226)(4);
  VNStageIntLLRInputS3xD(367)(4) <= CNStageIntLLROutputS3xD(226)(5);
  VNStageIntLLRInputS3xD(16)(3) <= CNStageIntLLROutputS3xD(227)(0);
  VNStageIntLLRInputS3xD(119)(3) <= CNStageIntLLROutputS3xD(227)(1);
  VNStageIntLLRInputS3xD(181)(4) <= CNStageIntLLROutputS3xD(227)(2);
  VNStageIntLLRInputS3xD(217)(4) <= CNStageIntLLROutputS3xD(227)(3);
  VNStageIntLLRInputS3xD(302)(4) <= CNStageIntLLROutputS3xD(227)(4);
  VNStageIntLLRInputS3xD(353)(4) <= CNStageIntLLROutputS3xD(227)(5);
  VNStageIntLLRInputS3xD(15)(4) <= CNStageIntLLROutputS3xD(228)(0);
  VNStageIntLLRInputS3xD(116)(3) <= CNStageIntLLROutputS3xD(228)(1);
  VNStageIntLLRInputS3xD(152)(4) <= CNStageIntLLROutputS3xD(228)(2);
  VNStageIntLLRInputS3xD(237)(3) <= CNStageIntLLROutputS3xD(228)(3);
  VNStageIntLLRInputS3xD(288)(4) <= CNStageIntLLROutputS3xD(228)(4);
  VNStageIntLLRInputS3xD(343)(4) <= CNStageIntLLROutputS3xD(228)(5);
  VNStageIntLLRInputS3xD(14)(4) <= CNStageIntLLROutputS3xD(229)(0);
  VNStageIntLLRInputS3xD(87)(4) <= CNStageIntLLROutputS3xD(229)(1);
  VNStageIntLLRInputS3xD(172)(3) <= CNStageIntLLROutputS3xD(229)(2);
  VNStageIntLLRInputS3xD(223)(4) <= CNStageIntLLROutputS3xD(229)(3);
  VNStageIntLLRInputS3xD(278)(3) <= CNStageIntLLROutputS3xD(229)(4);
  VNStageIntLLRInputS3xD(372)(3) <= CNStageIntLLROutputS3xD(229)(5);
  VNStageIntLLRInputS3xD(13)(3) <= CNStageIntLLROutputS3xD(230)(0);
  VNStageIntLLRInputS3xD(107)(3) <= CNStageIntLLROutputS3xD(230)(1);
  VNStageIntLLRInputS3xD(158)(4) <= CNStageIntLLROutputS3xD(230)(2);
  VNStageIntLLRInputS3xD(213)(3) <= CNStageIntLLROutputS3xD(230)(3);
  VNStageIntLLRInputS3xD(307)(4) <= CNStageIntLLROutputS3xD(230)(4);
  VNStageIntLLRInputS3xD(355)(4) <= CNStageIntLLROutputS3xD(230)(5);
  VNStageIntLLRInputS3xD(12)(4) <= CNStageIntLLROutputS3xD(231)(0);
  VNStageIntLLRInputS3xD(93)(4) <= CNStageIntLLROutputS3xD(231)(1);
  VNStageIntLLRInputS3xD(148)(4) <= CNStageIntLLROutputS3xD(231)(2);
  VNStageIntLLRInputS3xD(242)(4) <= CNStageIntLLROutputS3xD(231)(3);
  VNStageIntLLRInputS3xD(290)(4) <= CNStageIntLLROutputS3xD(231)(4);
  VNStageIntLLRInputS3xD(322)(3) <= CNStageIntLLROutputS3xD(231)(5);
  VNStageIntLLRInputS3xD(11)(4) <= CNStageIntLLROutputS3xD(232)(0);
  VNStageIntLLRInputS3xD(83)(4) <= CNStageIntLLROutputS3xD(232)(1);
  VNStageIntLLRInputS3xD(177)(4) <= CNStageIntLLROutputS3xD(232)(2);
  VNStageIntLLRInputS3xD(225)(4) <= CNStageIntLLROutputS3xD(232)(3);
  VNStageIntLLRInputS3xD(257)(4) <= CNStageIntLLROutputS3xD(232)(4);
  VNStageIntLLRInputS3xD(345)(3) <= CNStageIntLLROutputS3xD(232)(5);
  VNStageIntLLRInputS3xD(10)(3) <= CNStageIntLLROutputS3xD(233)(0);
  VNStageIntLLRInputS3xD(112)(4) <= CNStageIntLLROutputS3xD(233)(1);
  VNStageIntLLRInputS3xD(160)(4) <= CNStageIntLLROutputS3xD(233)(2);
  VNStageIntLLRInputS3xD(255)(4) <= CNStageIntLLROutputS3xD(233)(3);
  VNStageIntLLRInputS3xD(280)(4) <= CNStageIntLLROutputS3xD(233)(4);
  VNStageIntLLRInputS3xD(381)(3) <= CNStageIntLLROutputS3xD(233)(5);
  VNStageIntLLRInputS3xD(9)(4) <= CNStageIntLLROutputS3xD(234)(0);
  VNStageIntLLRInputS3xD(95)(4) <= CNStageIntLLROutputS3xD(234)(1);
  VNStageIntLLRInputS3xD(190)(2) <= CNStageIntLLROutputS3xD(234)(2);
  VNStageIntLLRInputS3xD(215)(4) <= CNStageIntLLROutputS3xD(234)(3);
  VNStageIntLLRInputS3xD(316)(2) <= CNStageIntLLROutputS3xD(234)(4);
  VNStageIntLLRInputS3xD(365)(4) <= CNStageIntLLROutputS3xD(234)(5);
  VNStageIntLLRInputS3xD(7)(4) <= CNStageIntLLROutputS3xD(235)(0);
  VNStageIntLLRInputS3xD(85)(3) <= CNStageIntLLROutputS3xD(235)(1);
  VNStageIntLLRInputS3xD(186)(3) <= CNStageIntLLROutputS3xD(235)(2);
  VNStageIntLLRInputS3xD(235)(3) <= CNStageIntLLROutputS3xD(235)(3);
  VNStageIntLLRInputS3xD(303)(4) <= CNStageIntLLROutputS3xD(235)(4);
  VNStageIntLLRInputS3xD(346)(4) <= CNStageIntLLROutputS3xD(235)(5);
  VNStageIntLLRInputS3xD(6)(4) <= CNStageIntLLROutputS3xD(236)(0);
  VNStageIntLLRInputS3xD(121)(3) <= CNStageIntLLROutputS3xD(236)(1);
  VNStageIntLLRInputS3xD(170)(3) <= CNStageIntLLROutputS3xD(236)(2);
  VNStageIntLLRInputS3xD(238)(4) <= CNStageIntLLROutputS3xD(236)(3);
  VNStageIntLLRInputS3xD(281)(4) <= CNStageIntLLROutputS3xD(236)(4);
  VNStageIntLLRInputS3xD(321)(4) <= CNStageIntLLROutputS3xD(236)(5);
  VNStageIntLLRInputS3xD(5)(4) <= CNStageIntLLROutputS3xD(237)(0);
  VNStageIntLLRInputS3xD(105)(3) <= CNStageIntLLROutputS3xD(237)(1);
  VNStageIntLLRInputS3xD(173)(4) <= CNStageIntLLROutputS3xD(237)(2);
  VNStageIntLLRInputS3xD(216)(4) <= CNStageIntLLROutputS3xD(237)(3);
  VNStageIntLLRInputS3xD(319)(4) <= CNStageIntLLROutputS3xD(237)(4);
  VNStageIntLLRInputS3xD(382)(3) <= CNStageIntLLROutputS3xD(237)(5);
  VNStageIntLLRInputS3xD(4)(3) <= CNStageIntLLROutputS3xD(238)(0);
  VNStageIntLLRInputS3xD(108)(4) <= CNStageIntLLROutputS3xD(238)(1);
  VNStageIntLLRInputS3xD(151)(4) <= CNStageIntLLROutputS3xD(238)(2);
  VNStageIntLLRInputS3xD(254)(2) <= CNStageIntLLROutputS3xD(238)(3);
  VNStageIntLLRInputS3xD(317)(1) <= CNStageIntLLROutputS3xD(238)(4);
  VNStageIntLLRInputS3xD(344)(4) <= CNStageIntLLROutputS3xD(238)(5);
  VNStageIntLLRInputS3xD(3)(3) <= CNStageIntLLROutputS3xD(239)(0);
  VNStageIntLLRInputS3xD(86)(2) <= CNStageIntLLROutputS3xD(239)(1);
  VNStageIntLLRInputS3xD(189)(3) <= CNStageIntLLROutputS3xD(239)(2);
  VNStageIntLLRInputS3xD(252)(3) <= CNStageIntLLROutputS3xD(239)(3);
  VNStageIntLLRInputS3xD(279)(4) <= CNStageIntLLROutputS3xD(239)(4);
  VNStageIntLLRInputS3xD(352)(4) <= CNStageIntLLROutputS3xD(239)(5);
  VNStageIntLLRInputS3xD(2)(4) <= CNStageIntLLROutputS3xD(240)(0);
  VNStageIntLLRInputS3xD(124)(2) <= CNStageIntLLROutputS3xD(240)(1);
  VNStageIntLLRInputS3xD(187)(3) <= CNStageIntLLROutputS3xD(240)(2);
  VNStageIntLLRInputS3xD(214)(4) <= CNStageIntLLROutputS3xD(240)(3);
  VNStageIntLLRInputS3xD(287)(4) <= CNStageIntLLROutputS3xD(240)(4);
  VNStageIntLLRInputS3xD(332)(4) <= CNStageIntLLROutputS3xD(240)(5);
  VNStageIntLLRInputS3xD(1)(3) <= CNStageIntLLROutputS3xD(241)(0);
  VNStageIntLLRInputS3xD(122)(3) <= CNStageIntLLROutputS3xD(241)(1);
  VNStageIntLLRInputS3xD(149)(4) <= CNStageIntLLROutputS3xD(241)(2);
  VNStageIntLLRInputS3xD(222)(2) <= CNStageIntLLROutputS3xD(241)(3);
  VNStageIntLLRInputS3xD(267)(4) <= CNStageIntLLROutputS3xD(241)(4);
  VNStageIntLLRInputS3xD(326)(3) <= CNStageIntLLROutputS3xD(241)(5);
  VNStageIntLLRInputS3xD(62)(3) <= CNStageIntLLROutputS3xD(242)(0);
  VNStageIntLLRInputS3xD(92)(4) <= CNStageIntLLROutputS3xD(242)(1);
  VNStageIntLLRInputS3xD(137)(4) <= CNStageIntLLROutputS3xD(242)(2);
  VNStageIntLLRInputS3xD(196)(4) <= CNStageIntLLROutputS3xD(242)(3);
  VNStageIntLLRInputS3xD(256)(3) <= CNStageIntLLROutputS3xD(242)(4);
  VNStageIntLLRInputS3xD(325)(4) <= CNStageIntLLROutputS3xD(242)(5);
  VNStageIntLLRInputS3xD(61)(3) <= CNStageIntLLROutputS3xD(243)(0);
  VNStageIntLLRInputS3xD(72)(4) <= CNStageIntLLROutputS3xD(243)(1);
  VNStageIntLLRInputS3xD(131)(3) <= CNStageIntLLROutputS3xD(243)(2);
  VNStageIntLLRInputS3xD(192)(4) <= CNStageIntLLROutputS3xD(243)(3);
  VNStageIntLLRInputS3xD(260)(4) <= CNStageIntLLROutputS3xD(243)(4);
  VNStageIntLLRInputS3xD(330)(4) <= CNStageIntLLROutputS3xD(243)(5);
  VNStageIntLLRInputS3xD(60)(3) <= CNStageIntLLROutputS3xD(244)(0);
  VNStageIntLLRInputS3xD(66)(3) <= CNStageIntLLROutputS3xD(244)(1);
  VNStageIntLLRInputS3xD(128)(4) <= CNStageIntLLROutputS3xD(244)(2);
  VNStageIntLLRInputS3xD(195)(3) <= CNStageIntLLROutputS3xD(244)(3);
  VNStageIntLLRInputS3xD(265)(3) <= CNStageIntLLROutputS3xD(244)(4);
  VNStageIntLLRInputS3xD(349)(3) <= CNStageIntLLROutputS3xD(244)(5);
  VNStageIntLLRInputS3xD(59)(2) <= CNStageIntLLROutputS3xD(245)(0);
  VNStageIntLLRInputS3xD(64)(3) <= CNStageIntLLROutputS3xD(245)(1);
  VNStageIntLLRInputS3xD(130)(4) <= CNStageIntLLROutputS3xD(245)(2);
  VNStageIntLLRInputS3xD(200)(4) <= CNStageIntLLROutputS3xD(245)(3);
  VNStageIntLLRInputS3xD(284)(4) <= CNStageIntLLROutputS3xD(245)(4);
  VNStageIntLLRInputS3xD(340)(4) <= CNStageIntLLROutputS3xD(245)(5);
  VNStageIntLLRInputS3xD(57)(3) <= CNStageIntLLROutputS3xD(246)(0);
  VNStageIntLLRInputS3xD(70)(4) <= CNStageIntLLROutputS3xD(246)(1);
  VNStageIntLLRInputS3xD(154)(3) <= CNStageIntLLROutputS3xD(246)(2);
  VNStageIntLLRInputS3xD(210)(4) <= CNStageIntLLROutputS3xD(246)(3);
  VNStageIntLLRInputS3xD(312)(3) <= CNStageIntLLROutputS3xD(246)(4);
  VNStageIntLLRInputS3xD(378)(3) <= CNStageIntLLROutputS3xD(246)(5);
  VNStageIntLLRInputS3xD(56)(4) <= CNStageIntLLROutputS3xD(247)(0);
  VNStageIntLLRInputS3xD(89)(4) <= CNStageIntLLROutputS3xD(247)(1);
  VNStageIntLLRInputS3xD(145)(4) <= CNStageIntLLROutputS3xD(247)(2);
  VNStageIntLLRInputS3xD(247)(4) <= CNStageIntLLROutputS3xD(247)(3);
  VNStageIntLLRInputS3xD(313)(2) <= CNStageIntLLROutputS3xD(247)(4);
  VNStageIntLLRInputS3xD(339)(4) <= CNStageIntLLROutputS3xD(247)(5);
  VNStageIntLLRInputS3xD(55)(4) <= CNStageIntLLROutputS3xD(248)(0);
  VNStageIntLLRInputS3xD(80)(4) <= CNStageIntLLROutputS3xD(248)(1);
  VNStageIntLLRInputS3xD(182)(4) <= CNStageIntLLROutputS3xD(248)(2);
  VNStageIntLLRInputS3xD(248)(4) <= CNStageIntLLROutputS3xD(248)(3);
  VNStageIntLLRInputS3xD(274)(3) <= CNStageIntLLROutputS3xD(248)(4);
  VNStageIntLLRInputS3xD(360)(4) <= CNStageIntLLROutputS3xD(248)(5);
  VNStageIntLLRInputS3xD(53)(3) <= CNStageIntLLROutputS3xD(249)(0);
  VNStageIntLLRInputS3xD(118)(3) <= CNStageIntLLROutputS3xD(249)(1);
  VNStageIntLLRInputS3xD(144)(4) <= CNStageIntLLROutputS3xD(249)(2);
  VNStageIntLLRInputS3xD(230)(3) <= CNStageIntLLROutputS3xD(249)(3);
  VNStageIntLLRInputS3xD(291)(4) <= CNStageIntLLROutputS3xD(249)(4);
  VNStageIntLLRInputS3xD(371)(3) <= CNStageIntLLROutputS3xD(249)(5);
  VNStageIntLLRInputS3xD(51)(3) <= CNStageIntLLROutputS3xD(250)(0);
  VNStageIntLLRInputS3xD(100)(4) <= CNStageIntLLROutputS3xD(250)(1);
  VNStageIntLLRInputS3xD(161)(4) <= CNStageIntLLROutputS3xD(250)(2);
  VNStageIntLLRInputS3xD(241)(3) <= CNStageIntLLROutputS3xD(250)(3);
  VNStageIntLLRInputS3xD(269)(3) <= CNStageIntLLROutputS3xD(250)(4);
  VNStageIntLLRInputS3xD(373)(2) <= CNStageIntLLROutputS3xD(250)(5);
  VNStageIntLLRInputS3xD(50)(4) <= CNStageIntLLROutputS3xD(251)(0);
  VNStageIntLLRInputS3xD(96)(4) <= CNStageIntLLROutputS3xD(251)(1);
  VNStageIntLLRInputS3xD(176)(4) <= CNStageIntLLROutputS3xD(251)(2);
  VNStageIntLLRInputS3xD(204)(4) <= CNStageIntLLROutputS3xD(251)(3);
  VNStageIntLLRInputS3xD(308)(2) <= CNStageIntLLROutputS3xD(251)(4);
  VNStageIntLLRInputS3xD(342)(3) <= CNStageIntLLROutputS3xD(251)(5);
  VNStageIntLLRInputS3xD(49)(4) <= CNStageIntLLROutputS3xD(252)(0);
  VNStageIntLLRInputS3xD(111)(4) <= CNStageIntLLROutputS3xD(252)(1);
  VNStageIntLLRInputS3xD(139)(4) <= CNStageIntLLROutputS3xD(252)(2);
  VNStageIntLLRInputS3xD(243)(4) <= CNStageIntLLROutputS3xD(252)(3);
  VNStageIntLLRInputS3xD(277)(4) <= CNStageIntLLROutputS3xD(252)(4);
  VNStageIntLLRInputS3xD(358)(3) <= CNStageIntLLROutputS3xD(252)(5);
  VNStageIntLLRInputS3xD(47)(2) <= CNStageIntLLROutputS3xD(253)(0);
  VNStageIntLLRInputS3xD(113)(4) <= CNStageIntLLROutputS3xD(253)(1);
  VNStageIntLLRInputS3xD(147)(4) <= CNStageIntLLROutputS3xD(253)(2);
  VNStageIntLLRInputS3xD(228)(4) <= CNStageIntLLROutputS3xD(253)(3);
  VNStageIntLLRInputS3xD(263)(4) <= CNStageIntLLROutputS3xD(253)(4);
  VNStageIntLLRInputS3xD(337)(4) <= CNStageIntLLROutputS3xD(253)(5);
  VNStageIntLLRInputS3xD(46)(4) <= CNStageIntLLROutputS3xD(254)(0);
  VNStageIntLLRInputS3xD(82)(4) <= CNStageIntLLROutputS3xD(254)(1);
  VNStageIntLLRInputS3xD(163)(3) <= CNStageIntLLROutputS3xD(254)(2);
  VNStageIntLLRInputS3xD(198)(4) <= CNStageIntLLROutputS3xD(254)(3);
  VNStageIntLLRInputS3xD(272)(4) <= CNStageIntLLROutputS3xD(254)(4);
  VNStageIntLLRInputS3xD(350)(4) <= CNStageIntLLROutputS3xD(254)(5);
  VNStageIntLLRInputS3xD(45)(4) <= CNStageIntLLROutputS3xD(255)(0);
  VNStageIntLLRInputS3xD(98)(3) <= CNStageIntLLROutputS3xD(255)(1);
  VNStageIntLLRInputS3xD(133)(2) <= CNStageIntLLROutputS3xD(255)(2);
  VNStageIntLLRInputS3xD(207)(3) <= CNStageIntLLROutputS3xD(255)(3);
  VNStageIntLLRInputS3xD(285)(4) <= CNStageIntLLROutputS3xD(255)(4);
  VNStageIntLLRInputS3xD(329)(4) <= CNStageIntLLROutputS3xD(255)(5);
  VNStageIntLLRInputS3xD(44)(4) <= CNStageIntLLROutputS3xD(256)(0);
  VNStageIntLLRInputS3xD(68)(3) <= CNStageIntLLROutputS3xD(256)(1);
  VNStageIntLLRInputS3xD(142)(3) <= CNStageIntLLROutputS3xD(256)(2);
  VNStageIntLLRInputS3xD(220)(4) <= CNStageIntLLROutputS3xD(256)(3);
  VNStageIntLLRInputS3xD(264)(4) <= CNStageIntLLROutputS3xD(256)(4);
  VNStageIntLLRInputS3xD(357)(4) <= CNStageIntLLROutputS3xD(256)(5);
  VNStageIntLLRInputS3xD(43)(3) <= CNStageIntLLROutputS3xD(257)(0);
  VNStageIntLLRInputS3xD(77)(2) <= CNStageIntLLROutputS3xD(257)(1);
  VNStageIntLLRInputS3xD(155)(4) <= CNStageIntLLROutputS3xD(257)(2);
  VNStageIntLLRInputS3xD(199)(4) <= CNStageIntLLROutputS3xD(257)(3);
  VNStageIntLLRInputS3xD(292)(4) <= CNStageIntLLROutputS3xD(257)(4);
  VNStageIntLLRInputS3xD(359)(4) <= CNStageIntLLROutputS3xD(257)(5);
  VNStageIntLLRInputS3xD(42)(4) <= CNStageIntLLROutputS3xD(258)(0);
  VNStageIntLLRInputS3xD(90)(4) <= CNStageIntLLROutputS3xD(258)(1);
  VNStageIntLLRInputS3xD(134)(3) <= CNStageIntLLROutputS3xD(258)(2);
  VNStageIntLLRInputS3xD(227)(4) <= CNStageIntLLROutputS3xD(258)(3);
  VNStageIntLLRInputS3xD(294)(4) <= CNStageIntLLROutputS3xD(258)(4);
  VNStageIntLLRInputS3xD(341)(4) <= CNStageIntLLROutputS3xD(258)(5);
  VNStageIntLLRInputS3xD(41)(4) <= CNStageIntLLROutputS3xD(259)(0);
  VNStageIntLLRInputS3xD(69)(4) <= CNStageIntLLROutputS3xD(259)(1);
  VNStageIntLLRInputS3xD(162)(4) <= CNStageIntLLROutputS3xD(259)(2);
  VNStageIntLLRInputS3xD(229)(3) <= CNStageIntLLROutputS3xD(259)(3);
  VNStageIntLLRInputS3xD(276)(4) <= CNStageIntLLROutputS3xD(259)(4);
  VNStageIntLLRInputS3xD(348)(4) <= CNStageIntLLROutputS3xD(259)(5);
  VNStageIntLLRInputS3xD(40)(3) <= CNStageIntLLROutputS3xD(260)(0);
  VNStageIntLLRInputS3xD(97)(4) <= CNStageIntLLROutputS3xD(260)(1);
  VNStageIntLLRInputS3xD(164)(4) <= CNStageIntLLROutputS3xD(260)(2);
  VNStageIntLLRInputS3xD(211)(4) <= CNStageIntLLROutputS3xD(260)(3);
  VNStageIntLLRInputS3xD(283)(4) <= CNStageIntLLROutputS3xD(260)(4);
  VNStageIntLLRInputS3xD(375)(3) <= CNStageIntLLROutputS3xD(260)(5);
  VNStageIntLLRInputS3xD(39)(4) <= CNStageIntLLROutputS3xD(261)(0);
  VNStageIntLLRInputS3xD(99)(4) <= CNStageIntLLROutputS3xD(261)(1);
  VNStageIntLLRInputS3xD(146)(3) <= CNStageIntLLROutputS3xD(261)(2);
  VNStageIntLLRInputS3xD(218)(4) <= CNStageIntLLROutputS3xD(261)(3);
  VNStageIntLLRInputS3xD(310)(3) <= CNStageIntLLROutputS3xD(261)(4);
  VNStageIntLLRInputS3xD(363)(3) <= CNStageIntLLROutputS3xD(261)(5);
  VNStageIntLLRInputS3xD(38)(4) <= CNStageIntLLROutputS3xD(262)(0);
  VNStageIntLLRInputS3xD(81)(3) <= CNStageIntLLROutputS3xD(262)(1);
  VNStageIntLLRInputS3xD(153)(4) <= CNStageIntLLROutputS3xD(262)(2);
  VNStageIntLLRInputS3xD(245)(4) <= CNStageIntLLROutputS3xD(262)(3);
  VNStageIntLLRInputS3xD(298)(4) <= CNStageIntLLROutputS3xD(262)(4);
  VNStageIntLLRInputS3xD(369)(3) <= CNStageIntLLROutputS3xD(262)(5);
  VNStageIntLLRInputS3xD(37)(4) <= CNStageIntLLROutputS3xD(263)(0);
  VNStageIntLLRInputS3xD(88)(4) <= CNStageIntLLROutputS3xD(263)(1);
  VNStageIntLLRInputS3xD(180)(2) <= CNStageIntLLROutputS3xD(263)(2);
  VNStageIntLLRInputS3xD(233)(3) <= CNStageIntLLROutputS3xD(263)(3);
  VNStageIntLLRInputS3xD(304)(4) <= CNStageIntLLROutputS3xD(263)(4);
  VNStageIntLLRInputS3xD(364)(4) <= CNStageIntLLROutputS3xD(263)(5);
  VNStageIntLLRInputS3xD(36)(3) <= CNStageIntLLROutputS3xD(264)(0);
  VNStageIntLLRInputS3xD(115)(4) <= CNStageIntLLROutputS3xD(264)(1);
  VNStageIntLLRInputS3xD(168)(3) <= CNStageIntLLROutputS3xD(264)(2);
  VNStageIntLLRInputS3xD(239)(4) <= CNStageIntLLROutputS3xD(264)(3);
  VNStageIntLLRInputS3xD(299)(3) <= CNStageIntLLROutputS3xD(264)(4);
  VNStageIntLLRInputS3xD(374)(4) <= CNStageIntLLROutputS3xD(264)(5);
  VNStageIntLLRInputS3xD(35)(4) <= CNStageIntLLROutputS3xD(265)(0);
  VNStageIntLLRInputS3xD(103)(4) <= CNStageIntLLROutputS3xD(265)(1);
  VNStageIntLLRInputS3xD(174)(3) <= CNStageIntLLROutputS3xD(265)(2);
  VNStageIntLLRInputS3xD(234)(4) <= CNStageIntLLROutputS3xD(265)(3);
  VNStageIntLLRInputS3xD(309)(4) <= CNStageIntLLROutputS3xD(265)(4);
  VNStageIntLLRInputS3xD(333)(3) <= CNStageIntLLROutputS3xD(265)(5);
  VNStageIntLLRInputS3xD(34)(4) <= CNStageIntLLROutputS3xD(266)(0);
  VNStageIntLLRInputS3xD(109)(4) <= CNStageIntLLROutputS3xD(266)(1);
  VNStageIntLLRInputS3xD(169)(4) <= CNStageIntLLROutputS3xD(266)(2);
  VNStageIntLLRInputS3xD(244)(1) <= CNStageIntLLROutputS3xD(266)(3);
  VNStageIntLLRInputS3xD(268)(4) <= CNStageIntLLROutputS3xD(266)(4);
  VNStageIntLLRInputS3xD(351)(3) <= CNStageIntLLROutputS3xD(266)(5);
  VNStageIntLLRInputS3xD(33)(4) <= CNStageIntLLROutputS3xD(267)(0);
  VNStageIntLLRInputS3xD(104)(4) <= CNStageIntLLROutputS3xD(267)(1);
  VNStageIntLLRInputS3xD(179)(4) <= CNStageIntLLROutputS3xD(267)(2);
  VNStageIntLLRInputS3xD(203)(4) <= CNStageIntLLROutputS3xD(267)(3);
  VNStageIntLLRInputS3xD(286)(4) <= CNStageIntLLROutputS3xD(267)(4);
  VNStageIntLLRInputS3xD(336)(3) <= CNStageIntLLROutputS3xD(267)(5);
  VNStageIntLLRInputS3xD(32)(3) <= CNStageIntLLROutputS3xD(268)(0);
  VNStageIntLLRInputS3xD(114)(4) <= CNStageIntLLROutputS3xD(268)(1);
  VNStageIntLLRInputS3xD(138)(4) <= CNStageIntLLROutputS3xD(268)(2);
  VNStageIntLLRInputS3xD(221)(4) <= CNStageIntLLROutputS3xD(268)(3);
  VNStageIntLLRInputS3xD(271)(3) <= CNStageIntLLROutputS3xD(268)(4);
  VNStageIntLLRInputS3xD(323)(3) <= CNStageIntLLROutputS3xD(268)(5);
  VNStageIntLLRInputS3xD(30)(4) <= CNStageIntLLROutputS3xD(269)(0);
  VNStageIntLLRInputS3xD(91)(4) <= CNStageIntLLROutputS3xD(269)(1);
  VNStageIntLLRInputS3xD(141)(2) <= CNStageIntLLROutputS3xD(269)(2);
  VNStageIntLLRInputS3xD(193)(3) <= CNStageIntLLROutputS3xD(269)(3);
  VNStageIntLLRInputS3xD(289)(4) <= CNStageIntLLROutputS3xD(269)(4);
  VNStageIntLLRInputS3xD(366)(4) <= CNStageIntLLROutputS3xD(269)(5);
  VNStageIntLLRInputS3xD(29)(3) <= CNStageIntLLROutputS3xD(270)(0);
  VNStageIntLLRInputS3xD(76)(4) <= CNStageIntLLROutputS3xD(270)(1);
  VNStageIntLLRInputS3xD(191)(4) <= CNStageIntLLROutputS3xD(270)(2);
  VNStageIntLLRInputS3xD(224)(4) <= CNStageIntLLROutputS3xD(270)(3);
  VNStageIntLLRInputS3xD(301)(4) <= CNStageIntLLROutputS3xD(270)(4);
  VNStageIntLLRInputS3xD(380)(3) <= CNStageIntLLROutputS3xD(270)(5);
  VNStageIntLLRInputS3xD(28)(4) <= CNStageIntLLROutputS3xD(271)(0);
  VNStageIntLLRInputS3xD(126)(3) <= CNStageIntLLROutputS3xD(271)(1);
  VNStageIntLLRInputS3xD(159)(3) <= CNStageIntLLROutputS3xD(271)(2);
  VNStageIntLLRInputS3xD(236)(4) <= CNStageIntLLROutputS3xD(271)(3);
  VNStageIntLLRInputS3xD(315)(3) <= CNStageIntLLROutputS3xD(271)(4);
  VNStageIntLLRInputS3xD(361)(4) <= CNStageIntLLROutputS3xD(271)(5);
  VNStageIntLLRInputS3xD(26)(4) <= CNStageIntLLROutputS3xD(272)(0);
  VNStageIntLLRInputS3xD(106)(3) <= CNStageIntLLROutputS3xD(272)(1);
  VNStageIntLLRInputS3xD(185)(1) <= CNStageIntLLROutputS3xD(272)(2);
  VNStageIntLLRInputS3xD(231)(3) <= CNStageIntLLROutputS3xD(272)(3);
  VNStageIntLLRInputS3xD(273)(3) <= CNStageIntLLROutputS3xD(272)(4);
  VNStageIntLLRInputS3xD(327)(4) <= CNStageIntLLROutputS3xD(272)(5);
  VNStageIntLLRInputS3xD(24)(4) <= CNStageIntLLROutputS3xD(273)(0);
  VNStageIntLLRInputS3xD(101)(4) <= CNStageIntLLROutputS3xD(273)(1);
  VNStageIntLLRInputS3xD(143)(4) <= CNStageIntLLROutputS3xD(273)(2);
  VNStageIntLLRInputS3xD(197)(4) <= CNStageIntLLROutputS3xD(273)(3);
  VNStageIntLLRInputS3xD(266)(3) <= CNStageIntLLROutputS3xD(273)(4);
  VNStageIntLLRInputS3xD(324)(4) <= CNStageIntLLROutputS3xD(273)(5);
  VNStageIntLLRInputS3xD(23)(4) <= CNStageIntLLROutputS3xD(274)(0);
  VNStageIntLLRInputS3xD(78)(4) <= CNStageIntLLROutputS3xD(274)(1);
  VNStageIntLLRInputS3xD(132)(3) <= CNStageIntLLROutputS3xD(274)(2);
  VNStageIntLLRInputS3xD(201)(4) <= CNStageIntLLROutputS3xD(274)(3);
  VNStageIntLLRInputS3xD(259)(2) <= CNStageIntLLROutputS3xD(274)(4);
  VNStageIntLLRInputS3xD(335)(4) <= CNStageIntLLROutputS3xD(274)(5);
  VNStageIntLLRInputS3xD(22)(4) <= CNStageIntLLROutputS3xD(275)(0);
  VNStageIntLLRInputS3xD(67)(1) <= CNStageIntLLROutputS3xD(275)(1);
  VNStageIntLLRInputS3xD(136)(4) <= CNStageIntLLROutputS3xD(275)(2);
  VNStageIntLLRInputS3xD(194)(4) <= CNStageIntLLROutputS3xD(275)(3);
  VNStageIntLLRInputS3xD(270)(4) <= CNStageIntLLROutputS3xD(275)(4);
  VNStageIntLLRInputS3xD(370)(3) <= CNStageIntLLROutputS3xD(275)(5);
  VNStageIntLLRInputS3xD(21)(4) <= CNStageIntLLROutputS3xD(276)(0);
  VNStageIntLLRInputS3xD(71)(3) <= CNStageIntLLROutputS3xD(276)(1);
  VNStageIntLLRInputS3xD(129)(4) <= CNStageIntLLROutputS3xD(276)(2);
  VNStageIntLLRInputS3xD(205)(1) <= CNStageIntLLROutputS3xD(276)(3);
  VNStageIntLLRInputS3xD(305)(4) <= CNStageIntLLROutputS3xD(276)(4);
  VNStageIntLLRInputS3xD(362)(4) <= CNStageIntLLROutputS3xD(276)(5);
  VNStageIntLLRInputS3xD(20)(2) <= CNStageIntLLROutputS3xD(277)(0);
  VNStageIntLLRInputS3xD(127)(4) <= CNStageIntLLROutputS3xD(277)(1);
  VNStageIntLLRInputS3xD(140)(4) <= CNStageIntLLROutputS3xD(277)(2);
  VNStageIntLLRInputS3xD(240)(4) <= CNStageIntLLROutputS3xD(277)(3);
  VNStageIntLLRInputS3xD(297)(4) <= CNStageIntLLROutputS3xD(277)(4);
  VNStageIntLLRInputS3xD(379)(2) <= CNStageIntLLROutputS3xD(277)(5);
  VNStageIntLLRInputS3xD(19)(3) <= CNStageIntLLROutputS3xD(278)(0);
  VNStageIntLLRInputS3xD(75)(4) <= CNStageIntLLROutputS3xD(278)(1);
  VNStageIntLLRInputS3xD(175)(4) <= CNStageIntLLROutputS3xD(278)(2);
  VNStageIntLLRInputS3xD(232)(3) <= CNStageIntLLROutputS3xD(278)(3);
  VNStageIntLLRInputS3xD(314)(1) <= CNStageIntLLROutputS3xD(278)(4);
  VNStageIntLLRInputS3xD(376)(3) <= CNStageIntLLROutputS3xD(278)(5);
  VNStageIntLLRInputS3xD(0)(4) <= CNStageIntLLROutputS3xD(279)(0);
  VNStageIntLLRInputS3xD(123)(3) <= CNStageIntLLROutputS3xD(279)(1);
  VNStageIntLLRInputS3xD(188)(2) <= CNStageIntLLROutputS3xD(279)(2);
  VNStageIntLLRInputS3xD(253)(3) <= CNStageIntLLROutputS3xD(279)(3);
  VNStageIntLLRInputS3xD(318)(2) <= CNStageIntLLROutputS3xD(279)(4);
  VNStageIntLLRInputS3xD(383)(4) <= CNStageIntLLROutputS3xD(279)(5);
  VNStageIntLLRInputS3xD(35)(5) <= CNStageIntLLROutputS3xD(280)(0);
  VNStageIntLLRInputS3xD(91)(5) <= CNStageIntLLROutputS3xD(280)(1);
  VNStageIntLLRInputS3xD(191)(5) <= CNStageIntLLROutputS3xD(280)(2);
  VNStageIntLLRInputS3xD(248)(5) <= CNStageIntLLROutputS3xD(280)(3);
  VNStageIntLLRInputS3xD(267)(5) <= CNStageIntLLROutputS3xD(280)(4);
  VNStageIntLLRInputS3xD(329)(5) <= CNStageIntLLROutputS3xD(280)(5);
  VNStageIntLLRInputS3xD(34)(5) <= CNStageIntLLROutputS3xD(281)(0);
  VNStageIntLLRInputS3xD(126)(4) <= CNStageIntLLROutputS3xD(281)(1);
  VNStageIntLLRInputS3xD(183)(3) <= CNStageIntLLROutputS3xD(281)(2);
  VNStageIntLLRInputS3xD(202)(4) <= CNStageIntLLROutputS3xD(281)(3);
  VNStageIntLLRInputS3xD(264)(5) <= CNStageIntLLROutputS3xD(281)(4);
  VNStageIntLLRInputS3xD(363)(4) <= CNStageIntLLROutputS3xD(281)(5);
  VNStageIntLLRInputS3xD(33)(5) <= CNStageIntLLROutputS3xD(282)(0);
  VNStageIntLLRInputS3xD(118)(4) <= CNStageIntLLROutputS3xD(282)(1);
  VNStageIntLLRInputS3xD(137)(5) <= CNStageIntLLROutputS3xD(282)(2);
  VNStageIntLLRInputS3xD(199)(5) <= CNStageIntLLROutputS3xD(282)(3);
  VNStageIntLLRInputS3xD(298)(5) <= CNStageIntLLROutputS3xD(282)(4);
  VNStageIntLLRInputS3xD(383)(5) <= CNStageIntLLROutputS3xD(282)(5);
  VNStageIntLLRInputS3xD(31)(3) <= CNStageIntLLROutputS3xD(283)(0);
  VNStageIntLLRInputS3xD(69)(5) <= CNStageIntLLROutputS3xD(283)(1);
  VNStageIntLLRInputS3xD(168)(4) <= CNStageIntLLROutputS3xD(283)(2);
  VNStageIntLLRInputS3xD(253)(4) <= CNStageIntLLROutputS3xD(283)(3);
  VNStageIntLLRInputS3xD(304)(5) <= CNStageIntLLROutputS3xD(283)(4);
  VNStageIntLLRInputS3xD(359)(5) <= CNStageIntLLROutputS3xD(283)(5);
  VNStageIntLLRInputS3xD(30)(5) <= CNStageIntLLROutputS3xD(284)(0);
  VNStageIntLLRInputS3xD(103)(5) <= CNStageIntLLROutputS3xD(284)(1);
  VNStageIntLLRInputS3xD(188)(3) <= CNStageIntLLROutputS3xD(284)(2);
  VNStageIntLLRInputS3xD(239)(5) <= CNStageIntLLROutputS3xD(284)(3);
  VNStageIntLLRInputS3xD(294)(5) <= CNStageIntLLROutputS3xD(284)(4);
  VNStageIntLLRInputS3xD(325)(5) <= CNStageIntLLROutputS3xD(284)(5);
  VNStageIntLLRInputS3xD(27)(4) <= CNStageIntLLROutputS3xD(285)(0);
  VNStageIntLLRInputS3xD(99)(5) <= CNStageIntLLROutputS3xD(285)(1);
  VNStageIntLLRInputS3xD(130)(5) <= CNStageIntLLROutputS3xD(285)(2);
  VNStageIntLLRInputS3xD(241)(4) <= CNStageIntLLROutputS3xD(285)(3);
  VNStageIntLLRInputS3xD(273)(4) <= CNStageIntLLROutputS3xD(285)(4);
  VNStageIntLLRInputS3xD(361)(5) <= CNStageIntLLROutputS3xD(285)(5);
  VNStageIntLLRInputS3xD(26)(5) <= CNStageIntLLROutputS3xD(286)(0);
  VNStageIntLLRInputS3xD(65)(4) <= CNStageIntLLROutputS3xD(286)(1);
  VNStageIntLLRInputS3xD(176)(5) <= CNStageIntLLROutputS3xD(286)(2);
  VNStageIntLLRInputS3xD(208)(4) <= CNStageIntLLROutputS3xD(286)(3);
  VNStageIntLLRInputS3xD(296)(4) <= CNStageIntLLROutputS3xD(286)(4);
  VNStageIntLLRInputS3xD(334)(3) <= CNStageIntLLROutputS3xD(286)(5);
  VNStageIntLLRInputS3xD(25)(4) <= CNStageIntLLROutputS3xD(287)(0);
  VNStageIntLLRInputS3xD(111)(5) <= CNStageIntLLROutputS3xD(287)(1);
  VNStageIntLLRInputS3xD(143)(5) <= CNStageIntLLROutputS3xD(287)(2);
  VNStageIntLLRInputS3xD(231)(4) <= CNStageIntLLROutputS3xD(287)(3);
  VNStageIntLLRInputS3xD(269)(4) <= CNStageIntLLROutputS3xD(287)(4);
  VNStageIntLLRInputS3xD(381)(4) <= CNStageIntLLROutputS3xD(287)(5);
  VNStageIntLLRInputS3xD(24)(5) <= CNStageIntLLROutputS3xD(288)(0);
  VNStageIntLLRInputS3xD(78)(5) <= CNStageIntLLROutputS3xD(288)(1);
  VNStageIntLLRInputS3xD(166)(4) <= CNStageIntLLROutputS3xD(288)(2);
  VNStageIntLLRInputS3xD(204)(5) <= CNStageIntLLROutputS3xD(288)(3);
  VNStageIntLLRInputS3xD(316)(3) <= CNStageIntLLROutputS3xD(288)(4);
  VNStageIntLLRInputS3xD(321)(5) <= CNStageIntLLROutputS3xD(288)(5);
  VNStageIntLLRInputS3xD(23)(5) <= CNStageIntLLROutputS3xD(289)(0);
  VNStageIntLLRInputS3xD(101)(5) <= CNStageIntLLROutputS3xD(289)(1);
  VNStageIntLLRInputS3xD(139)(5) <= CNStageIntLLROutputS3xD(289)(2);
  VNStageIntLLRInputS3xD(251)(3) <= CNStageIntLLROutputS3xD(289)(3);
  VNStageIntLLRInputS3xD(319)(5) <= CNStageIntLLROutputS3xD(289)(4);
  VNStageIntLLRInputS3xD(362)(5) <= CNStageIntLLROutputS3xD(289)(5);
  VNStageIntLLRInputS3xD(22)(5) <= CNStageIntLLROutputS3xD(290)(0);
  VNStageIntLLRInputS3xD(74)(4) <= CNStageIntLLROutputS3xD(290)(1);
  VNStageIntLLRInputS3xD(186)(4) <= CNStageIntLLROutputS3xD(290)(2);
  VNStageIntLLRInputS3xD(254)(3) <= CNStageIntLLROutputS3xD(290)(3);
  VNStageIntLLRInputS3xD(297)(5) <= CNStageIntLLROutputS3xD(290)(4);
  VNStageIntLLRInputS3xD(337)(5) <= CNStageIntLLROutputS3xD(290)(5);
  VNStageIntLLRInputS3xD(21)(5) <= CNStageIntLLROutputS3xD(291)(0);
  VNStageIntLLRInputS3xD(121)(4) <= CNStageIntLLROutputS3xD(291)(1);
  VNStageIntLLRInputS3xD(189)(4) <= CNStageIntLLROutputS3xD(291)(2);
  VNStageIntLLRInputS3xD(232)(4) <= CNStageIntLLROutputS3xD(291)(3);
  VNStageIntLLRInputS3xD(272)(5) <= CNStageIntLLROutputS3xD(291)(4);
  VNStageIntLLRInputS3xD(335)(5) <= CNStageIntLLROutputS3xD(291)(5);
  VNStageIntLLRInputS3xD(20)(3) <= CNStageIntLLROutputS3xD(292)(0);
  VNStageIntLLRInputS3xD(124)(3) <= CNStageIntLLROutputS3xD(292)(1);
  VNStageIntLLRInputS3xD(167)(5) <= CNStageIntLLROutputS3xD(292)(2);
  VNStageIntLLRInputS3xD(207)(4) <= CNStageIntLLROutputS3xD(292)(3);
  VNStageIntLLRInputS3xD(270)(5) <= CNStageIntLLROutputS3xD(292)(4);
  VNStageIntLLRInputS3xD(360)(5) <= CNStageIntLLROutputS3xD(292)(5);
  VNStageIntLLRInputS3xD(18)(5) <= CNStageIntLLROutputS3xD(293)(0);
  VNStageIntLLRInputS3xD(77)(3) <= CNStageIntLLROutputS3xD(293)(1);
  VNStageIntLLRInputS3xD(140)(5) <= CNStageIntLLROutputS3xD(293)(2);
  VNStageIntLLRInputS3xD(230)(4) <= CNStageIntLLROutputS3xD(293)(3);
  VNStageIntLLRInputS3xD(303)(5) <= CNStageIntLLROutputS3xD(293)(4);
  VNStageIntLLRInputS3xD(348)(5) <= CNStageIntLLROutputS3xD(293)(5);
  VNStageIntLLRInputS3xD(17)(5) <= CNStageIntLLROutputS3xD(294)(0);
  VNStageIntLLRInputS3xD(75)(5) <= CNStageIntLLROutputS3xD(294)(1);
  VNStageIntLLRInputS3xD(165)(4) <= CNStageIntLLROutputS3xD(294)(2);
  VNStageIntLLRInputS3xD(238)(5) <= CNStageIntLLROutputS3xD(294)(3);
  VNStageIntLLRInputS3xD(283)(5) <= CNStageIntLLROutputS3xD(294)(4);
  VNStageIntLLRInputS3xD(342)(4) <= CNStageIntLLROutputS3xD(294)(5);
  VNStageIntLLRInputS3xD(16)(4) <= CNStageIntLLROutputS3xD(295)(0);
  VNStageIntLLRInputS3xD(100)(5) <= CNStageIntLLROutputS3xD(295)(1);
  VNStageIntLLRInputS3xD(173)(5) <= CNStageIntLLROutputS3xD(295)(2);
  VNStageIntLLRInputS3xD(218)(5) <= CNStageIntLLROutputS3xD(295)(3);
  VNStageIntLLRInputS3xD(277)(5) <= CNStageIntLLROutputS3xD(295)(4);
  VNStageIntLLRInputS3xD(320)(3) <= CNStageIntLLROutputS3xD(295)(5);
  VNStageIntLLRInputS3xD(15)(5) <= CNStageIntLLROutputS3xD(296)(0);
  VNStageIntLLRInputS3xD(108)(5) <= CNStageIntLLROutputS3xD(296)(1);
  VNStageIntLLRInputS3xD(153)(5) <= CNStageIntLLROutputS3xD(296)(2);
  VNStageIntLLRInputS3xD(212)(4) <= CNStageIntLLROutputS3xD(296)(3);
  VNStageIntLLRInputS3xD(256)(4) <= CNStageIntLLROutputS3xD(296)(4);
  VNStageIntLLRInputS3xD(341)(5) <= CNStageIntLLROutputS3xD(296)(5);
  VNStageIntLLRInputS3xD(14)(5) <= CNStageIntLLROutputS3xD(297)(0);
  VNStageIntLLRInputS3xD(88)(5) <= CNStageIntLLROutputS3xD(297)(1);
  VNStageIntLLRInputS3xD(147)(5) <= CNStageIntLLROutputS3xD(297)(2);
  VNStageIntLLRInputS3xD(192)(5) <= CNStageIntLLROutputS3xD(297)(3);
  VNStageIntLLRInputS3xD(276)(5) <= CNStageIntLLROutputS3xD(297)(4);
  VNStageIntLLRInputS3xD(346)(5) <= CNStageIntLLROutputS3xD(297)(5);
  VNStageIntLLRInputS3xD(13)(4) <= CNStageIntLLROutputS3xD(298)(0);
  VNStageIntLLRInputS3xD(82)(5) <= CNStageIntLLROutputS3xD(298)(1);
  VNStageIntLLRInputS3xD(128)(5) <= CNStageIntLLROutputS3xD(298)(2);
  VNStageIntLLRInputS3xD(211)(5) <= CNStageIntLLROutputS3xD(298)(3);
  VNStageIntLLRInputS3xD(281)(5) <= CNStageIntLLROutputS3xD(298)(4);
  VNStageIntLLRInputS3xD(365)(5) <= CNStageIntLLROutputS3xD(298)(5);
  VNStageIntLLRInputS3xD(12)(5) <= CNStageIntLLROutputS3xD(299)(0);
  VNStageIntLLRInputS3xD(64)(4) <= CNStageIntLLROutputS3xD(299)(1);
  VNStageIntLLRInputS3xD(146)(4) <= CNStageIntLLROutputS3xD(299)(2);
  VNStageIntLLRInputS3xD(216)(5) <= CNStageIntLLROutputS3xD(299)(3);
  VNStageIntLLRInputS3xD(300)(4) <= CNStageIntLLROutputS3xD(299)(4);
  VNStageIntLLRInputS3xD(356)(4) <= CNStageIntLLROutputS3xD(299)(5);
  VNStageIntLLRInputS3xD(9)(5) <= CNStageIntLLROutputS3xD(300)(0);
  VNStageIntLLRInputS3xD(105)(4) <= CNStageIntLLROutputS3xD(300)(1);
  VNStageIntLLRInputS3xD(161)(5) <= CNStageIntLLROutputS3xD(300)(2);
  VNStageIntLLRInputS3xD(200)(5) <= CNStageIntLLROutputS3xD(300)(3);
  VNStageIntLLRInputS3xD(266)(4) <= CNStageIntLLROutputS3xD(300)(4);
  VNStageIntLLRInputS3xD(355)(5) <= CNStageIntLLROutputS3xD(300)(5);
  VNStageIntLLRInputS3xD(7)(5) <= CNStageIntLLROutputS3xD(301)(0);
  VNStageIntLLRInputS3xD(70)(5) <= CNStageIntLLROutputS3xD(301)(1);
  VNStageIntLLRInputS3xD(136)(5) <= CNStageIntLLROutputS3xD(301)(2);
  VNStageIntLLRInputS3xD(225)(5) <= CNStageIntLLROutputS3xD(301)(3);
  VNStageIntLLRInputS3xD(311)(4) <= CNStageIntLLROutputS3xD(301)(4);
  VNStageIntLLRInputS3xD(372)(4) <= CNStageIntLLROutputS3xD(301)(5);
  VNStageIntLLRInputS3xD(6)(5) <= CNStageIntLLROutputS3xD(302)(0);
  VNStageIntLLRInputS3xD(71)(4) <= CNStageIntLLROutputS3xD(302)(1);
  VNStageIntLLRInputS3xD(160)(5) <= CNStageIntLLROutputS3xD(302)(2);
  VNStageIntLLRInputS3xD(246)(5) <= CNStageIntLLROutputS3xD(302)(3);
  VNStageIntLLRInputS3xD(307)(5) <= CNStageIntLLROutputS3xD(302)(4);
  VNStageIntLLRInputS3xD(324)(5) <= CNStageIntLLROutputS3xD(302)(5);
  VNStageIntLLRInputS3xD(5)(5) <= CNStageIntLLROutputS3xD(303)(0);
  VNStageIntLLRInputS3xD(95)(5) <= CNStageIntLLROutputS3xD(303)(1);
  VNStageIntLLRInputS3xD(181)(5) <= CNStageIntLLROutputS3xD(303)(2);
  VNStageIntLLRInputS3xD(242)(5) <= CNStageIntLLROutputS3xD(303)(3);
  VNStageIntLLRInputS3xD(259)(3) <= CNStageIntLLROutputS3xD(303)(4);
  VNStageIntLLRInputS3xD(350)(5) <= CNStageIntLLROutputS3xD(303)(5);
  VNStageIntLLRInputS3xD(4)(4) <= CNStageIntLLROutputS3xD(304)(0);
  VNStageIntLLRInputS3xD(116)(4) <= CNStageIntLLROutputS3xD(304)(1);
  VNStageIntLLRInputS3xD(177)(5) <= CNStageIntLLROutputS3xD(304)(2);
  VNStageIntLLRInputS3xD(194)(5) <= CNStageIntLLROutputS3xD(304)(3);
  VNStageIntLLRInputS3xD(285)(5) <= CNStageIntLLROutputS3xD(304)(4);
  VNStageIntLLRInputS3xD(326)(4) <= CNStageIntLLROutputS3xD(304)(5);
  VNStageIntLLRInputS3xD(3)(4) <= CNStageIntLLROutputS3xD(305)(0);
  VNStageIntLLRInputS3xD(112)(5) <= CNStageIntLLROutputS3xD(305)(1);
  VNStageIntLLRInputS3xD(129)(5) <= CNStageIntLLROutputS3xD(305)(2);
  VNStageIntLLRInputS3xD(220)(5) <= CNStageIntLLROutputS3xD(305)(3);
  VNStageIntLLRInputS3xD(261)(4) <= CNStageIntLLROutputS3xD(305)(4);
  VNStageIntLLRInputS3xD(358)(4) <= CNStageIntLLROutputS3xD(305)(5);
  VNStageIntLLRInputS3xD(2)(5) <= CNStageIntLLROutputS3xD(306)(0);
  VNStageIntLLRInputS3xD(127)(5) <= CNStageIntLLROutputS3xD(306)(1);
  VNStageIntLLRInputS3xD(155)(5) <= CNStageIntLLROutputS3xD(306)(2);
  VNStageIntLLRInputS3xD(196)(5) <= CNStageIntLLROutputS3xD(306)(3);
  VNStageIntLLRInputS3xD(293)(4) <= CNStageIntLLROutputS3xD(306)(4);
  VNStageIntLLRInputS3xD(374)(5) <= CNStageIntLLROutputS3xD(306)(5);
  VNStageIntLLRInputS3xD(1)(4) <= CNStageIntLLROutputS3xD(307)(0);
  VNStageIntLLRInputS3xD(90)(5) <= CNStageIntLLROutputS3xD(307)(1);
  VNStageIntLLRInputS3xD(131)(4) <= CNStageIntLLROutputS3xD(307)(2);
  VNStageIntLLRInputS3xD(228)(5) <= CNStageIntLLROutputS3xD(307)(3);
  VNStageIntLLRInputS3xD(309)(5) <= CNStageIntLLROutputS3xD(307)(4);
  VNStageIntLLRInputS3xD(344)(5) <= CNStageIntLLROutputS3xD(307)(5);
  VNStageIntLLRInputS3xD(62)(4) <= CNStageIntLLROutputS3xD(308)(0);
  VNStageIntLLRInputS3xD(98)(4) <= CNStageIntLLROutputS3xD(308)(1);
  VNStageIntLLRInputS3xD(179)(5) <= CNStageIntLLROutputS3xD(308)(2);
  VNStageIntLLRInputS3xD(214)(5) <= CNStageIntLLROutputS3xD(308)(3);
  VNStageIntLLRInputS3xD(288)(5) <= CNStageIntLLROutputS3xD(308)(4);
  VNStageIntLLRInputS3xD(366)(5) <= CNStageIntLLROutputS3xD(308)(5);
  VNStageIntLLRInputS3xD(61)(4) <= CNStageIntLLROutputS3xD(309)(0);
  VNStageIntLLRInputS3xD(114)(5) <= CNStageIntLLROutputS3xD(309)(1);
  VNStageIntLLRInputS3xD(149)(5) <= CNStageIntLLROutputS3xD(309)(2);
  VNStageIntLLRInputS3xD(223)(5) <= CNStageIntLLROutputS3xD(309)(3);
  VNStageIntLLRInputS3xD(301)(5) <= CNStageIntLLROutputS3xD(309)(4);
  VNStageIntLLRInputS3xD(345)(4) <= CNStageIntLLROutputS3xD(309)(5);
  VNStageIntLLRInputS3xD(60)(4) <= CNStageIntLLROutputS3xD(310)(0);
  VNStageIntLLRInputS3xD(84)(4) <= CNStageIntLLROutputS3xD(310)(1);
  VNStageIntLLRInputS3xD(158)(5) <= CNStageIntLLROutputS3xD(310)(2);
  VNStageIntLLRInputS3xD(236)(5) <= CNStageIntLLROutputS3xD(310)(3);
  VNStageIntLLRInputS3xD(280)(5) <= CNStageIntLLROutputS3xD(310)(4);
  VNStageIntLLRInputS3xD(373)(3) <= CNStageIntLLROutputS3xD(310)(5);
  VNStageIntLLRInputS3xD(59)(3) <= CNStageIntLLROutputS3xD(311)(0);
  VNStageIntLLRInputS3xD(93)(5) <= CNStageIntLLROutputS3xD(311)(1);
  VNStageIntLLRInputS3xD(171)(3) <= CNStageIntLLROutputS3xD(311)(2);
  VNStageIntLLRInputS3xD(215)(5) <= CNStageIntLLROutputS3xD(311)(3);
  VNStageIntLLRInputS3xD(308)(3) <= CNStageIntLLROutputS3xD(311)(4);
  VNStageIntLLRInputS3xD(375)(4) <= CNStageIntLLROutputS3xD(311)(5);
  VNStageIntLLRInputS3xD(58)(3) <= CNStageIntLLROutputS3xD(312)(0);
  VNStageIntLLRInputS3xD(106)(4) <= CNStageIntLLROutputS3xD(312)(1);
  VNStageIntLLRInputS3xD(150)(4) <= CNStageIntLLROutputS3xD(312)(2);
  VNStageIntLLRInputS3xD(243)(5) <= CNStageIntLLROutputS3xD(312)(3);
  VNStageIntLLRInputS3xD(310)(4) <= CNStageIntLLROutputS3xD(312)(4);
  VNStageIntLLRInputS3xD(357)(5) <= CNStageIntLLROutputS3xD(312)(5);
  VNStageIntLLRInputS3xD(57)(4) <= CNStageIntLLROutputS3xD(313)(0);
  VNStageIntLLRInputS3xD(85)(4) <= CNStageIntLLROutputS3xD(313)(1);
  VNStageIntLLRInputS3xD(178)(4) <= CNStageIntLLROutputS3xD(313)(2);
  VNStageIntLLRInputS3xD(245)(5) <= CNStageIntLLROutputS3xD(313)(3);
  VNStageIntLLRInputS3xD(292)(5) <= CNStageIntLLROutputS3xD(313)(4);
  VNStageIntLLRInputS3xD(364)(5) <= CNStageIntLLROutputS3xD(313)(5);
  VNStageIntLLRInputS3xD(56)(5) <= CNStageIntLLROutputS3xD(314)(0);
  VNStageIntLLRInputS3xD(113)(5) <= CNStageIntLLROutputS3xD(314)(1);
  VNStageIntLLRInputS3xD(180)(3) <= CNStageIntLLROutputS3xD(314)(2);
  VNStageIntLLRInputS3xD(227)(5) <= CNStageIntLLROutputS3xD(314)(3);
  VNStageIntLLRInputS3xD(299)(4) <= CNStageIntLLROutputS3xD(314)(4);
  VNStageIntLLRInputS3xD(328)(3) <= CNStageIntLLROutputS3xD(314)(5);
  VNStageIntLLRInputS3xD(55)(5) <= CNStageIntLLROutputS3xD(315)(0);
  VNStageIntLLRInputS3xD(115)(5) <= CNStageIntLLROutputS3xD(315)(1);
  VNStageIntLLRInputS3xD(162)(5) <= CNStageIntLLROutputS3xD(315)(2);
  VNStageIntLLRInputS3xD(234)(5) <= CNStageIntLLROutputS3xD(315)(3);
  VNStageIntLLRInputS3xD(263)(5) <= CNStageIntLLROutputS3xD(315)(4);
  VNStageIntLLRInputS3xD(379)(3) <= CNStageIntLLROutputS3xD(315)(5);
  VNStageIntLLRInputS3xD(54)(4) <= CNStageIntLLROutputS3xD(316)(0);
  VNStageIntLLRInputS3xD(97)(5) <= CNStageIntLLROutputS3xD(316)(1);
  VNStageIntLLRInputS3xD(169)(5) <= CNStageIntLLROutputS3xD(316)(2);
  VNStageIntLLRInputS3xD(198)(5) <= CNStageIntLLROutputS3xD(316)(3);
  VNStageIntLLRInputS3xD(314)(2) <= CNStageIntLLROutputS3xD(316)(4);
  VNStageIntLLRInputS3xD(322)(4) <= CNStageIntLLROutputS3xD(316)(5);
  VNStageIntLLRInputS3xD(53)(4) <= CNStageIntLLROutputS3xD(317)(0);
  VNStageIntLLRInputS3xD(104)(5) <= CNStageIntLLROutputS3xD(317)(1);
  VNStageIntLLRInputS3xD(133)(3) <= CNStageIntLLROutputS3xD(317)(2);
  VNStageIntLLRInputS3xD(249)(3) <= CNStageIntLLROutputS3xD(317)(3);
  VNStageIntLLRInputS3xD(257)(5) <= CNStageIntLLROutputS3xD(317)(4);
  VNStageIntLLRInputS3xD(380)(4) <= CNStageIntLLROutputS3xD(317)(5);
  VNStageIntLLRInputS3xD(52)(3) <= CNStageIntLLROutputS3xD(318)(0);
  VNStageIntLLRInputS3xD(68)(4) <= CNStageIntLLROutputS3xD(318)(1);
  VNStageIntLLRInputS3xD(184)(5) <= CNStageIntLLROutputS3xD(318)(2);
  VNStageIntLLRInputS3xD(255)(5) <= CNStageIntLLROutputS3xD(318)(3);
  VNStageIntLLRInputS3xD(315)(4) <= CNStageIntLLROutputS3xD(318)(4);
  VNStageIntLLRInputS3xD(327)(5) <= CNStageIntLLROutputS3xD(318)(5);
  VNStageIntLLRInputS3xD(51)(4) <= CNStageIntLLROutputS3xD(319)(0);
  VNStageIntLLRInputS3xD(119)(4) <= CNStageIntLLROutputS3xD(319)(1);
  VNStageIntLLRInputS3xD(190)(3) <= CNStageIntLLROutputS3xD(319)(2);
  VNStageIntLLRInputS3xD(250)(3) <= CNStageIntLLROutputS3xD(319)(3);
  VNStageIntLLRInputS3xD(262)(4) <= CNStageIntLLROutputS3xD(319)(4);
  VNStageIntLLRInputS3xD(349)(4) <= CNStageIntLLROutputS3xD(319)(5);
  VNStageIntLLRInputS3xD(50)(5) <= CNStageIntLLROutputS3xD(320)(0);
  VNStageIntLLRInputS3xD(125)(2) <= CNStageIntLLROutputS3xD(320)(1);
  VNStageIntLLRInputS3xD(185)(2) <= CNStageIntLLROutputS3xD(320)(2);
  VNStageIntLLRInputS3xD(197)(5) <= CNStageIntLLROutputS3xD(320)(3);
  VNStageIntLLRInputS3xD(284)(5) <= CNStageIntLLROutputS3xD(320)(4);
  VNStageIntLLRInputS3xD(367)(5) <= CNStageIntLLROutputS3xD(320)(5);
  VNStageIntLLRInputS3xD(49)(5) <= CNStageIntLLROutputS3xD(321)(0);
  VNStageIntLLRInputS3xD(120)(2) <= CNStageIntLLROutputS3xD(321)(1);
  VNStageIntLLRInputS3xD(132)(4) <= CNStageIntLLROutputS3xD(321)(2);
  VNStageIntLLRInputS3xD(219)(4) <= CNStageIntLLROutputS3xD(321)(3);
  VNStageIntLLRInputS3xD(302)(5) <= CNStageIntLLROutputS3xD(321)(4);
  VNStageIntLLRInputS3xD(352)(5) <= CNStageIntLLROutputS3xD(321)(5);
  VNStageIntLLRInputS3xD(48)(2) <= CNStageIntLLROutputS3xD(322)(0);
  VNStageIntLLRInputS3xD(67)(2) <= CNStageIntLLROutputS3xD(322)(1);
  VNStageIntLLRInputS3xD(154)(4) <= CNStageIntLLROutputS3xD(322)(2);
  VNStageIntLLRInputS3xD(237)(4) <= CNStageIntLLROutputS3xD(322)(3);
  VNStageIntLLRInputS3xD(287)(5) <= CNStageIntLLROutputS3xD(322)(4);
  VNStageIntLLRInputS3xD(339)(5) <= CNStageIntLLROutputS3xD(322)(5);
  VNStageIntLLRInputS3xD(46)(5) <= CNStageIntLLROutputS3xD(323)(0);
  VNStageIntLLRInputS3xD(107)(4) <= CNStageIntLLROutputS3xD(323)(1);
  VNStageIntLLRInputS3xD(157)(4) <= CNStageIntLLROutputS3xD(323)(2);
  VNStageIntLLRInputS3xD(209)(4) <= CNStageIntLLROutputS3xD(323)(3);
  VNStageIntLLRInputS3xD(305)(5) <= CNStageIntLLROutputS3xD(323)(4);
  VNStageIntLLRInputS3xD(382)(4) <= CNStageIntLLROutputS3xD(323)(5);
  VNStageIntLLRInputS3xD(45)(5) <= CNStageIntLLROutputS3xD(324)(0);
  VNStageIntLLRInputS3xD(92)(5) <= CNStageIntLLROutputS3xD(324)(1);
  VNStageIntLLRInputS3xD(144)(5) <= CNStageIntLLROutputS3xD(324)(2);
  VNStageIntLLRInputS3xD(240)(5) <= CNStageIntLLROutputS3xD(324)(3);
  VNStageIntLLRInputS3xD(317)(2) <= CNStageIntLLROutputS3xD(324)(4);
  VNStageIntLLRInputS3xD(333)(4) <= CNStageIntLLROutputS3xD(324)(5);
  VNStageIntLLRInputS3xD(44)(5) <= CNStageIntLLROutputS3xD(325)(0);
  VNStageIntLLRInputS3xD(79)(4) <= CNStageIntLLROutputS3xD(325)(1);
  VNStageIntLLRInputS3xD(175)(5) <= CNStageIntLLROutputS3xD(325)(2);
  VNStageIntLLRInputS3xD(252)(4) <= CNStageIntLLROutputS3xD(325)(3);
  VNStageIntLLRInputS3xD(268)(5) <= CNStageIntLLROutputS3xD(325)(4);
  VNStageIntLLRInputS3xD(377)(3) <= CNStageIntLLROutputS3xD(325)(5);
  VNStageIntLLRInputS3xD(43)(4) <= CNStageIntLLROutputS3xD(326)(0);
  VNStageIntLLRInputS3xD(110)(5) <= CNStageIntLLROutputS3xD(326)(1);
  VNStageIntLLRInputS3xD(187)(4) <= CNStageIntLLROutputS3xD(326)(2);
  VNStageIntLLRInputS3xD(203)(5) <= CNStageIntLLROutputS3xD(326)(3);
  VNStageIntLLRInputS3xD(312)(4) <= CNStageIntLLROutputS3xD(326)(4);
  VNStageIntLLRInputS3xD(354)(4) <= CNStageIntLLROutputS3xD(326)(5);
  VNStageIntLLRInputS3xD(42)(5) <= CNStageIntLLROutputS3xD(327)(0);
  VNStageIntLLRInputS3xD(122)(4) <= CNStageIntLLROutputS3xD(327)(1);
  VNStageIntLLRInputS3xD(138)(5) <= CNStageIntLLROutputS3xD(327)(2);
  VNStageIntLLRInputS3xD(247)(5) <= CNStageIntLLROutputS3xD(327)(3);
  VNStageIntLLRInputS3xD(289)(5) <= CNStageIntLLROutputS3xD(327)(4);
  VNStageIntLLRInputS3xD(343)(5) <= CNStageIntLLROutputS3xD(327)(5);
  VNStageIntLLRInputS3xD(41)(5) <= CNStageIntLLROutputS3xD(328)(0);
  VNStageIntLLRInputS3xD(73)(4) <= CNStageIntLLROutputS3xD(328)(1);
  VNStageIntLLRInputS3xD(182)(5) <= CNStageIntLLROutputS3xD(328)(2);
  VNStageIntLLRInputS3xD(224)(5) <= CNStageIntLLROutputS3xD(328)(3);
  VNStageIntLLRInputS3xD(278)(4) <= CNStageIntLLROutputS3xD(328)(4);
  VNStageIntLLRInputS3xD(347)(5) <= CNStageIntLLROutputS3xD(328)(5);
  VNStageIntLLRInputS3xD(39)(5) <= CNStageIntLLROutputS3xD(329)(0);
  VNStageIntLLRInputS3xD(94)(3) <= CNStageIntLLROutputS3xD(329)(1);
  VNStageIntLLRInputS3xD(148)(5) <= CNStageIntLLROutputS3xD(329)(2);
  VNStageIntLLRInputS3xD(217)(5) <= CNStageIntLLROutputS3xD(329)(3);
  VNStageIntLLRInputS3xD(275)(4) <= CNStageIntLLROutputS3xD(329)(4);
  VNStageIntLLRInputS3xD(351)(4) <= CNStageIntLLROutputS3xD(329)(5);
  VNStageIntLLRInputS3xD(38)(5) <= CNStageIntLLROutputS3xD(330)(0);
  VNStageIntLLRInputS3xD(83)(5) <= CNStageIntLLROutputS3xD(330)(1);
  VNStageIntLLRInputS3xD(152)(5) <= CNStageIntLLROutputS3xD(330)(2);
  VNStageIntLLRInputS3xD(210)(5) <= CNStageIntLLROutputS3xD(330)(3);
  VNStageIntLLRInputS3xD(286)(5) <= CNStageIntLLROutputS3xD(330)(4);
  VNStageIntLLRInputS3xD(323)(4) <= CNStageIntLLROutputS3xD(330)(5);
  VNStageIntLLRInputS3xD(37)(5) <= CNStageIntLLROutputS3xD(331)(0);
  VNStageIntLLRInputS3xD(87)(5) <= CNStageIntLLROutputS3xD(331)(1);
  VNStageIntLLRInputS3xD(145)(5) <= CNStageIntLLROutputS3xD(331)(2);
  VNStageIntLLRInputS3xD(221)(5) <= CNStageIntLLROutputS3xD(331)(3);
  VNStageIntLLRInputS3xD(258)(2) <= CNStageIntLLROutputS3xD(331)(4);
  VNStageIntLLRInputS3xD(378)(4) <= CNStageIntLLROutputS3xD(331)(5);
  VNStageIntLLRInputS3xD(0)(5) <= CNStageIntLLROutputS3xD(332)(0);
  VNStageIntLLRInputS3xD(76)(5) <= CNStageIntLLROutputS3xD(332)(1);
  VNStageIntLLRInputS3xD(141)(3) <= CNStageIntLLROutputS3xD(332)(2);
  VNStageIntLLRInputS3xD(206)(3) <= CNStageIntLLROutputS3xD(332)(3);
  VNStageIntLLRInputS3xD(271)(4) <= CNStageIntLLROutputS3xD(332)(4);
  VNStageIntLLRInputS3xD(336)(4) <= CNStageIntLLROutputS3xD(332)(5);
  VNStageIntLLRInputS3xD(28)(5) <= CNStageIntLLROutputS3xD(333)(0);
  VNStageIntLLRInputS3xD(106)(5) <= CNStageIntLLROutputS3xD(333)(1);
  VNStageIntLLRInputS3xD(144)(6) <= CNStageIntLLROutputS3xD(333)(2);
  VNStageIntLLRInputS3xD(193)(4) <= CNStageIntLLROutputS3xD(333)(3);
  VNStageIntLLRInputS3xD(261)(5) <= CNStageIntLLROutputS3xD(333)(4);
  VNStageIntLLRInputS3xD(367)(6) <= CNStageIntLLROutputS3xD(333)(5);
  VNStageIntLLRInputS3xD(26)(6) <= CNStageIntLLROutputS3xD(334)(0);
  VNStageIntLLRInputS3xD(126)(5) <= CNStageIntLLROutputS3xD(334)(1);
  VNStageIntLLRInputS3xD(131)(5) <= CNStageIntLLROutputS3xD(334)(2);
  VNStageIntLLRInputS3xD(237)(5) <= CNStageIntLLROutputS3xD(334)(3);
  VNStageIntLLRInputS3xD(277)(6) <= CNStageIntLLROutputS3xD(334)(4);
  VNStageIntLLRInputS3xD(340)(5) <= CNStageIntLLROutputS3xD(334)(5);
  VNStageIntLLRInputS3xD(24)(6) <= CNStageIntLLROutputS3xD(335)(0);
  VNStageIntLLRInputS3xD(107)(5) <= CNStageIntLLROutputS3xD(335)(1);
  VNStageIntLLRInputS3xD(147)(6) <= CNStageIntLLROutputS3xD(335)(2);
  VNStageIntLLRInputS3xD(210)(6) <= CNStageIntLLROutputS3xD(335)(3);
  VNStageIntLLRInputS3xD(300)(5) <= CNStageIntLLROutputS3xD(335)(4);
  VNStageIntLLRInputS3xD(373)(4) <= CNStageIntLLROutputS3xD(335)(5);
  VNStageIntLLRInputS3xD(23)(6) <= CNStageIntLLROutputS3xD(336)(0);
  VNStageIntLLRInputS3xD(82)(6) <= CNStageIntLLROutputS3xD(336)(1);
  VNStageIntLLRInputS3xD(145)(6) <= CNStageIntLLROutputS3xD(336)(2);
  VNStageIntLLRInputS3xD(235)(4) <= CNStageIntLLROutputS3xD(336)(3);
  VNStageIntLLRInputS3xD(308)(4) <= CNStageIntLLROutputS3xD(336)(4);
  VNStageIntLLRInputS3xD(353)(5) <= CNStageIntLLROutputS3xD(336)(5);
  VNStageIntLLRInputS3xD(22)(6) <= CNStageIntLLROutputS3xD(337)(0);
  VNStageIntLLRInputS3xD(80)(5) <= CNStageIntLLROutputS3xD(337)(1);
  VNStageIntLLRInputS3xD(170)(4) <= CNStageIntLLROutputS3xD(337)(2);
  VNStageIntLLRInputS3xD(243)(6) <= CNStageIntLLROutputS3xD(337)(3);
  VNStageIntLLRInputS3xD(288)(6) <= CNStageIntLLROutputS3xD(337)(4);
  VNStageIntLLRInputS3xD(347)(6) <= CNStageIntLLROutputS3xD(337)(5);
  VNStageIntLLRInputS3xD(21)(6) <= CNStageIntLLROutputS3xD(338)(0);
  VNStageIntLLRInputS3xD(105)(5) <= CNStageIntLLROutputS3xD(338)(1);
  VNStageIntLLRInputS3xD(178)(5) <= CNStageIntLLROutputS3xD(338)(2);
  VNStageIntLLRInputS3xD(223)(6) <= CNStageIntLLROutputS3xD(338)(3);
  VNStageIntLLRInputS3xD(282)(5) <= CNStageIntLLROutputS3xD(338)(4);
  VNStageIntLLRInputS3xD(320)(4) <= CNStageIntLLROutputS3xD(338)(5);
  VNStageIntLLRInputS3xD(20)(4) <= CNStageIntLLROutputS3xD(339)(0);
  VNStageIntLLRInputS3xD(113)(6) <= CNStageIntLLROutputS3xD(339)(1);
  VNStageIntLLRInputS3xD(158)(6) <= CNStageIntLLROutputS3xD(339)(2);
  VNStageIntLLRInputS3xD(217)(6) <= CNStageIntLLROutputS3xD(339)(3);
  VNStageIntLLRInputS3xD(256)(5) <= CNStageIntLLROutputS3xD(339)(4);
  VNStageIntLLRInputS3xD(346)(6) <= CNStageIntLLROutputS3xD(339)(5);
  VNStageIntLLRInputS3xD(19)(4) <= CNStageIntLLROutputS3xD(340)(0);
  VNStageIntLLRInputS3xD(93)(6) <= CNStageIntLLROutputS3xD(340)(1);
  VNStageIntLLRInputS3xD(152)(6) <= CNStageIntLLROutputS3xD(340)(2);
  VNStageIntLLRInputS3xD(192)(6) <= CNStageIntLLROutputS3xD(340)(3);
  VNStageIntLLRInputS3xD(281)(6) <= CNStageIntLLROutputS3xD(340)(4);
  VNStageIntLLRInputS3xD(351)(5) <= CNStageIntLLROutputS3xD(340)(5);
  VNStageIntLLRInputS3xD(18)(6) <= CNStageIntLLROutputS3xD(341)(0);
  VNStageIntLLRInputS3xD(87)(6) <= CNStageIntLLROutputS3xD(341)(1);
  VNStageIntLLRInputS3xD(128)(6) <= CNStageIntLLROutputS3xD(341)(2);
  VNStageIntLLRInputS3xD(216)(6) <= CNStageIntLLROutputS3xD(341)(3);
  VNStageIntLLRInputS3xD(286)(6) <= CNStageIntLLROutputS3xD(341)(4);
  VNStageIntLLRInputS3xD(370)(4) <= CNStageIntLLROutputS3xD(341)(5);
  VNStageIntLLRInputS3xD(17)(6) <= CNStageIntLLROutputS3xD(342)(0);
  VNStageIntLLRInputS3xD(64)(5) <= CNStageIntLLROutputS3xD(342)(1);
  VNStageIntLLRInputS3xD(151)(5) <= CNStageIntLLROutputS3xD(342)(2);
  VNStageIntLLRInputS3xD(221)(6) <= CNStageIntLLROutputS3xD(342)(3);
  VNStageIntLLRInputS3xD(305)(6) <= CNStageIntLLROutputS3xD(342)(4);
  VNStageIntLLRInputS3xD(361)(6) <= CNStageIntLLROutputS3xD(342)(5);
  VNStageIntLLRInputS3xD(16)(5) <= CNStageIntLLROutputS3xD(343)(0);
  VNStageIntLLRInputS3xD(86)(3) <= CNStageIntLLROutputS3xD(343)(1);
  VNStageIntLLRInputS3xD(156)(3) <= CNStageIntLLROutputS3xD(343)(2);
  VNStageIntLLRInputS3xD(240)(6) <= CNStageIntLLROutputS3xD(343)(3);
  VNStageIntLLRInputS3xD(296)(5) <= CNStageIntLLROutputS3xD(343)(4);
  VNStageIntLLRInputS3xD(335)(6) <= CNStageIntLLROutputS3xD(343)(5);
  VNStageIntLLRInputS3xD(15)(6) <= CNStageIntLLROutputS3xD(344)(0);
  VNStageIntLLRInputS3xD(91)(6) <= CNStageIntLLROutputS3xD(344)(1);
  VNStageIntLLRInputS3xD(175)(6) <= CNStageIntLLROutputS3xD(344)(2);
  VNStageIntLLRInputS3xD(231)(5) <= CNStageIntLLROutputS3xD(344)(3);
  VNStageIntLLRInputS3xD(270)(6) <= CNStageIntLLROutputS3xD(344)(4);
  VNStageIntLLRInputS3xD(336)(5) <= CNStageIntLLROutputS3xD(344)(5);
  VNStageIntLLRInputS3xD(14)(6) <= CNStageIntLLROutputS3xD(345)(0);
  VNStageIntLLRInputS3xD(110)(6) <= CNStageIntLLROutputS3xD(345)(1);
  VNStageIntLLRInputS3xD(166)(5) <= CNStageIntLLROutputS3xD(345)(2);
  VNStageIntLLRInputS3xD(205)(2) <= CNStageIntLLROutputS3xD(345)(3);
  VNStageIntLLRInputS3xD(271)(5) <= CNStageIntLLROutputS3xD(345)(4);
  VNStageIntLLRInputS3xD(360)(6) <= CNStageIntLLROutputS3xD(345)(5);
  VNStageIntLLRInputS3xD(13)(5) <= CNStageIntLLROutputS3xD(346)(0);
  VNStageIntLLRInputS3xD(101)(6) <= CNStageIntLLROutputS3xD(346)(1);
  VNStageIntLLRInputS3xD(140)(6) <= CNStageIntLLROutputS3xD(346)(2);
  VNStageIntLLRInputS3xD(206)(4) <= CNStageIntLLROutputS3xD(346)(3);
  VNStageIntLLRInputS3xD(295)(4) <= CNStageIntLLROutputS3xD(346)(4);
  VNStageIntLLRInputS3xD(381)(5) <= CNStageIntLLROutputS3xD(346)(5);
  VNStageIntLLRInputS3xD(12)(6) <= CNStageIntLLROutputS3xD(347)(0);
  VNStageIntLLRInputS3xD(75)(6) <= CNStageIntLLROutputS3xD(347)(1);
  VNStageIntLLRInputS3xD(141)(4) <= CNStageIntLLROutputS3xD(347)(2);
  VNStageIntLLRInputS3xD(230)(5) <= CNStageIntLLROutputS3xD(347)(3);
  VNStageIntLLRInputS3xD(316)(4) <= CNStageIntLLROutputS3xD(347)(4);
  VNStageIntLLRInputS3xD(377)(4) <= CNStageIntLLROutputS3xD(347)(5);
  VNStageIntLLRInputS3xD(11)(5) <= CNStageIntLLROutputS3xD(348)(0);
  VNStageIntLLRInputS3xD(76)(6) <= CNStageIntLLROutputS3xD(348)(1);
  VNStageIntLLRInputS3xD(165)(5) <= CNStageIntLLROutputS3xD(348)(2);
  VNStageIntLLRInputS3xD(251)(4) <= CNStageIntLLROutputS3xD(348)(3);
  VNStageIntLLRInputS3xD(312)(5) <= CNStageIntLLROutputS3xD(348)(4);
  VNStageIntLLRInputS3xD(329)(6) <= CNStageIntLLROutputS3xD(348)(5);
  VNStageIntLLRInputS3xD(10)(4) <= CNStageIntLLROutputS3xD(349)(0);
  VNStageIntLLRInputS3xD(100)(6) <= CNStageIntLLROutputS3xD(349)(1);
  VNStageIntLLRInputS3xD(186)(5) <= CNStageIntLLROutputS3xD(349)(2);
  VNStageIntLLRInputS3xD(247)(6) <= CNStageIntLLROutputS3xD(349)(3);
  VNStageIntLLRInputS3xD(264)(6) <= CNStageIntLLROutputS3xD(349)(4);
  VNStageIntLLRInputS3xD(355)(6) <= CNStageIntLLROutputS3xD(349)(5);
  VNStageIntLLRInputS3xD(9)(6) <= CNStageIntLLROutputS3xD(350)(0);
  VNStageIntLLRInputS3xD(121)(5) <= CNStageIntLLROutputS3xD(350)(1);
  VNStageIntLLRInputS3xD(182)(6) <= CNStageIntLLROutputS3xD(350)(2);
  VNStageIntLLRInputS3xD(199)(6) <= CNStageIntLLROutputS3xD(350)(3);
  VNStageIntLLRInputS3xD(290)(5) <= CNStageIntLLROutputS3xD(350)(4);
  VNStageIntLLRInputS3xD(331)(4) <= CNStageIntLLROutputS3xD(350)(5);
  VNStageIntLLRInputS3xD(7)(6) <= CNStageIntLLROutputS3xD(351)(0);
  VNStageIntLLRInputS3xD(69)(6) <= CNStageIntLLROutputS3xD(351)(1);
  VNStageIntLLRInputS3xD(160)(6) <= CNStageIntLLROutputS3xD(351)(2);
  VNStageIntLLRInputS3xD(201)(5) <= CNStageIntLLROutputS3xD(351)(3);
  VNStageIntLLRInputS3xD(298)(6) <= CNStageIntLLROutputS3xD(351)(4);
  VNStageIntLLRInputS3xD(379)(4) <= CNStageIntLLROutputS3xD(351)(5);
  VNStageIntLLRInputS3xD(6)(6) <= CNStageIntLLROutputS3xD(352)(0);
  VNStageIntLLRInputS3xD(95)(6) <= CNStageIntLLROutputS3xD(352)(1);
  VNStageIntLLRInputS3xD(136)(6) <= CNStageIntLLROutputS3xD(352)(2);
  VNStageIntLLRInputS3xD(233)(4) <= CNStageIntLLROutputS3xD(352)(3);
  VNStageIntLLRInputS3xD(314)(3) <= CNStageIntLLROutputS3xD(352)(4);
  VNStageIntLLRInputS3xD(349)(5) <= CNStageIntLLROutputS3xD(352)(5);
  VNStageIntLLRInputS3xD(5)(6) <= CNStageIntLLROutputS3xD(353)(0);
  VNStageIntLLRInputS3xD(71)(5) <= CNStageIntLLROutputS3xD(353)(1);
  VNStageIntLLRInputS3xD(168)(5) <= CNStageIntLLROutputS3xD(353)(2);
  VNStageIntLLRInputS3xD(249)(4) <= CNStageIntLLROutputS3xD(353)(3);
  VNStageIntLLRInputS3xD(284)(6) <= CNStageIntLLROutputS3xD(353)(4);
  VNStageIntLLRInputS3xD(358)(5) <= CNStageIntLLROutputS3xD(353)(5);
  VNStageIntLLRInputS3xD(4)(5) <= CNStageIntLLROutputS3xD(354)(0);
  VNStageIntLLRInputS3xD(103)(6) <= CNStageIntLLROutputS3xD(354)(1);
  VNStageIntLLRInputS3xD(184)(6) <= CNStageIntLLROutputS3xD(354)(2);
  VNStageIntLLRInputS3xD(219)(5) <= CNStageIntLLROutputS3xD(354)(3);
  VNStageIntLLRInputS3xD(293)(5) <= CNStageIntLLROutputS3xD(354)(4);
  VNStageIntLLRInputS3xD(371)(4) <= CNStageIntLLROutputS3xD(354)(5);
  VNStageIntLLRInputS3xD(2)(6) <= CNStageIntLLROutputS3xD(355)(0);
  VNStageIntLLRInputS3xD(89)(5) <= CNStageIntLLROutputS3xD(355)(1);
  VNStageIntLLRInputS3xD(163)(4) <= CNStageIntLLROutputS3xD(355)(2);
  VNStageIntLLRInputS3xD(241)(5) <= CNStageIntLLROutputS3xD(355)(3);
  VNStageIntLLRInputS3xD(285)(6) <= CNStageIntLLROutputS3xD(355)(4);
  VNStageIntLLRInputS3xD(378)(5) <= CNStageIntLLROutputS3xD(355)(5);
  VNStageIntLLRInputS3xD(1)(5) <= CNStageIntLLROutputS3xD(356)(0);
  VNStageIntLLRInputS3xD(98)(5) <= CNStageIntLLROutputS3xD(356)(1);
  VNStageIntLLRInputS3xD(176)(6) <= CNStageIntLLROutputS3xD(356)(2);
  VNStageIntLLRInputS3xD(220)(6) <= CNStageIntLLROutputS3xD(356)(3);
  VNStageIntLLRInputS3xD(313)(3) <= CNStageIntLLROutputS3xD(356)(4);
  VNStageIntLLRInputS3xD(380)(5) <= CNStageIntLLROutputS3xD(356)(5);
  VNStageIntLLRInputS3xD(63)(3) <= CNStageIntLLROutputS3xD(357)(0);
  VNStageIntLLRInputS3xD(111)(6) <= CNStageIntLLROutputS3xD(357)(1);
  VNStageIntLLRInputS3xD(155)(6) <= CNStageIntLLROutputS3xD(357)(2);
  VNStageIntLLRInputS3xD(248)(6) <= CNStageIntLLROutputS3xD(357)(3);
  VNStageIntLLRInputS3xD(315)(5) <= CNStageIntLLROutputS3xD(357)(4);
  VNStageIntLLRInputS3xD(362)(6) <= CNStageIntLLROutputS3xD(357)(5);
  VNStageIntLLRInputS3xD(62)(5) <= CNStageIntLLROutputS3xD(358)(0);
  VNStageIntLLRInputS3xD(90)(6) <= CNStageIntLLROutputS3xD(358)(1);
  VNStageIntLLRInputS3xD(183)(4) <= CNStageIntLLROutputS3xD(358)(2);
  VNStageIntLLRInputS3xD(250)(4) <= CNStageIntLLROutputS3xD(358)(3);
  VNStageIntLLRInputS3xD(297)(6) <= CNStageIntLLROutputS3xD(358)(4);
  VNStageIntLLRInputS3xD(369)(4) <= CNStageIntLLROutputS3xD(358)(5);
  VNStageIntLLRInputS3xD(61)(5) <= CNStageIntLLROutputS3xD(359)(0);
  VNStageIntLLRInputS3xD(118)(5) <= CNStageIntLLROutputS3xD(359)(1);
  VNStageIntLLRInputS3xD(185)(3) <= CNStageIntLLROutputS3xD(359)(2);
  VNStageIntLLRInputS3xD(232)(5) <= CNStageIntLLROutputS3xD(359)(3);
  VNStageIntLLRInputS3xD(304)(6) <= CNStageIntLLROutputS3xD(359)(4);
  VNStageIntLLRInputS3xD(333)(5) <= CNStageIntLLROutputS3xD(359)(5);
  VNStageIntLLRInputS3xD(60)(5) <= CNStageIntLLROutputS3xD(360)(0);
  VNStageIntLLRInputS3xD(120)(3) <= CNStageIntLLROutputS3xD(360)(1);
  VNStageIntLLRInputS3xD(167)(6) <= CNStageIntLLROutputS3xD(360)(2);
  VNStageIntLLRInputS3xD(239)(6) <= CNStageIntLLROutputS3xD(360)(3);
  VNStageIntLLRInputS3xD(268)(6) <= CNStageIntLLROutputS3xD(360)(4);
  VNStageIntLLRInputS3xD(321)(6) <= CNStageIntLLROutputS3xD(360)(5);
  VNStageIntLLRInputS3xD(59)(4) <= CNStageIntLLROutputS3xD(361)(0);
  VNStageIntLLRInputS3xD(102)(5) <= CNStageIntLLROutputS3xD(361)(1);
  VNStageIntLLRInputS3xD(174)(4) <= CNStageIntLLROutputS3xD(361)(2);
  VNStageIntLLRInputS3xD(203)(6) <= CNStageIntLLROutputS3xD(361)(3);
  VNStageIntLLRInputS3xD(319)(6) <= CNStageIntLLROutputS3xD(361)(4);
  VNStageIntLLRInputS3xD(327)(6) <= CNStageIntLLROutputS3xD(361)(5);
  VNStageIntLLRInputS3xD(58)(4) <= CNStageIntLLROutputS3xD(362)(0);
  VNStageIntLLRInputS3xD(109)(5) <= CNStageIntLLROutputS3xD(362)(1);
  VNStageIntLLRInputS3xD(138)(6) <= CNStageIntLLROutputS3xD(362)(2);
  VNStageIntLLRInputS3xD(254)(4) <= CNStageIntLLROutputS3xD(362)(3);
  VNStageIntLLRInputS3xD(262)(5) <= CNStageIntLLROutputS3xD(362)(4);
  VNStageIntLLRInputS3xD(322)(5) <= CNStageIntLLROutputS3xD(362)(5);
  VNStageIntLLRInputS3xD(57)(5) <= CNStageIntLLROutputS3xD(363)(0);
  VNStageIntLLRInputS3xD(73)(5) <= CNStageIntLLROutputS3xD(363)(1);
  VNStageIntLLRInputS3xD(189)(5) <= CNStageIntLLROutputS3xD(363)(2);
  VNStageIntLLRInputS3xD(197)(6) <= CNStageIntLLROutputS3xD(363)(3);
  VNStageIntLLRInputS3xD(257)(6) <= CNStageIntLLROutputS3xD(363)(4);
  VNStageIntLLRInputS3xD(332)(5) <= CNStageIntLLROutputS3xD(363)(5);
  VNStageIntLLRInputS3xD(56)(6) <= CNStageIntLLROutputS3xD(364)(0);
  VNStageIntLLRInputS3xD(124)(4) <= CNStageIntLLROutputS3xD(364)(1);
  VNStageIntLLRInputS3xD(132)(5) <= CNStageIntLLROutputS3xD(364)(2);
  VNStageIntLLRInputS3xD(255)(6) <= CNStageIntLLROutputS3xD(364)(3);
  VNStageIntLLRInputS3xD(267)(6) <= CNStageIntLLROutputS3xD(364)(4);
  VNStageIntLLRInputS3xD(354)(5) <= CNStageIntLLROutputS3xD(364)(5);
  VNStageIntLLRInputS3xD(55)(6) <= CNStageIntLLROutputS3xD(365)(0);
  VNStageIntLLRInputS3xD(67)(3) <= CNStageIntLLROutputS3xD(365)(1);
  VNStageIntLLRInputS3xD(190)(4) <= CNStageIntLLROutputS3xD(365)(2);
  VNStageIntLLRInputS3xD(202)(5) <= CNStageIntLLROutputS3xD(365)(3);
  VNStageIntLLRInputS3xD(289)(6) <= CNStageIntLLROutputS3xD(365)(4);
  VNStageIntLLRInputS3xD(372)(5) <= CNStageIntLLROutputS3xD(365)(5);
  VNStageIntLLRInputS3xD(54)(5) <= CNStageIntLLROutputS3xD(366)(0);
  VNStageIntLLRInputS3xD(125)(3) <= CNStageIntLLROutputS3xD(366)(1);
  VNStageIntLLRInputS3xD(137)(6) <= CNStageIntLLROutputS3xD(366)(2);
  VNStageIntLLRInputS3xD(224)(6) <= CNStageIntLLROutputS3xD(366)(3);
  VNStageIntLLRInputS3xD(307)(6) <= CNStageIntLLROutputS3xD(366)(4);
  VNStageIntLLRInputS3xD(357)(6) <= CNStageIntLLROutputS3xD(366)(5);
  VNStageIntLLRInputS3xD(53)(5) <= CNStageIntLLROutputS3xD(367)(0);
  VNStageIntLLRInputS3xD(72)(5) <= CNStageIntLLROutputS3xD(367)(1);
  VNStageIntLLRInputS3xD(159)(4) <= CNStageIntLLROutputS3xD(367)(2);
  VNStageIntLLRInputS3xD(242)(6) <= CNStageIntLLROutputS3xD(367)(3);
  VNStageIntLLRInputS3xD(292)(6) <= CNStageIntLLROutputS3xD(367)(4);
  VNStageIntLLRInputS3xD(344)(6) <= CNStageIntLLROutputS3xD(367)(5);
  VNStageIntLLRInputS3xD(52)(4) <= CNStageIntLLROutputS3xD(368)(0);
  VNStageIntLLRInputS3xD(94)(4) <= CNStageIntLLROutputS3xD(368)(1);
  VNStageIntLLRInputS3xD(177)(6) <= CNStageIntLLROutputS3xD(368)(2);
  VNStageIntLLRInputS3xD(227)(6) <= CNStageIntLLROutputS3xD(368)(3);
  VNStageIntLLRInputS3xD(279)(5) <= CNStageIntLLROutputS3xD(368)(4);
  VNStageIntLLRInputS3xD(375)(5) <= CNStageIntLLROutputS3xD(368)(5);
  VNStageIntLLRInputS3xD(51)(5) <= CNStageIntLLROutputS3xD(369)(0);
  VNStageIntLLRInputS3xD(112)(6) <= CNStageIntLLROutputS3xD(369)(1);
  VNStageIntLLRInputS3xD(162)(6) <= CNStageIntLLROutputS3xD(369)(2);
  VNStageIntLLRInputS3xD(214)(6) <= CNStageIntLLROutputS3xD(369)(3);
  VNStageIntLLRInputS3xD(310)(5) <= CNStageIntLLROutputS3xD(369)(4);
  VNStageIntLLRInputS3xD(324)(6) <= CNStageIntLLROutputS3xD(369)(5);
  VNStageIntLLRInputS3xD(50)(6) <= CNStageIntLLROutputS3xD(370)(0);
  VNStageIntLLRInputS3xD(97)(6) <= CNStageIntLLROutputS3xD(370)(1);
  VNStageIntLLRInputS3xD(149)(6) <= CNStageIntLLROutputS3xD(370)(2);
  VNStageIntLLRInputS3xD(245)(6) <= CNStageIntLLROutputS3xD(370)(3);
  VNStageIntLLRInputS3xD(259)(4) <= CNStageIntLLROutputS3xD(370)(4);
  VNStageIntLLRInputS3xD(338)(4) <= CNStageIntLLROutputS3xD(370)(5);
  VNStageIntLLRInputS3xD(49)(6) <= CNStageIntLLROutputS3xD(371)(0);
  VNStageIntLLRInputS3xD(84)(5) <= CNStageIntLLROutputS3xD(371)(1);
  VNStageIntLLRInputS3xD(180)(4) <= CNStageIntLLROutputS3xD(371)(2);
  VNStageIntLLRInputS3xD(194)(6) <= CNStageIntLLROutputS3xD(371)(3);
  VNStageIntLLRInputS3xD(273)(5) <= CNStageIntLLROutputS3xD(371)(4);
  VNStageIntLLRInputS3xD(382)(5) <= CNStageIntLLROutputS3xD(371)(5);
  VNStageIntLLRInputS3xD(48)(3) <= CNStageIntLLROutputS3xD(372)(0);
  VNStageIntLLRInputS3xD(115)(6) <= CNStageIntLLROutputS3xD(372)(1);
  VNStageIntLLRInputS3xD(129)(6) <= CNStageIntLLROutputS3xD(372)(2);
  VNStageIntLLRInputS3xD(208)(5) <= CNStageIntLLROutputS3xD(372)(3);
  VNStageIntLLRInputS3xD(317)(3) <= CNStageIntLLROutputS3xD(372)(4);
  VNStageIntLLRInputS3xD(359)(6) <= CNStageIntLLROutputS3xD(372)(5);
  VNStageIntLLRInputS3xD(47)(3) <= CNStageIntLLROutputS3xD(373)(0);
  VNStageIntLLRInputS3xD(127)(6) <= CNStageIntLLROutputS3xD(373)(1);
  VNStageIntLLRInputS3xD(143)(6) <= CNStageIntLLROutputS3xD(373)(2);
  VNStageIntLLRInputS3xD(252)(5) <= CNStageIntLLROutputS3xD(373)(3);
  VNStageIntLLRInputS3xD(294)(6) <= CNStageIntLLROutputS3xD(373)(4);
  VNStageIntLLRInputS3xD(348)(6) <= CNStageIntLLROutputS3xD(373)(5);
  VNStageIntLLRInputS3xD(46)(6) <= CNStageIntLLROutputS3xD(374)(0);
  VNStageIntLLRInputS3xD(78)(6) <= CNStageIntLLROutputS3xD(374)(1);
  VNStageIntLLRInputS3xD(187)(5) <= CNStageIntLLROutputS3xD(374)(2);
  VNStageIntLLRInputS3xD(229)(4) <= CNStageIntLLROutputS3xD(374)(3);
  VNStageIntLLRInputS3xD(283)(6) <= CNStageIntLLROutputS3xD(374)(4);
  VNStageIntLLRInputS3xD(352)(6) <= CNStageIntLLROutputS3xD(374)(5);
  VNStageIntLLRInputS3xD(45)(6) <= CNStageIntLLROutputS3xD(375)(0);
  VNStageIntLLRInputS3xD(122)(5) <= CNStageIntLLROutputS3xD(375)(1);
  VNStageIntLLRInputS3xD(164)(5) <= CNStageIntLLROutputS3xD(375)(2);
  VNStageIntLLRInputS3xD(218)(6) <= CNStageIntLLROutputS3xD(375)(3);
  VNStageIntLLRInputS3xD(287)(6) <= CNStageIntLLROutputS3xD(375)(4);
  VNStageIntLLRInputS3xD(345)(5) <= CNStageIntLLROutputS3xD(375)(5);
  VNStageIntLLRInputS3xD(44)(6) <= CNStageIntLLROutputS3xD(376)(0);
  VNStageIntLLRInputS3xD(99)(6) <= CNStageIntLLROutputS3xD(376)(1);
  VNStageIntLLRInputS3xD(153)(6) <= CNStageIntLLROutputS3xD(376)(2);
  VNStageIntLLRInputS3xD(222)(3) <= CNStageIntLLROutputS3xD(376)(3);
  VNStageIntLLRInputS3xD(280)(6) <= CNStageIntLLROutputS3xD(376)(4);
  VNStageIntLLRInputS3xD(356)(5) <= CNStageIntLLROutputS3xD(376)(5);
  VNStageIntLLRInputS3xD(43)(5) <= CNStageIntLLROutputS3xD(377)(0);
  VNStageIntLLRInputS3xD(88)(6) <= CNStageIntLLROutputS3xD(377)(1);
  VNStageIntLLRInputS3xD(157)(5) <= CNStageIntLLROutputS3xD(377)(2);
  VNStageIntLLRInputS3xD(215)(6) <= CNStageIntLLROutputS3xD(377)(3);
  VNStageIntLLRInputS3xD(291)(5) <= CNStageIntLLROutputS3xD(377)(4);
  VNStageIntLLRInputS3xD(328)(4) <= CNStageIntLLROutputS3xD(377)(5);
  VNStageIntLLRInputS3xD(42)(6) <= CNStageIntLLROutputS3xD(378)(0);
  VNStageIntLLRInputS3xD(92)(6) <= CNStageIntLLROutputS3xD(378)(1);
  VNStageIntLLRInputS3xD(150)(5) <= CNStageIntLLROutputS3xD(378)(2);
  VNStageIntLLRInputS3xD(226)(2) <= CNStageIntLLROutputS3xD(378)(3);
  VNStageIntLLRInputS3xD(263)(6) <= CNStageIntLLROutputS3xD(378)(4);
  VNStageIntLLRInputS3xD(383)(6) <= CNStageIntLLROutputS3xD(378)(5);
  VNStageIntLLRInputS3xD(41)(6) <= CNStageIntLLROutputS3xD(379)(0);
  VNStageIntLLRInputS3xD(85)(5) <= CNStageIntLLROutputS3xD(379)(1);
  VNStageIntLLRInputS3xD(161)(6) <= CNStageIntLLROutputS3xD(379)(2);
  VNStageIntLLRInputS3xD(198)(6) <= CNStageIntLLROutputS3xD(379)(3);
  VNStageIntLLRInputS3xD(318)(3) <= CNStageIntLLROutputS3xD(379)(4);
  VNStageIntLLRInputS3xD(337)(6) <= CNStageIntLLROutputS3xD(379)(5);
  VNStageIntLLRInputS3xD(40)(4) <= CNStageIntLLROutputS3xD(380)(0);
  VNStageIntLLRInputS3xD(96)(5) <= CNStageIntLLROutputS3xD(380)(1);
  VNStageIntLLRInputS3xD(133)(4) <= CNStageIntLLROutputS3xD(380)(2);
  VNStageIntLLRInputS3xD(253)(5) <= CNStageIntLLROutputS3xD(380)(3);
  VNStageIntLLRInputS3xD(272)(6) <= CNStageIntLLROutputS3xD(380)(4);
  VNStageIntLLRInputS3xD(334)(4) <= CNStageIntLLROutputS3xD(380)(5);
  VNStageIntLLRInputS3xD(39)(6) <= CNStageIntLLROutputS3xD(381)(0);
  VNStageIntLLRInputS3xD(68)(5) <= CNStageIntLLROutputS3xD(381)(1);
  VNStageIntLLRInputS3xD(188)(4) <= CNStageIntLLROutputS3xD(381)(2);
  VNStageIntLLRInputS3xD(207)(5) <= CNStageIntLLROutputS3xD(381)(3);
  VNStageIntLLRInputS3xD(269)(5) <= CNStageIntLLROutputS3xD(381)(4);
  VNStageIntLLRInputS3xD(368)(2) <= CNStageIntLLROutputS3xD(381)(5);
  VNStageIntLLRInputS3xD(38)(6) <= CNStageIntLLROutputS3xD(382)(0);
  VNStageIntLLRInputS3xD(123)(4) <= CNStageIntLLROutputS3xD(382)(1);
  VNStageIntLLRInputS3xD(142)(4) <= CNStageIntLLROutputS3xD(382)(2);
  VNStageIntLLRInputS3xD(204)(6) <= CNStageIntLLROutputS3xD(382)(3);
  VNStageIntLLRInputS3xD(303)(6) <= CNStageIntLLROutputS3xD(382)(4);
  VNStageIntLLRInputS3xD(325)(6) <= CNStageIntLLROutputS3xD(382)(5);
  VNStageIntLLRInputS3xD(37)(6) <= CNStageIntLLROutputS3xD(383)(0);
  VNStageIntLLRInputS3xD(77)(4) <= CNStageIntLLROutputS3xD(383)(1);
  VNStageIntLLRInputS3xD(139)(6) <= CNStageIntLLROutputS3xD(383)(2);
  VNStageIntLLRInputS3xD(238)(6) <= CNStageIntLLROutputS3xD(383)(3);
  VNStageIntLLRInputS3xD(260)(5) <= CNStageIntLLROutputS3xD(383)(4);
  VNStageIntLLRInputS3xD(374)(6) <= CNStageIntLLROutputS3xD(383)(5);

  -- Check Nodes (Iteration 4)
  CNStageIntLLRInputS4xD(53)(0) <= VNStageIntLLROutputS3xD(0)(0);
  CNStageIntLLRInputS4xD(110)(0) <= VNStageIntLLROutputS3xD(0)(1);
  CNStageIntLLRInputS4xD(170)(0) <= VNStageIntLLROutputS3xD(0)(2);
  CNStageIntLLRInputS4xD(224)(0) <= VNStageIntLLROutputS3xD(0)(3);
  CNStageIntLLRInputS4xD(279)(0) <= VNStageIntLLROutputS3xD(0)(4);
  CNStageIntLLRInputS4xD(332)(0) <= VNStageIntLLROutputS3xD(0)(5);
  CNStageIntLLRInputS4xD(51)(0) <= VNStageIntLLROutputS3xD(1)(0);
  CNStageIntLLRInputS4xD(139)(0) <= VNStageIntLLROutputS3xD(1)(1);
  CNStageIntLLRInputS4xD(223)(0) <= VNStageIntLLROutputS3xD(1)(2);
  CNStageIntLLRInputS4xD(241)(0) <= VNStageIntLLROutputS3xD(1)(3);
  CNStageIntLLRInputS4xD(307)(0) <= VNStageIntLLROutputS3xD(1)(4);
  CNStageIntLLRInputS4xD(356)(0) <= VNStageIntLLROutputS3xD(1)(5);
  CNStageIntLLRInputS4xD(50)(0) <= VNStageIntLLROutputS3xD(2)(0);
  CNStageIntLLRInputS4xD(92)(0) <= VNStageIntLLROutputS3xD(2)(1);
  CNStageIntLLRInputS4xD(138)(0) <= VNStageIntLLROutputS3xD(2)(2);
  CNStageIntLLRInputS4xD(222)(0) <= VNStageIntLLROutputS3xD(2)(3);
  CNStageIntLLRInputS4xD(240)(0) <= VNStageIntLLROutputS3xD(2)(4);
  CNStageIntLLRInputS4xD(306)(0) <= VNStageIntLLROutputS3xD(2)(5);
  CNStageIntLLRInputS4xD(355)(0) <= VNStageIntLLROutputS3xD(2)(6);
  CNStageIntLLRInputS4xD(91)(0) <= VNStageIntLLROutputS3xD(3)(0);
  CNStageIntLLRInputS4xD(137)(0) <= VNStageIntLLROutputS3xD(3)(1);
  CNStageIntLLRInputS4xD(221)(0) <= VNStageIntLLROutputS3xD(3)(2);
  CNStageIntLLRInputS4xD(239)(0) <= VNStageIntLLROutputS3xD(3)(3);
  CNStageIntLLRInputS4xD(305)(0) <= VNStageIntLLROutputS3xD(3)(4);
  CNStageIntLLRInputS4xD(49)(0) <= VNStageIntLLROutputS3xD(4)(0);
  CNStageIntLLRInputS4xD(90)(0) <= VNStageIntLLROutputS3xD(4)(1);
  CNStageIntLLRInputS4xD(220)(0) <= VNStageIntLLROutputS3xD(4)(2);
  CNStageIntLLRInputS4xD(238)(0) <= VNStageIntLLROutputS3xD(4)(3);
  CNStageIntLLRInputS4xD(304)(0) <= VNStageIntLLROutputS3xD(4)(4);
  CNStageIntLLRInputS4xD(354)(0) <= VNStageIntLLROutputS3xD(4)(5);
  CNStageIntLLRInputS4xD(48)(0) <= VNStageIntLLROutputS3xD(5)(0);
  CNStageIntLLRInputS4xD(89)(0) <= VNStageIntLLROutputS3xD(5)(1);
  CNStageIntLLRInputS4xD(136)(0) <= VNStageIntLLROutputS3xD(5)(2);
  CNStageIntLLRInputS4xD(219)(0) <= VNStageIntLLROutputS3xD(5)(3);
  CNStageIntLLRInputS4xD(237)(0) <= VNStageIntLLROutputS3xD(5)(4);
  CNStageIntLLRInputS4xD(303)(0) <= VNStageIntLLROutputS3xD(5)(5);
  CNStageIntLLRInputS4xD(353)(0) <= VNStageIntLLROutputS3xD(5)(6);
  CNStageIntLLRInputS4xD(47)(0) <= VNStageIntLLROutputS3xD(6)(0);
  CNStageIntLLRInputS4xD(88)(0) <= VNStageIntLLROutputS3xD(6)(1);
  CNStageIntLLRInputS4xD(135)(0) <= VNStageIntLLROutputS3xD(6)(2);
  CNStageIntLLRInputS4xD(218)(0) <= VNStageIntLLROutputS3xD(6)(3);
  CNStageIntLLRInputS4xD(236)(0) <= VNStageIntLLROutputS3xD(6)(4);
  CNStageIntLLRInputS4xD(302)(0) <= VNStageIntLLROutputS3xD(6)(5);
  CNStageIntLLRInputS4xD(352)(0) <= VNStageIntLLROutputS3xD(6)(6);
  CNStageIntLLRInputS4xD(46)(0) <= VNStageIntLLROutputS3xD(7)(0);
  CNStageIntLLRInputS4xD(87)(0) <= VNStageIntLLROutputS3xD(7)(1);
  CNStageIntLLRInputS4xD(134)(0) <= VNStageIntLLROutputS3xD(7)(2);
  CNStageIntLLRInputS4xD(217)(0) <= VNStageIntLLROutputS3xD(7)(3);
  CNStageIntLLRInputS4xD(235)(0) <= VNStageIntLLROutputS3xD(7)(4);
  CNStageIntLLRInputS4xD(301)(0) <= VNStageIntLLROutputS3xD(7)(5);
  CNStageIntLLRInputS4xD(351)(0) <= VNStageIntLLROutputS3xD(7)(6);
  CNStageIntLLRInputS4xD(45)(0) <= VNStageIntLLROutputS3xD(8)(0);
  CNStageIntLLRInputS4xD(133)(0) <= VNStageIntLLROutputS3xD(8)(1);
  CNStageIntLLRInputS4xD(216)(0) <= VNStageIntLLROutputS3xD(8)(2);
  CNStageIntLLRInputS4xD(44)(0) <= VNStageIntLLROutputS3xD(9)(0);
  CNStageIntLLRInputS4xD(86)(0) <= VNStageIntLLROutputS3xD(9)(1);
  CNStageIntLLRInputS4xD(132)(0) <= VNStageIntLLROutputS3xD(9)(2);
  CNStageIntLLRInputS4xD(215)(0) <= VNStageIntLLROutputS3xD(9)(3);
  CNStageIntLLRInputS4xD(234)(0) <= VNStageIntLLROutputS3xD(9)(4);
  CNStageIntLLRInputS4xD(300)(0) <= VNStageIntLLROutputS3xD(9)(5);
  CNStageIntLLRInputS4xD(350)(0) <= VNStageIntLLROutputS3xD(9)(6);
  CNStageIntLLRInputS4xD(43)(0) <= VNStageIntLLROutputS3xD(10)(0);
  CNStageIntLLRInputS4xD(85)(0) <= VNStageIntLLROutputS3xD(10)(1);
  CNStageIntLLRInputS4xD(131)(0) <= VNStageIntLLROutputS3xD(10)(2);
  CNStageIntLLRInputS4xD(233)(0) <= VNStageIntLLROutputS3xD(10)(3);
  CNStageIntLLRInputS4xD(349)(0) <= VNStageIntLLROutputS3xD(10)(4);
  CNStageIntLLRInputS4xD(42)(0) <= VNStageIntLLROutputS3xD(11)(0);
  CNStageIntLLRInputS4xD(84)(0) <= VNStageIntLLROutputS3xD(11)(1);
  CNStageIntLLRInputS4xD(130)(0) <= VNStageIntLLROutputS3xD(11)(2);
  CNStageIntLLRInputS4xD(214)(0) <= VNStageIntLLROutputS3xD(11)(3);
  CNStageIntLLRInputS4xD(232)(0) <= VNStageIntLLROutputS3xD(11)(4);
  CNStageIntLLRInputS4xD(348)(0) <= VNStageIntLLROutputS3xD(11)(5);
  CNStageIntLLRInputS4xD(41)(0) <= VNStageIntLLROutputS3xD(12)(0);
  CNStageIntLLRInputS4xD(83)(0) <= VNStageIntLLROutputS3xD(12)(1);
  CNStageIntLLRInputS4xD(129)(0) <= VNStageIntLLROutputS3xD(12)(2);
  CNStageIntLLRInputS4xD(213)(0) <= VNStageIntLLROutputS3xD(12)(3);
  CNStageIntLLRInputS4xD(231)(0) <= VNStageIntLLROutputS3xD(12)(4);
  CNStageIntLLRInputS4xD(299)(0) <= VNStageIntLLROutputS3xD(12)(5);
  CNStageIntLLRInputS4xD(347)(0) <= VNStageIntLLROutputS3xD(12)(6);
  CNStageIntLLRInputS4xD(82)(0) <= VNStageIntLLROutputS3xD(13)(0);
  CNStageIntLLRInputS4xD(128)(0) <= VNStageIntLLROutputS3xD(13)(1);
  CNStageIntLLRInputS4xD(212)(0) <= VNStageIntLLROutputS3xD(13)(2);
  CNStageIntLLRInputS4xD(230)(0) <= VNStageIntLLROutputS3xD(13)(3);
  CNStageIntLLRInputS4xD(298)(0) <= VNStageIntLLROutputS3xD(13)(4);
  CNStageIntLLRInputS4xD(346)(0) <= VNStageIntLLROutputS3xD(13)(5);
  CNStageIntLLRInputS4xD(40)(0) <= VNStageIntLLROutputS3xD(14)(0);
  CNStageIntLLRInputS4xD(81)(0) <= VNStageIntLLROutputS3xD(14)(1);
  CNStageIntLLRInputS4xD(127)(0) <= VNStageIntLLROutputS3xD(14)(2);
  CNStageIntLLRInputS4xD(211)(0) <= VNStageIntLLROutputS3xD(14)(3);
  CNStageIntLLRInputS4xD(229)(0) <= VNStageIntLLROutputS3xD(14)(4);
  CNStageIntLLRInputS4xD(297)(0) <= VNStageIntLLROutputS3xD(14)(5);
  CNStageIntLLRInputS4xD(345)(0) <= VNStageIntLLROutputS3xD(14)(6);
  CNStageIntLLRInputS4xD(39)(0) <= VNStageIntLLROutputS3xD(15)(0);
  CNStageIntLLRInputS4xD(80)(0) <= VNStageIntLLROutputS3xD(15)(1);
  CNStageIntLLRInputS4xD(126)(0) <= VNStageIntLLROutputS3xD(15)(2);
  CNStageIntLLRInputS4xD(210)(0) <= VNStageIntLLROutputS3xD(15)(3);
  CNStageIntLLRInputS4xD(228)(0) <= VNStageIntLLROutputS3xD(15)(4);
  CNStageIntLLRInputS4xD(296)(0) <= VNStageIntLLROutputS3xD(15)(5);
  CNStageIntLLRInputS4xD(344)(0) <= VNStageIntLLROutputS3xD(15)(6);
  CNStageIntLLRInputS4xD(38)(0) <= VNStageIntLLROutputS3xD(16)(0);
  CNStageIntLLRInputS4xD(125)(0) <= VNStageIntLLROutputS3xD(16)(1);
  CNStageIntLLRInputS4xD(209)(0) <= VNStageIntLLROutputS3xD(16)(2);
  CNStageIntLLRInputS4xD(227)(0) <= VNStageIntLLROutputS3xD(16)(3);
  CNStageIntLLRInputS4xD(295)(0) <= VNStageIntLLROutputS3xD(16)(4);
  CNStageIntLLRInputS4xD(343)(0) <= VNStageIntLLROutputS3xD(16)(5);
  CNStageIntLLRInputS4xD(37)(0) <= VNStageIntLLROutputS3xD(17)(0);
  CNStageIntLLRInputS4xD(79)(0) <= VNStageIntLLROutputS3xD(17)(1);
  CNStageIntLLRInputS4xD(124)(0) <= VNStageIntLLROutputS3xD(17)(2);
  CNStageIntLLRInputS4xD(208)(0) <= VNStageIntLLROutputS3xD(17)(3);
  CNStageIntLLRInputS4xD(226)(0) <= VNStageIntLLROutputS3xD(17)(4);
  CNStageIntLLRInputS4xD(294)(0) <= VNStageIntLLROutputS3xD(17)(5);
  CNStageIntLLRInputS4xD(342)(0) <= VNStageIntLLROutputS3xD(17)(6);
  CNStageIntLLRInputS4xD(36)(0) <= VNStageIntLLROutputS3xD(18)(0);
  CNStageIntLLRInputS4xD(78)(0) <= VNStageIntLLROutputS3xD(18)(1);
  CNStageIntLLRInputS4xD(123)(0) <= VNStageIntLLROutputS3xD(18)(2);
  CNStageIntLLRInputS4xD(207)(0) <= VNStageIntLLROutputS3xD(18)(3);
  CNStageIntLLRInputS4xD(225)(0) <= VNStageIntLLROutputS3xD(18)(4);
  CNStageIntLLRInputS4xD(293)(0) <= VNStageIntLLROutputS3xD(18)(5);
  CNStageIntLLRInputS4xD(341)(0) <= VNStageIntLLROutputS3xD(18)(6);
  CNStageIntLLRInputS4xD(35)(0) <= VNStageIntLLROutputS3xD(19)(0);
  CNStageIntLLRInputS4xD(77)(0) <= VNStageIntLLROutputS3xD(19)(1);
  CNStageIntLLRInputS4xD(122)(0) <= VNStageIntLLROutputS3xD(19)(2);
  CNStageIntLLRInputS4xD(278)(0) <= VNStageIntLLROutputS3xD(19)(3);
  CNStageIntLLRInputS4xD(340)(0) <= VNStageIntLLROutputS3xD(19)(4);
  CNStageIntLLRInputS4xD(34)(0) <= VNStageIntLLROutputS3xD(20)(0);
  CNStageIntLLRInputS4xD(76)(0) <= VNStageIntLLROutputS3xD(20)(1);
  CNStageIntLLRInputS4xD(277)(0) <= VNStageIntLLROutputS3xD(20)(2);
  CNStageIntLLRInputS4xD(292)(0) <= VNStageIntLLROutputS3xD(20)(3);
  CNStageIntLLRInputS4xD(339)(0) <= VNStageIntLLROutputS3xD(20)(4);
  CNStageIntLLRInputS4xD(33)(0) <= VNStageIntLLROutputS3xD(21)(0);
  CNStageIntLLRInputS4xD(75)(0) <= VNStageIntLLROutputS3xD(21)(1);
  CNStageIntLLRInputS4xD(121)(0) <= VNStageIntLLROutputS3xD(21)(2);
  CNStageIntLLRInputS4xD(206)(0) <= VNStageIntLLROutputS3xD(21)(3);
  CNStageIntLLRInputS4xD(276)(0) <= VNStageIntLLROutputS3xD(21)(4);
  CNStageIntLLRInputS4xD(291)(0) <= VNStageIntLLROutputS3xD(21)(5);
  CNStageIntLLRInputS4xD(338)(0) <= VNStageIntLLROutputS3xD(21)(6);
  CNStageIntLLRInputS4xD(32)(0) <= VNStageIntLLROutputS3xD(22)(0);
  CNStageIntLLRInputS4xD(74)(0) <= VNStageIntLLROutputS3xD(22)(1);
  CNStageIntLLRInputS4xD(120)(0) <= VNStageIntLLROutputS3xD(22)(2);
  CNStageIntLLRInputS4xD(205)(0) <= VNStageIntLLROutputS3xD(22)(3);
  CNStageIntLLRInputS4xD(275)(0) <= VNStageIntLLROutputS3xD(22)(4);
  CNStageIntLLRInputS4xD(290)(0) <= VNStageIntLLROutputS3xD(22)(5);
  CNStageIntLLRInputS4xD(337)(0) <= VNStageIntLLROutputS3xD(22)(6);
  CNStageIntLLRInputS4xD(31)(0) <= VNStageIntLLROutputS3xD(23)(0);
  CNStageIntLLRInputS4xD(73)(0) <= VNStageIntLLROutputS3xD(23)(1);
  CNStageIntLLRInputS4xD(119)(0) <= VNStageIntLLROutputS3xD(23)(2);
  CNStageIntLLRInputS4xD(204)(0) <= VNStageIntLLROutputS3xD(23)(3);
  CNStageIntLLRInputS4xD(274)(0) <= VNStageIntLLROutputS3xD(23)(4);
  CNStageIntLLRInputS4xD(289)(0) <= VNStageIntLLROutputS3xD(23)(5);
  CNStageIntLLRInputS4xD(336)(0) <= VNStageIntLLROutputS3xD(23)(6);
  CNStageIntLLRInputS4xD(30)(0) <= VNStageIntLLROutputS3xD(24)(0);
  CNStageIntLLRInputS4xD(72)(0) <= VNStageIntLLROutputS3xD(24)(1);
  CNStageIntLLRInputS4xD(118)(0) <= VNStageIntLLROutputS3xD(24)(2);
  CNStageIntLLRInputS4xD(203)(0) <= VNStageIntLLROutputS3xD(24)(3);
  CNStageIntLLRInputS4xD(273)(0) <= VNStageIntLLROutputS3xD(24)(4);
  CNStageIntLLRInputS4xD(288)(0) <= VNStageIntLLROutputS3xD(24)(5);
  CNStageIntLLRInputS4xD(335)(0) <= VNStageIntLLROutputS3xD(24)(6);
  CNStageIntLLRInputS4xD(29)(0) <= VNStageIntLLROutputS3xD(25)(0);
  CNStageIntLLRInputS4xD(71)(0) <= VNStageIntLLROutputS3xD(25)(1);
  CNStageIntLLRInputS4xD(117)(0) <= VNStageIntLLROutputS3xD(25)(2);
  CNStageIntLLRInputS4xD(202)(0) <= VNStageIntLLROutputS3xD(25)(3);
  CNStageIntLLRInputS4xD(287)(0) <= VNStageIntLLROutputS3xD(25)(4);
  CNStageIntLLRInputS4xD(28)(0) <= VNStageIntLLROutputS3xD(26)(0);
  CNStageIntLLRInputS4xD(70)(0) <= VNStageIntLLROutputS3xD(26)(1);
  CNStageIntLLRInputS4xD(116)(0) <= VNStageIntLLROutputS3xD(26)(2);
  CNStageIntLLRInputS4xD(201)(0) <= VNStageIntLLROutputS3xD(26)(3);
  CNStageIntLLRInputS4xD(272)(0) <= VNStageIntLLROutputS3xD(26)(4);
  CNStageIntLLRInputS4xD(286)(0) <= VNStageIntLLROutputS3xD(26)(5);
  CNStageIntLLRInputS4xD(334)(0) <= VNStageIntLLROutputS3xD(26)(6);
  CNStageIntLLRInputS4xD(27)(0) <= VNStageIntLLROutputS3xD(27)(0);
  CNStageIntLLRInputS4xD(69)(0) <= VNStageIntLLROutputS3xD(27)(1);
  CNStageIntLLRInputS4xD(115)(0) <= VNStageIntLLROutputS3xD(27)(2);
  CNStageIntLLRInputS4xD(200)(0) <= VNStageIntLLROutputS3xD(27)(3);
  CNStageIntLLRInputS4xD(285)(0) <= VNStageIntLLROutputS3xD(27)(4);
  CNStageIntLLRInputS4xD(26)(0) <= VNStageIntLLROutputS3xD(28)(0);
  CNStageIntLLRInputS4xD(68)(0) <= VNStageIntLLROutputS3xD(28)(1);
  CNStageIntLLRInputS4xD(114)(0) <= VNStageIntLLROutputS3xD(28)(2);
  CNStageIntLLRInputS4xD(199)(0) <= VNStageIntLLROutputS3xD(28)(3);
  CNStageIntLLRInputS4xD(271)(0) <= VNStageIntLLROutputS3xD(28)(4);
  CNStageIntLLRInputS4xD(333)(0) <= VNStageIntLLROutputS3xD(28)(5);
  CNStageIntLLRInputS4xD(25)(0) <= VNStageIntLLROutputS3xD(29)(0);
  CNStageIntLLRInputS4xD(67)(0) <= VNStageIntLLROutputS3xD(29)(1);
  CNStageIntLLRInputS4xD(113)(0) <= VNStageIntLLROutputS3xD(29)(2);
  CNStageIntLLRInputS4xD(270)(0) <= VNStageIntLLROutputS3xD(29)(3);
  CNStageIntLLRInputS4xD(24)(0) <= VNStageIntLLROutputS3xD(30)(0);
  CNStageIntLLRInputS4xD(66)(0) <= VNStageIntLLROutputS3xD(30)(1);
  CNStageIntLLRInputS4xD(112)(0) <= VNStageIntLLROutputS3xD(30)(2);
  CNStageIntLLRInputS4xD(198)(0) <= VNStageIntLLROutputS3xD(30)(3);
  CNStageIntLLRInputS4xD(269)(0) <= VNStageIntLLROutputS3xD(30)(4);
  CNStageIntLLRInputS4xD(284)(0) <= VNStageIntLLROutputS3xD(30)(5);
  CNStageIntLLRInputS4xD(23)(0) <= VNStageIntLLROutputS3xD(31)(0);
  CNStageIntLLRInputS4xD(65)(0) <= VNStageIntLLROutputS3xD(31)(1);
  CNStageIntLLRInputS4xD(197)(0) <= VNStageIntLLROutputS3xD(31)(2);
  CNStageIntLLRInputS4xD(283)(0) <= VNStageIntLLROutputS3xD(31)(3);
  CNStageIntLLRInputS4xD(22)(0) <= VNStageIntLLROutputS3xD(32)(0);
  CNStageIntLLRInputS4xD(64)(0) <= VNStageIntLLROutputS3xD(32)(1);
  CNStageIntLLRInputS4xD(111)(0) <= VNStageIntLLROutputS3xD(32)(2);
  CNStageIntLLRInputS4xD(268)(0) <= VNStageIntLLROutputS3xD(32)(3);
  CNStageIntLLRInputS4xD(21)(0) <= VNStageIntLLROutputS3xD(33)(0);
  CNStageIntLLRInputS4xD(63)(0) <= VNStageIntLLROutputS3xD(33)(1);
  CNStageIntLLRInputS4xD(169)(0) <= VNStageIntLLROutputS3xD(33)(2);
  CNStageIntLLRInputS4xD(196)(0) <= VNStageIntLLROutputS3xD(33)(3);
  CNStageIntLLRInputS4xD(267)(0) <= VNStageIntLLROutputS3xD(33)(4);
  CNStageIntLLRInputS4xD(282)(0) <= VNStageIntLLROutputS3xD(33)(5);
  CNStageIntLLRInputS4xD(20)(0) <= VNStageIntLLROutputS3xD(34)(0);
  CNStageIntLLRInputS4xD(62)(0) <= VNStageIntLLROutputS3xD(34)(1);
  CNStageIntLLRInputS4xD(168)(0) <= VNStageIntLLROutputS3xD(34)(2);
  CNStageIntLLRInputS4xD(195)(0) <= VNStageIntLLROutputS3xD(34)(3);
  CNStageIntLLRInputS4xD(266)(0) <= VNStageIntLLROutputS3xD(34)(4);
  CNStageIntLLRInputS4xD(281)(0) <= VNStageIntLLROutputS3xD(34)(5);
  CNStageIntLLRInputS4xD(19)(0) <= VNStageIntLLROutputS3xD(35)(0);
  CNStageIntLLRInputS4xD(61)(0) <= VNStageIntLLROutputS3xD(35)(1);
  CNStageIntLLRInputS4xD(167)(0) <= VNStageIntLLROutputS3xD(35)(2);
  CNStageIntLLRInputS4xD(194)(0) <= VNStageIntLLROutputS3xD(35)(3);
  CNStageIntLLRInputS4xD(265)(0) <= VNStageIntLLROutputS3xD(35)(4);
  CNStageIntLLRInputS4xD(280)(0) <= VNStageIntLLROutputS3xD(35)(5);
  CNStageIntLLRInputS4xD(18)(0) <= VNStageIntLLROutputS3xD(36)(0);
  CNStageIntLLRInputS4xD(60)(0) <= VNStageIntLLROutputS3xD(36)(1);
  CNStageIntLLRInputS4xD(166)(0) <= VNStageIntLLROutputS3xD(36)(2);
  CNStageIntLLRInputS4xD(264)(0) <= VNStageIntLLROutputS3xD(36)(3);
  CNStageIntLLRInputS4xD(17)(0) <= VNStageIntLLROutputS3xD(37)(0);
  CNStageIntLLRInputS4xD(59)(0) <= VNStageIntLLROutputS3xD(37)(1);
  CNStageIntLLRInputS4xD(165)(0) <= VNStageIntLLROutputS3xD(37)(2);
  CNStageIntLLRInputS4xD(193)(0) <= VNStageIntLLROutputS3xD(37)(3);
  CNStageIntLLRInputS4xD(263)(0) <= VNStageIntLLROutputS3xD(37)(4);
  CNStageIntLLRInputS4xD(331)(0) <= VNStageIntLLROutputS3xD(37)(5);
  CNStageIntLLRInputS4xD(383)(0) <= VNStageIntLLROutputS3xD(37)(6);
  CNStageIntLLRInputS4xD(16)(0) <= VNStageIntLLROutputS3xD(38)(0);
  CNStageIntLLRInputS4xD(58)(0) <= VNStageIntLLROutputS3xD(38)(1);
  CNStageIntLLRInputS4xD(164)(0) <= VNStageIntLLROutputS3xD(38)(2);
  CNStageIntLLRInputS4xD(192)(0) <= VNStageIntLLROutputS3xD(38)(3);
  CNStageIntLLRInputS4xD(262)(0) <= VNStageIntLLROutputS3xD(38)(4);
  CNStageIntLLRInputS4xD(330)(0) <= VNStageIntLLROutputS3xD(38)(5);
  CNStageIntLLRInputS4xD(382)(0) <= VNStageIntLLROutputS3xD(38)(6);
  CNStageIntLLRInputS4xD(15)(0) <= VNStageIntLLROutputS3xD(39)(0);
  CNStageIntLLRInputS4xD(57)(0) <= VNStageIntLLROutputS3xD(39)(1);
  CNStageIntLLRInputS4xD(163)(0) <= VNStageIntLLROutputS3xD(39)(2);
  CNStageIntLLRInputS4xD(191)(0) <= VNStageIntLLROutputS3xD(39)(3);
  CNStageIntLLRInputS4xD(261)(0) <= VNStageIntLLROutputS3xD(39)(4);
  CNStageIntLLRInputS4xD(329)(0) <= VNStageIntLLROutputS3xD(39)(5);
  CNStageIntLLRInputS4xD(381)(0) <= VNStageIntLLROutputS3xD(39)(6);
  CNStageIntLLRInputS4xD(14)(0) <= VNStageIntLLROutputS3xD(40)(0);
  CNStageIntLLRInputS4xD(56)(0) <= VNStageIntLLROutputS3xD(40)(1);
  CNStageIntLLRInputS4xD(162)(0) <= VNStageIntLLROutputS3xD(40)(2);
  CNStageIntLLRInputS4xD(260)(0) <= VNStageIntLLROutputS3xD(40)(3);
  CNStageIntLLRInputS4xD(380)(0) <= VNStageIntLLROutputS3xD(40)(4);
  CNStageIntLLRInputS4xD(13)(0) <= VNStageIntLLROutputS3xD(41)(0);
  CNStageIntLLRInputS4xD(55)(0) <= VNStageIntLLROutputS3xD(41)(1);
  CNStageIntLLRInputS4xD(161)(0) <= VNStageIntLLROutputS3xD(41)(2);
  CNStageIntLLRInputS4xD(190)(0) <= VNStageIntLLROutputS3xD(41)(3);
  CNStageIntLLRInputS4xD(259)(0) <= VNStageIntLLROutputS3xD(41)(4);
  CNStageIntLLRInputS4xD(328)(0) <= VNStageIntLLROutputS3xD(41)(5);
  CNStageIntLLRInputS4xD(379)(0) <= VNStageIntLLROutputS3xD(41)(6);
  CNStageIntLLRInputS4xD(12)(0) <= VNStageIntLLROutputS3xD(42)(0);
  CNStageIntLLRInputS4xD(54)(0) <= VNStageIntLLROutputS3xD(42)(1);
  CNStageIntLLRInputS4xD(160)(0) <= VNStageIntLLROutputS3xD(42)(2);
  CNStageIntLLRInputS4xD(189)(0) <= VNStageIntLLROutputS3xD(42)(3);
  CNStageIntLLRInputS4xD(258)(0) <= VNStageIntLLROutputS3xD(42)(4);
  CNStageIntLLRInputS4xD(327)(0) <= VNStageIntLLROutputS3xD(42)(5);
  CNStageIntLLRInputS4xD(378)(0) <= VNStageIntLLROutputS3xD(42)(6);
  CNStageIntLLRInputS4xD(109)(0) <= VNStageIntLLROutputS3xD(43)(0);
  CNStageIntLLRInputS4xD(159)(0) <= VNStageIntLLROutputS3xD(43)(1);
  CNStageIntLLRInputS4xD(188)(0) <= VNStageIntLLROutputS3xD(43)(2);
  CNStageIntLLRInputS4xD(257)(0) <= VNStageIntLLROutputS3xD(43)(3);
  CNStageIntLLRInputS4xD(326)(0) <= VNStageIntLLROutputS3xD(43)(4);
  CNStageIntLLRInputS4xD(377)(0) <= VNStageIntLLROutputS3xD(43)(5);
  CNStageIntLLRInputS4xD(11)(0) <= VNStageIntLLROutputS3xD(44)(0);
  CNStageIntLLRInputS4xD(108)(0) <= VNStageIntLLROutputS3xD(44)(1);
  CNStageIntLLRInputS4xD(158)(0) <= VNStageIntLLROutputS3xD(44)(2);
  CNStageIntLLRInputS4xD(187)(0) <= VNStageIntLLROutputS3xD(44)(3);
  CNStageIntLLRInputS4xD(256)(0) <= VNStageIntLLROutputS3xD(44)(4);
  CNStageIntLLRInputS4xD(325)(0) <= VNStageIntLLROutputS3xD(44)(5);
  CNStageIntLLRInputS4xD(376)(0) <= VNStageIntLLROutputS3xD(44)(6);
  CNStageIntLLRInputS4xD(10)(0) <= VNStageIntLLROutputS3xD(45)(0);
  CNStageIntLLRInputS4xD(107)(0) <= VNStageIntLLROutputS3xD(45)(1);
  CNStageIntLLRInputS4xD(157)(0) <= VNStageIntLLROutputS3xD(45)(2);
  CNStageIntLLRInputS4xD(186)(0) <= VNStageIntLLROutputS3xD(45)(3);
  CNStageIntLLRInputS4xD(255)(0) <= VNStageIntLLROutputS3xD(45)(4);
  CNStageIntLLRInputS4xD(324)(0) <= VNStageIntLLROutputS3xD(45)(5);
  CNStageIntLLRInputS4xD(375)(0) <= VNStageIntLLROutputS3xD(45)(6);
  CNStageIntLLRInputS4xD(9)(0) <= VNStageIntLLROutputS3xD(46)(0);
  CNStageIntLLRInputS4xD(106)(0) <= VNStageIntLLROutputS3xD(46)(1);
  CNStageIntLLRInputS4xD(156)(0) <= VNStageIntLLROutputS3xD(46)(2);
  CNStageIntLLRInputS4xD(185)(0) <= VNStageIntLLROutputS3xD(46)(3);
  CNStageIntLLRInputS4xD(254)(0) <= VNStageIntLLROutputS3xD(46)(4);
  CNStageIntLLRInputS4xD(323)(0) <= VNStageIntLLROutputS3xD(46)(5);
  CNStageIntLLRInputS4xD(374)(0) <= VNStageIntLLROutputS3xD(46)(6);
  CNStageIntLLRInputS4xD(8)(0) <= VNStageIntLLROutputS3xD(47)(0);
  CNStageIntLLRInputS4xD(155)(0) <= VNStageIntLLROutputS3xD(47)(1);
  CNStageIntLLRInputS4xD(253)(0) <= VNStageIntLLROutputS3xD(47)(2);
  CNStageIntLLRInputS4xD(373)(0) <= VNStageIntLLROutputS3xD(47)(3);
  CNStageIntLLRInputS4xD(7)(0) <= VNStageIntLLROutputS3xD(48)(0);
  CNStageIntLLRInputS4xD(154)(0) <= VNStageIntLLROutputS3xD(48)(1);
  CNStageIntLLRInputS4xD(322)(0) <= VNStageIntLLROutputS3xD(48)(2);
  CNStageIntLLRInputS4xD(372)(0) <= VNStageIntLLROutputS3xD(48)(3);
  CNStageIntLLRInputS4xD(6)(0) <= VNStageIntLLROutputS3xD(49)(0);
  CNStageIntLLRInputS4xD(105)(0) <= VNStageIntLLROutputS3xD(49)(1);
  CNStageIntLLRInputS4xD(153)(0) <= VNStageIntLLROutputS3xD(49)(2);
  CNStageIntLLRInputS4xD(184)(0) <= VNStageIntLLROutputS3xD(49)(3);
  CNStageIntLLRInputS4xD(252)(0) <= VNStageIntLLROutputS3xD(49)(4);
  CNStageIntLLRInputS4xD(321)(0) <= VNStageIntLLROutputS3xD(49)(5);
  CNStageIntLLRInputS4xD(371)(0) <= VNStageIntLLROutputS3xD(49)(6);
  CNStageIntLLRInputS4xD(5)(0) <= VNStageIntLLROutputS3xD(50)(0);
  CNStageIntLLRInputS4xD(104)(0) <= VNStageIntLLROutputS3xD(50)(1);
  CNStageIntLLRInputS4xD(152)(0) <= VNStageIntLLROutputS3xD(50)(2);
  CNStageIntLLRInputS4xD(183)(0) <= VNStageIntLLROutputS3xD(50)(3);
  CNStageIntLLRInputS4xD(251)(0) <= VNStageIntLLROutputS3xD(50)(4);
  CNStageIntLLRInputS4xD(320)(0) <= VNStageIntLLROutputS3xD(50)(5);
  CNStageIntLLRInputS4xD(370)(0) <= VNStageIntLLROutputS3xD(50)(6);
  CNStageIntLLRInputS4xD(4)(0) <= VNStageIntLLROutputS3xD(51)(0);
  CNStageIntLLRInputS4xD(103)(0) <= VNStageIntLLROutputS3xD(51)(1);
  CNStageIntLLRInputS4xD(182)(0) <= VNStageIntLLROutputS3xD(51)(2);
  CNStageIntLLRInputS4xD(250)(0) <= VNStageIntLLROutputS3xD(51)(3);
  CNStageIntLLRInputS4xD(319)(0) <= VNStageIntLLROutputS3xD(51)(4);
  CNStageIntLLRInputS4xD(369)(0) <= VNStageIntLLROutputS3xD(51)(5);
  CNStageIntLLRInputS4xD(102)(0) <= VNStageIntLLROutputS3xD(52)(0);
  CNStageIntLLRInputS4xD(151)(0) <= VNStageIntLLROutputS3xD(52)(1);
  CNStageIntLLRInputS4xD(181)(0) <= VNStageIntLLROutputS3xD(52)(2);
  CNStageIntLLRInputS4xD(318)(0) <= VNStageIntLLROutputS3xD(52)(3);
  CNStageIntLLRInputS4xD(368)(0) <= VNStageIntLLROutputS3xD(52)(4);
  CNStageIntLLRInputS4xD(3)(0) <= VNStageIntLLROutputS3xD(53)(0);
  CNStageIntLLRInputS4xD(150)(0) <= VNStageIntLLROutputS3xD(53)(1);
  CNStageIntLLRInputS4xD(180)(0) <= VNStageIntLLROutputS3xD(53)(2);
  CNStageIntLLRInputS4xD(249)(0) <= VNStageIntLLROutputS3xD(53)(3);
  CNStageIntLLRInputS4xD(317)(0) <= VNStageIntLLROutputS3xD(53)(4);
  CNStageIntLLRInputS4xD(367)(0) <= VNStageIntLLROutputS3xD(53)(5);
  CNStageIntLLRInputS4xD(2)(0) <= VNStageIntLLROutputS3xD(54)(0);
  CNStageIntLLRInputS4xD(101)(0) <= VNStageIntLLROutputS3xD(54)(1);
  CNStageIntLLRInputS4xD(149)(0) <= VNStageIntLLROutputS3xD(54)(2);
  CNStageIntLLRInputS4xD(179)(0) <= VNStageIntLLROutputS3xD(54)(3);
  CNStageIntLLRInputS4xD(316)(0) <= VNStageIntLLROutputS3xD(54)(4);
  CNStageIntLLRInputS4xD(366)(0) <= VNStageIntLLROutputS3xD(54)(5);
  CNStageIntLLRInputS4xD(1)(0) <= VNStageIntLLROutputS3xD(55)(0);
  CNStageIntLLRInputS4xD(100)(0) <= VNStageIntLLROutputS3xD(55)(1);
  CNStageIntLLRInputS4xD(148)(0) <= VNStageIntLLROutputS3xD(55)(2);
  CNStageIntLLRInputS4xD(178)(0) <= VNStageIntLLROutputS3xD(55)(3);
  CNStageIntLLRInputS4xD(248)(0) <= VNStageIntLLROutputS3xD(55)(4);
  CNStageIntLLRInputS4xD(315)(0) <= VNStageIntLLROutputS3xD(55)(5);
  CNStageIntLLRInputS4xD(365)(0) <= VNStageIntLLROutputS3xD(55)(6);
  CNStageIntLLRInputS4xD(0)(0) <= VNStageIntLLROutputS3xD(56)(0);
  CNStageIntLLRInputS4xD(99)(0) <= VNStageIntLLROutputS3xD(56)(1);
  CNStageIntLLRInputS4xD(147)(0) <= VNStageIntLLROutputS3xD(56)(2);
  CNStageIntLLRInputS4xD(177)(0) <= VNStageIntLLROutputS3xD(56)(3);
  CNStageIntLLRInputS4xD(247)(0) <= VNStageIntLLROutputS3xD(56)(4);
  CNStageIntLLRInputS4xD(314)(0) <= VNStageIntLLROutputS3xD(56)(5);
  CNStageIntLLRInputS4xD(364)(0) <= VNStageIntLLROutputS3xD(56)(6);
  CNStageIntLLRInputS4xD(98)(0) <= VNStageIntLLROutputS3xD(57)(0);
  CNStageIntLLRInputS4xD(146)(0) <= VNStageIntLLROutputS3xD(57)(1);
  CNStageIntLLRInputS4xD(176)(0) <= VNStageIntLLROutputS3xD(57)(2);
  CNStageIntLLRInputS4xD(246)(0) <= VNStageIntLLROutputS3xD(57)(3);
  CNStageIntLLRInputS4xD(313)(0) <= VNStageIntLLROutputS3xD(57)(4);
  CNStageIntLLRInputS4xD(363)(0) <= VNStageIntLLROutputS3xD(57)(5);
  CNStageIntLLRInputS4xD(97)(0) <= VNStageIntLLROutputS3xD(58)(0);
  CNStageIntLLRInputS4xD(145)(0) <= VNStageIntLLROutputS3xD(58)(1);
  CNStageIntLLRInputS4xD(175)(0) <= VNStageIntLLROutputS3xD(58)(2);
  CNStageIntLLRInputS4xD(312)(0) <= VNStageIntLLROutputS3xD(58)(3);
  CNStageIntLLRInputS4xD(362)(0) <= VNStageIntLLROutputS3xD(58)(4);
  CNStageIntLLRInputS4xD(144)(0) <= VNStageIntLLROutputS3xD(59)(0);
  CNStageIntLLRInputS4xD(174)(0) <= VNStageIntLLROutputS3xD(59)(1);
  CNStageIntLLRInputS4xD(245)(0) <= VNStageIntLLROutputS3xD(59)(2);
  CNStageIntLLRInputS4xD(311)(0) <= VNStageIntLLROutputS3xD(59)(3);
  CNStageIntLLRInputS4xD(361)(0) <= VNStageIntLLROutputS3xD(59)(4);
  CNStageIntLLRInputS4xD(96)(0) <= VNStageIntLLROutputS3xD(60)(0);
  CNStageIntLLRInputS4xD(143)(0) <= VNStageIntLLROutputS3xD(60)(1);
  CNStageIntLLRInputS4xD(173)(0) <= VNStageIntLLROutputS3xD(60)(2);
  CNStageIntLLRInputS4xD(244)(0) <= VNStageIntLLROutputS3xD(60)(3);
  CNStageIntLLRInputS4xD(310)(0) <= VNStageIntLLROutputS3xD(60)(4);
  CNStageIntLLRInputS4xD(360)(0) <= VNStageIntLLROutputS3xD(60)(5);
  CNStageIntLLRInputS4xD(95)(0) <= VNStageIntLLROutputS3xD(61)(0);
  CNStageIntLLRInputS4xD(142)(0) <= VNStageIntLLROutputS3xD(61)(1);
  CNStageIntLLRInputS4xD(172)(0) <= VNStageIntLLROutputS3xD(61)(2);
  CNStageIntLLRInputS4xD(243)(0) <= VNStageIntLLROutputS3xD(61)(3);
  CNStageIntLLRInputS4xD(309)(0) <= VNStageIntLLROutputS3xD(61)(4);
  CNStageIntLLRInputS4xD(359)(0) <= VNStageIntLLROutputS3xD(61)(5);
  CNStageIntLLRInputS4xD(94)(0) <= VNStageIntLLROutputS3xD(62)(0);
  CNStageIntLLRInputS4xD(141)(0) <= VNStageIntLLROutputS3xD(62)(1);
  CNStageIntLLRInputS4xD(171)(0) <= VNStageIntLLROutputS3xD(62)(2);
  CNStageIntLLRInputS4xD(242)(0) <= VNStageIntLLROutputS3xD(62)(3);
  CNStageIntLLRInputS4xD(308)(0) <= VNStageIntLLROutputS3xD(62)(4);
  CNStageIntLLRInputS4xD(358)(0) <= VNStageIntLLROutputS3xD(62)(5);
  CNStageIntLLRInputS4xD(52)(0) <= VNStageIntLLROutputS3xD(63)(0);
  CNStageIntLLRInputS4xD(93)(0) <= VNStageIntLLROutputS3xD(63)(1);
  CNStageIntLLRInputS4xD(140)(0) <= VNStageIntLLROutputS3xD(63)(2);
  CNStageIntLLRInputS4xD(357)(0) <= VNStageIntLLROutputS3xD(63)(3);
  CNStageIntLLRInputS4xD(53)(1) <= VNStageIntLLROutputS3xD(64)(0);
  CNStageIntLLRInputS4xD(109)(1) <= VNStageIntLLROutputS3xD(64)(1);
  CNStageIntLLRInputS4xD(130)(1) <= VNStageIntLLROutputS3xD(64)(2);
  CNStageIntLLRInputS4xD(245)(1) <= VNStageIntLLROutputS3xD(64)(3);
  CNStageIntLLRInputS4xD(299)(1) <= VNStageIntLLROutputS3xD(64)(4);
  CNStageIntLLRInputS4xD(342)(1) <= VNStageIntLLROutputS3xD(64)(5);
  CNStageIntLLRInputS4xD(51)(1) <= VNStageIntLLROutputS3xD(65)(0);
  CNStageIntLLRInputS4xD(74)(1) <= VNStageIntLLROutputS3xD(65)(1);
  CNStageIntLLRInputS4xD(141)(1) <= VNStageIntLLROutputS3xD(65)(2);
  CNStageIntLLRInputS4xD(189)(1) <= VNStageIntLLROutputS3xD(65)(3);
  CNStageIntLLRInputS4xD(286)(1) <= VNStageIntLLROutputS3xD(65)(4);
  CNStageIntLLRInputS4xD(50)(1) <= VNStageIntLLROutputS3xD(66)(0);
  CNStageIntLLRInputS4xD(66)(1) <= VNStageIntLLROutputS3xD(66)(1);
  CNStageIntLLRInputS4xD(155)(1) <= VNStageIntLLROutputS3xD(66)(2);
  CNStageIntLLRInputS4xD(244)(1) <= VNStageIntLLROutputS3xD(66)(3);
  CNStageIntLLRInputS4xD(97)(1) <= VNStageIntLLROutputS3xD(67)(0);
  CNStageIntLLRInputS4xD(275)(1) <= VNStageIntLLROutputS3xD(67)(1);
  CNStageIntLLRInputS4xD(322)(1) <= VNStageIntLLROutputS3xD(67)(2);
  CNStageIntLLRInputS4xD(365)(1) <= VNStageIntLLROutputS3xD(67)(3);
  CNStageIntLLRInputS4xD(49)(1) <= VNStageIntLLROutputS3xD(68)(0);
  CNStageIntLLRInputS4xD(112)(1) <= VNStageIntLLROutputS3xD(68)(1);
  CNStageIntLLRInputS4xD(210)(1) <= VNStageIntLLROutputS3xD(68)(2);
  CNStageIntLLRInputS4xD(256)(1) <= VNStageIntLLROutputS3xD(68)(3);
  CNStageIntLLRInputS4xD(318)(1) <= VNStageIntLLROutputS3xD(68)(4);
  CNStageIntLLRInputS4xD(381)(1) <= VNStageIntLLROutputS3xD(68)(5);
  CNStageIntLLRInputS4xD(48)(1) <= VNStageIntLLROutputS3xD(69)(0);
  CNStageIntLLRInputS4xD(101)(1) <= VNStageIntLLROutputS3xD(69)(1);
  CNStageIntLLRInputS4xD(135)(1) <= VNStageIntLLROutputS3xD(69)(2);
  CNStageIntLLRInputS4xD(215)(1) <= VNStageIntLLROutputS3xD(69)(3);
  CNStageIntLLRInputS4xD(259)(1) <= VNStageIntLLROutputS3xD(69)(4);
  CNStageIntLLRInputS4xD(283)(1) <= VNStageIntLLROutputS3xD(69)(5);
  CNStageIntLLRInputS4xD(351)(1) <= VNStageIntLLROutputS3xD(69)(6);
  CNStageIntLLRInputS4xD(47)(1) <= VNStageIntLLROutputS3xD(70)(0);
  CNStageIntLLRInputS4xD(104)(1) <= VNStageIntLLROutputS3xD(70)(1);
  CNStageIntLLRInputS4xD(136)(1) <= VNStageIntLLROutputS3xD(70)(2);
  CNStageIntLLRInputS4xD(206)(1) <= VNStageIntLLROutputS3xD(70)(3);
  CNStageIntLLRInputS4xD(246)(1) <= VNStageIntLLROutputS3xD(70)(4);
  CNStageIntLLRInputS4xD(301)(1) <= VNStageIntLLROutputS3xD(70)(5);
  CNStageIntLLRInputS4xD(46)(1) <= VNStageIntLLROutputS3xD(71)(0);
  CNStageIntLLRInputS4xD(95)(1) <= VNStageIntLLROutputS3xD(71)(1);
  CNStageIntLLRInputS4xD(176)(1) <= VNStageIntLLROutputS3xD(71)(2);
  CNStageIntLLRInputS4xD(276)(1) <= VNStageIntLLROutputS3xD(71)(3);
  CNStageIntLLRInputS4xD(302)(1) <= VNStageIntLLROutputS3xD(71)(4);
  CNStageIntLLRInputS4xD(353)(1) <= VNStageIntLLROutputS3xD(71)(5);
  CNStageIntLLRInputS4xD(45)(1) <= VNStageIntLLROutputS3xD(72)(0);
  CNStageIntLLRInputS4xD(75)(1) <= VNStageIntLLROutputS3xD(72)(1);
  CNStageIntLLRInputS4xD(162)(1) <= VNStageIntLLROutputS3xD(72)(2);
  CNStageIntLLRInputS4xD(183)(1) <= VNStageIntLLROutputS3xD(72)(3);
  CNStageIntLLRInputS4xD(243)(1) <= VNStageIntLLROutputS3xD(72)(4);
  CNStageIntLLRInputS4xD(367)(1) <= VNStageIntLLROutputS3xD(72)(5);
  CNStageIntLLRInputS4xD(44)(1) <= VNStageIntLLROutputS3xD(73)(0);
  CNStageIntLLRInputS4xD(56)(1) <= VNStageIntLLROutputS3xD(73)(1);
  CNStageIntLLRInputS4xD(121)(1) <= VNStageIntLLROutputS3xD(73)(2);
  CNStageIntLLRInputS4xD(219)(1) <= VNStageIntLLROutputS3xD(73)(3);
  CNStageIntLLRInputS4xD(328)(1) <= VNStageIntLLROutputS3xD(73)(4);
  CNStageIntLLRInputS4xD(363)(1) <= VNStageIntLLROutputS3xD(73)(5);
  CNStageIntLLRInputS4xD(43)(1) <= VNStageIntLLROutputS3xD(74)(0);
  CNStageIntLLRInputS4xD(70)(1) <= VNStageIntLLROutputS3xD(74)(1);
  CNStageIntLLRInputS4xD(125)(1) <= VNStageIntLLROutputS3xD(74)(2);
  CNStageIntLLRInputS4xD(221)(1) <= VNStageIntLLROutputS3xD(74)(3);
  CNStageIntLLRInputS4xD(290)(1) <= VNStageIntLLROutputS3xD(74)(4);
  CNStageIntLLRInputS4xD(42)(1) <= VNStageIntLLROutputS3xD(75)(0);
  CNStageIntLLRInputS4xD(81)(1) <= VNStageIntLLROutputS3xD(75)(1);
  CNStageIntLLRInputS4xD(170)(1) <= VNStageIntLLROutputS3xD(75)(2);
  CNStageIntLLRInputS4xD(192)(1) <= VNStageIntLLROutputS3xD(75)(3);
  CNStageIntLLRInputS4xD(278)(1) <= VNStageIntLLROutputS3xD(75)(4);
  CNStageIntLLRInputS4xD(294)(1) <= VNStageIntLLROutputS3xD(75)(5);
  CNStageIntLLRInputS4xD(347)(1) <= VNStageIntLLROutputS3xD(75)(6);
  CNStageIntLLRInputS4xD(41)(1) <= VNStageIntLLROutputS3xD(76)(0);
  CNStageIntLLRInputS4xD(106)(1) <= VNStageIntLLROutputS3xD(76)(1);
  CNStageIntLLRInputS4xD(124)(1) <= VNStageIntLLROutputS3xD(76)(2);
  CNStageIntLLRInputS4xD(174)(1) <= VNStageIntLLROutputS3xD(76)(3);
  CNStageIntLLRInputS4xD(270)(1) <= VNStageIntLLROutputS3xD(76)(4);
  CNStageIntLLRInputS4xD(332)(1) <= VNStageIntLLROutputS3xD(76)(5);
  CNStageIntLLRInputS4xD(348)(1) <= VNStageIntLLROutputS3xD(76)(6);
  CNStageIntLLRInputS4xD(119)(1) <= VNStageIntLLROutputS3xD(77)(0);
  CNStageIntLLRInputS4xD(185)(1) <= VNStageIntLLROutputS3xD(77)(1);
  CNStageIntLLRInputS4xD(257)(1) <= VNStageIntLLROutputS3xD(77)(2);
  CNStageIntLLRInputS4xD(293)(1) <= VNStageIntLLROutputS3xD(77)(3);
  CNStageIntLLRInputS4xD(383)(1) <= VNStageIntLLROutputS3xD(77)(4);
  CNStageIntLLRInputS4xD(40)(1) <= VNStageIntLLROutputS3xD(78)(0);
  CNStageIntLLRInputS4xD(84)(1) <= VNStageIntLLROutputS3xD(78)(1);
  CNStageIntLLRInputS4xD(159)(1) <= VNStageIntLLROutputS3xD(78)(2);
  CNStageIntLLRInputS4xD(193)(1) <= VNStageIntLLROutputS3xD(78)(3);
  CNStageIntLLRInputS4xD(274)(1) <= VNStageIntLLROutputS3xD(78)(4);
  CNStageIntLLRInputS4xD(288)(1) <= VNStageIntLLROutputS3xD(78)(5);
  CNStageIntLLRInputS4xD(374)(1) <= VNStageIntLLROutputS3xD(78)(6);
  CNStageIntLLRInputS4xD(39)(1) <= VNStageIntLLROutputS3xD(79)(0);
  CNStageIntLLRInputS4xD(99)(1) <= VNStageIntLLROutputS3xD(79)(1);
  CNStageIntLLRInputS4xD(167)(1) <= VNStageIntLLROutputS3xD(79)(2);
  CNStageIntLLRInputS4xD(220)(1) <= VNStageIntLLROutputS3xD(79)(3);
  CNStageIntLLRInputS4xD(325)(1) <= VNStageIntLLROutputS3xD(79)(4);
  CNStageIntLLRInputS4xD(38)(1) <= VNStageIntLLROutputS3xD(80)(0);
  CNStageIntLLRInputS4xD(62)(1) <= VNStageIntLLROutputS3xD(80)(1);
  CNStageIntLLRInputS4xD(131)(1) <= VNStageIntLLROutputS3xD(80)(2);
  CNStageIntLLRInputS4xD(182)(1) <= VNStageIntLLROutputS3xD(80)(3);
  CNStageIntLLRInputS4xD(248)(1) <= VNStageIntLLROutputS3xD(80)(4);
  CNStageIntLLRInputS4xD(337)(1) <= VNStageIntLLROutputS3xD(80)(5);
  CNStageIntLLRInputS4xD(37)(1) <= VNStageIntLLROutputS3xD(81)(0);
  CNStageIntLLRInputS4xD(72)(1) <= VNStageIntLLROutputS3xD(81)(1);
  CNStageIntLLRInputS4xD(129)(1) <= VNStageIntLLROutputS3xD(81)(2);
  CNStageIntLLRInputS4xD(262)(1) <= VNStageIntLLROutputS3xD(81)(3);
  CNStageIntLLRInputS4xD(36)(1) <= VNStageIntLLROutputS3xD(82)(0);
  CNStageIntLLRInputS4xD(67)(1) <= VNStageIntLLROutputS3xD(82)(1);
  CNStageIntLLRInputS4xD(165)(1) <= VNStageIntLLROutputS3xD(82)(2);
  CNStageIntLLRInputS4xD(188)(1) <= VNStageIntLLROutputS3xD(82)(3);
  CNStageIntLLRInputS4xD(254)(1) <= VNStageIntLLROutputS3xD(82)(4);
  CNStageIntLLRInputS4xD(298)(1) <= VNStageIntLLROutputS3xD(82)(5);
  CNStageIntLLRInputS4xD(336)(1) <= VNStageIntLLROutputS3xD(82)(6);
  CNStageIntLLRInputS4xD(35)(1) <= VNStageIntLLROutputS3xD(83)(0);
  CNStageIntLLRInputS4xD(73)(1) <= VNStageIntLLROutputS3xD(83)(1);
  CNStageIntLLRInputS4xD(144)(1) <= VNStageIntLLROutputS3xD(83)(2);
  CNStageIntLLRInputS4xD(208)(1) <= VNStageIntLLROutputS3xD(83)(3);
  CNStageIntLLRInputS4xD(232)(1) <= VNStageIntLLROutputS3xD(83)(4);
  CNStageIntLLRInputS4xD(330)(1) <= VNStageIntLLROutputS3xD(83)(5);
  CNStageIntLLRInputS4xD(34)(1) <= VNStageIntLLROutputS3xD(84)(0);
  CNStageIntLLRInputS4xD(61)(1) <= VNStageIntLLROutputS3xD(84)(1);
  CNStageIntLLRInputS4xD(147)(1) <= VNStageIntLLROutputS3xD(84)(2);
  CNStageIntLLRInputS4xD(222)(1) <= VNStageIntLLROutputS3xD(84)(3);
  CNStageIntLLRInputS4xD(310)(1) <= VNStageIntLLROutputS3xD(84)(4);
  CNStageIntLLRInputS4xD(371)(1) <= VNStageIntLLROutputS3xD(84)(5);
  CNStageIntLLRInputS4xD(33)(1) <= VNStageIntLLROutputS3xD(85)(0);
  CNStageIntLLRInputS4xD(132)(1) <= VNStageIntLLROutputS3xD(85)(1);
  CNStageIntLLRInputS4xD(218)(1) <= VNStageIntLLROutputS3xD(85)(2);
  CNStageIntLLRInputS4xD(235)(1) <= VNStageIntLLROutputS3xD(85)(3);
  CNStageIntLLRInputS4xD(313)(1) <= VNStageIntLLROutputS3xD(85)(4);
  CNStageIntLLRInputS4xD(379)(1) <= VNStageIntLLROutputS3xD(85)(5);
  CNStageIntLLRInputS4xD(32)(1) <= VNStageIntLLROutputS3xD(86)(0);
  CNStageIntLLRInputS4xD(166)(1) <= VNStageIntLLROutputS3xD(86)(1);
  CNStageIntLLRInputS4xD(239)(1) <= VNStageIntLLROutputS3xD(86)(2);
  CNStageIntLLRInputS4xD(343)(1) <= VNStageIntLLROutputS3xD(86)(3);
  CNStageIntLLRInputS4xD(31)(1) <= VNStageIntLLROutputS3xD(87)(0);
  CNStageIntLLRInputS4xD(77)(1) <= VNStageIntLLROutputS3xD(87)(1);
  CNStageIntLLRInputS4xD(128)(1) <= VNStageIntLLROutputS3xD(87)(2);
  CNStageIntLLRInputS4xD(203)(1) <= VNStageIntLLROutputS3xD(87)(3);
  CNStageIntLLRInputS4xD(229)(1) <= VNStageIntLLROutputS3xD(87)(4);
  CNStageIntLLRInputS4xD(331)(1) <= VNStageIntLLROutputS3xD(87)(5);
  CNStageIntLLRInputS4xD(341)(1) <= VNStageIntLLROutputS3xD(87)(6);
  CNStageIntLLRInputS4xD(30)(1) <= VNStageIntLLROutputS3xD(88)(0);
  CNStageIntLLRInputS4xD(79)(1) <= VNStageIntLLROutputS3xD(88)(1);
  CNStageIntLLRInputS4xD(156)(1) <= VNStageIntLLROutputS3xD(88)(2);
  CNStageIntLLRInputS4xD(204)(1) <= VNStageIntLLROutputS3xD(88)(3);
  CNStageIntLLRInputS4xD(263)(1) <= VNStageIntLLROutputS3xD(88)(4);
  CNStageIntLLRInputS4xD(297)(1) <= VNStageIntLLROutputS3xD(88)(5);
  CNStageIntLLRInputS4xD(377)(1) <= VNStageIntLLROutputS3xD(88)(6);
  CNStageIntLLRInputS4xD(29)(1) <= VNStageIntLLROutputS3xD(89)(0);
  CNStageIntLLRInputS4xD(102)(1) <= VNStageIntLLROutputS3xD(89)(1);
  CNStageIntLLRInputS4xD(140)(1) <= VNStageIntLLROutputS3xD(89)(2);
  CNStageIntLLRInputS4xD(184)(1) <= VNStageIntLLROutputS3xD(89)(3);
  CNStageIntLLRInputS4xD(247)(1) <= VNStageIntLLROutputS3xD(89)(4);
  CNStageIntLLRInputS4xD(355)(1) <= VNStageIntLLROutputS3xD(89)(5);
  CNStageIntLLRInputS4xD(28)(1) <= VNStageIntLLROutputS3xD(90)(0);
  CNStageIntLLRInputS4xD(85)(1) <= VNStageIntLLROutputS3xD(90)(1);
  CNStageIntLLRInputS4xD(168)(1) <= VNStageIntLLROutputS3xD(90)(2);
  CNStageIntLLRInputS4xD(175)(1) <= VNStageIntLLROutputS3xD(90)(3);
  CNStageIntLLRInputS4xD(258)(1) <= VNStageIntLLROutputS3xD(90)(4);
  CNStageIntLLRInputS4xD(307)(1) <= VNStageIntLLROutputS3xD(90)(5);
  CNStageIntLLRInputS4xD(358)(1) <= VNStageIntLLROutputS3xD(90)(6);
  CNStageIntLLRInputS4xD(27)(1) <= VNStageIntLLROutputS3xD(91)(0);
  CNStageIntLLRInputS4xD(96)(1) <= VNStageIntLLROutputS3xD(91)(1);
  CNStageIntLLRInputS4xD(158)(1) <= VNStageIntLLROutputS3xD(91)(2);
  CNStageIntLLRInputS4xD(191)(1) <= VNStageIntLLROutputS3xD(91)(3);
  CNStageIntLLRInputS4xD(269)(1) <= VNStageIntLLROutputS3xD(91)(4);
  CNStageIntLLRInputS4xD(280)(1) <= VNStageIntLLROutputS3xD(91)(5);
  CNStageIntLLRInputS4xD(344)(1) <= VNStageIntLLROutputS3xD(91)(6);
  CNStageIntLLRInputS4xD(26)(1) <= VNStageIntLLROutputS3xD(92)(0);
  CNStageIntLLRInputS4xD(103)(1) <= VNStageIntLLROutputS3xD(92)(1);
  CNStageIntLLRInputS4xD(145)(1) <= VNStageIntLLROutputS3xD(92)(2);
  CNStageIntLLRInputS4xD(195)(1) <= VNStageIntLLROutputS3xD(92)(3);
  CNStageIntLLRInputS4xD(242)(1) <= VNStageIntLLROutputS3xD(92)(4);
  CNStageIntLLRInputS4xD(324)(1) <= VNStageIntLLROutputS3xD(92)(5);
  CNStageIntLLRInputS4xD(378)(1) <= VNStageIntLLROutputS3xD(92)(6);
  CNStageIntLLRInputS4xD(25)(1) <= VNStageIntLLROutputS3xD(93)(0);
  CNStageIntLLRInputS4xD(78)(1) <= VNStageIntLLROutputS3xD(93)(1);
  CNStageIntLLRInputS4xD(164)(1) <= VNStageIntLLROutputS3xD(93)(2);
  CNStageIntLLRInputS4xD(224)(1) <= VNStageIntLLROutputS3xD(93)(3);
  CNStageIntLLRInputS4xD(231)(1) <= VNStageIntLLROutputS3xD(93)(4);
  CNStageIntLLRInputS4xD(311)(1) <= VNStageIntLLROutputS3xD(93)(5);
  CNStageIntLLRInputS4xD(340)(1) <= VNStageIntLLROutputS3xD(93)(6);
  CNStageIntLLRInputS4xD(24)(1) <= VNStageIntLLROutputS3xD(94)(0);
  CNStageIntLLRInputS4xD(92)(1) <= VNStageIntLLROutputS3xD(94)(1);
  CNStageIntLLRInputS4xD(194)(1) <= VNStageIntLLROutputS3xD(94)(2);
  CNStageIntLLRInputS4xD(329)(1) <= VNStageIntLLROutputS3xD(94)(3);
  CNStageIntLLRInputS4xD(368)(1) <= VNStageIntLLROutputS3xD(94)(4);
  CNStageIntLLRInputS4xD(23)(1) <= VNStageIntLLROutputS3xD(95)(0);
  CNStageIntLLRInputS4xD(63)(1) <= VNStageIntLLROutputS3xD(95)(1);
  CNStageIntLLRInputS4xD(134)(1) <= VNStageIntLLROutputS3xD(95)(2);
  CNStageIntLLRInputS4xD(190)(1) <= VNStageIntLLROutputS3xD(95)(3);
  CNStageIntLLRInputS4xD(234)(1) <= VNStageIntLLROutputS3xD(95)(4);
  CNStageIntLLRInputS4xD(303)(1) <= VNStageIntLLROutputS3xD(95)(5);
  CNStageIntLLRInputS4xD(352)(1) <= VNStageIntLLROutputS3xD(95)(6);
  CNStageIntLLRInputS4xD(22)(1) <= VNStageIntLLROutputS3xD(96)(0);
  CNStageIntLLRInputS4xD(98)(1) <= VNStageIntLLROutputS3xD(96)(1);
  CNStageIntLLRInputS4xD(150)(1) <= VNStageIntLLROutputS3xD(96)(2);
  CNStageIntLLRInputS4xD(172)(1) <= VNStageIntLLROutputS3xD(96)(3);
  CNStageIntLLRInputS4xD(251)(1) <= VNStageIntLLROutputS3xD(96)(4);
  CNStageIntLLRInputS4xD(380)(1) <= VNStageIntLLROutputS3xD(96)(5);
  CNStageIntLLRInputS4xD(21)(1) <= VNStageIntLLROutputS3xD(97)(0);
  CNStageIntLLRInputS4xD(65)(1) <= VNStageIntLLROutputS3xD(97)(1);
  CNStageIntLLRInputS4xD(142)(1) <= VNStageIntLLROutputS3xD(97)(2);
  CNStageIntLLRInputS4xD(180)(1) <= VNStageIntLLROutputS3xD(97)(3);
  CNStageIntLLRInputS4xD(260)(1) <= VNStageIntLLROutputS3xD(97)(4);
  CNStageIntLLRInputS4xD(316)(1) <= VNStageIntLLROutputS3xD(97)(5);
  CNStageIntLLRInputS4xD(370)(1) <= VNStageIntLLROutputS3xD(97)(6);
  CNStageIntLLRInputS4xD(20)(1) <= VNStageIntLLROutputS3xD(98)(0);
  CNStageIntLLRInputS4xD(116)(1) <= VNStageIntLLROutputS3xD(98)(1);
  CNStageIntLLRInputS4xD(199)(1) <= VNStageIntLLROutputS3xD(98)(2);
  CNStageIntLLRInputS4xD(255)(1) <= VNStageIntLLROutputS3xD(98)(3);
  CNStageIntLLRInputS4xD(308)(1) <= VNStageIntLLROutputS3xD(98)(4);
  CNStageIntLLRInputS4xD(356)(1) <= VNStageIntLLROutputS3xD(98)(5);
  CNStageIntLLRInputS4xD(19)(1) <= VNStageIntLLROutputS3xD(99)(0);
  CNStageIntLLRInputS4xD(76)(1) <= VNStageIntLLROutputS3xD(99)(1);
  CNStageIntLLRInputS4xD(126)(1) <= VNStageIntLLROutputS3xD(99)(2);
  CNStageIntLLRInputS4xD(198)(1) <= VNStageIntLLROutputS3xD(99)(3);
  CNStageIntLLRInputS4xD(261)(1) <= VNStageIntLLROutputS3xD(99)(4);
  CNStageIntLLRInputS4xD(285)(1) <= VNStageIntLLROutputS3xD(99)(5);
  CNStageIntLLRInputS4xD(376)(1) <= VNStageIntLLROutputS3xD(99)(6);
  CNStageIntLLRInputS4xD(18)(1) <= VNStageIntLLROutputS3xD(100)(0);
  CNStageIntLLRInputS4xD(94)(1) <= VNStageIntLLROutputS3xD(100)(1);
  CNStageIntLLRInputS4xD(120)(1) <= VNStageIntLLROutputS3xD(100)(2);
  CNStageIntLLRInputS4xD(178)(1) <= VNStageIntLLROutputS3xD(100)(3);
  CNStageIntLLRInputS4xD(250)(1) <= VNStageIntLLROutputS3xD(100)(4);
  CNStageIntLLRInputS4xD(295)(1) <= VNStageIntLLROutputS3xD(100)(5);
  CNStageIntLLRInputS4xD(349)(1) <= VNStageIntLLROutputS3xD(100)(6);
  CNStageIntLLRInputS4xD(17)(1) <= VNStageIntLLROutputS3xD(101)(0);
  CNStageIntLLRInputS4xD(58)(1) <= VNStageIntLLROutputS3xD(101)(1);
  CNStageIntLLRInputS4xD(123)(1) <= VNStageIntLLROutputS3xD(101)(2);
  CNStageIntLLRInputS4xD(211)(1) <= VNStageIntLLROutputS3xD(101)(3);
  CNStageIntLLRInputS4xD(273)(1) <= VNStageIntLLROutputS3xD(101)(4);
  CNStageIntLLRInputS4xD(289)(1) <= VNStageIntLLROutputS3xD(101)(5);
  CNStageIntLLRInputS4xD(346)(1) <= VNStageIntLLROutputS3xD(101)(6);
  CNStageIntLLRInputS4xD(16)(1) <= VNStageIntLLROutputS3xD(102)(0);
  CNStageIntLLRInputS4xD(59)(1) <= VNStageIntLLROutputS3xD(102)(1);
  CNStageIntLLRInputS4xD(113)(1) <= VNStageIntLLROutputS3xD(102)(2);
  CNStageIntLLRInputS4xD(214)(1) <= VNStageIntLLROutputS3xD(102)(3);
  CNStageIntLLRInputS4xD(226)(1) <= VNStageIntLLROutputS3xD(102)(4);
  CNStageIntLLRInputS4xD(361)(1) <= VNStageIntLLROutputS3xD(102)(5);
  CNStageIntLLRInputS4xD(15)(1) <= VNStageIntLLROutputS3xD(103)(0);
  CNStageIntLLRInputS4xD(93)(1) <= VNStageIntLLROutputS3xD(103)(1);
  CNStageIntLLRInputS4xD(151)(1) <= VNStageIntLLROutputS3xD(103)(2);
  CNStageIntLLRInputS4xD(200)(1) <= VNStageIntLLROutputS3xD(103)(3);
  CNStageIntLLRInputS4xD(265)(1) <= VNStageIntLLROutputS3xD(103)(4);
  CNStageIntLLRInputS4xD(284)(1) <= VNStageIntLLROutputS3xD(103)(5);
  CNStageIntLLRInputS4xD(354)(1) <= VNStageIntLLROutputS3xD(103)(6);
  CNStageIntLLRInputS4xD(14)(1) <= VNStageIntLLROutputS3xD(104)(0);
  CNStageIntLLRInputS4xD(86)(1) <= VNStageIntLLROutputS3xD(104)(1);
  CNStageIntLLRInputS4xD(133)(1) <= VNStageIntLLROutputS3xD(104)(2);
  CNStageIntLLRInputS4xD(179)(1) <= VNStageIntLLROutputS3xD(104)(3);
  CNStageIntLLRInputS4xD(267)(1) <= VNStageIntLLROutputS3xD(104)(4);
  CNStageIntLLRInputS4xD(317)(1) <= VNStageIntLLROutputS3xD(104)(5);
  CNStageIntLLRInputS4xD(13)(1) <= VNStageIntLLROutputS3xD(105)(0);
  CNStageIntLLRInputS4xD(146)(1) <= VNStageIntLLROutputS3xD(105)(1);
  CNStageIntLLRInputS4xD(197)(1) <= VNStageIntLLROutputS3xD(105)(2);
  CNStageIntLLRInputS4xD(237)(1) <= VNStageIntLLROutputS3xD(105)(3);
  CNStageIntLLRInputS4xD(300)(1) <= VNStageIntLLROutputS3xD(105)(4);
  CNStageIntLLRInputS4xD(338)(1) <= VNStageIntLLROutputS3xD(105)(5);
  CNStageIntLLRInputS4xD(12)(1) <= VNStageIntLLROutputS3xD(106)(0);
  CNStageIntLLRInputS4xD(157)(1) <= VNStageIntLLROutputS3xD(106)(1);
  CNStageIntLLRInputS4xD(223)(1) <= VNStageIntLLROutputS3xD(106)(2);
  CNStageIntLLRInputS4xD(272)(1) <= VNStageIntLLROutputS3xD(106)(3);
  CNStageIntLLRInputS4xD(312)(1) <= VNStageIntLLROutputS3xD(106)(4);
  CNStageIntLLRInputS4xD(333)(1) <= VNStageIntLLROutputS3xD(106)(5);
  CNStageIntLLRInputS4xD(110)(1) <= VNStageIntLLROutputS3xD(107)(0);
  CNStageIntLLRInputS4xD(127)(1) <= VNStageIntLLROutputS3xD(107)(1);
  CNStageIntLLRInputS4xD(207)(1) <= VNStageIntLLROutputS3xD(107)(2);
  CNStageIntLLRInputS4xD(230)(1) <= VNStageIntLLROutputS3xD(107)(3);
  CNStageIntLLRInputS4xD(323)(1) <= VNStageIntLLROutputS3xD(107)(4);
  CNStageIntLLRInputS4xD(335)(1) <= VNStageIntLLROutputS3xD(107)(5);
  CNStageIntLLRInputS4xD(11)(1) <= VNStageIntLLROutputS3xD(108)(0);
  CNStageIntLLRInputS4xD(105)(1) <= VNStageIntLLROutputS3xD(108)(1);
  CNStageIntLLRInputS4xD(115)(1) <= VNStageIntLLROutputS3xD(108)(2);
  CNStageIntLLRInputS4xD(181)(1) <= VNStageIntLLROutputS3xD(108)(3);
  CNStageIntLLRInputS4xD(238)(1) <= VNStageIntLLROutputS3xD(108)(4);
  CNStageIntLLRInputS4xD(296)(1) <= VNStageIntLLROutputS3xD(108)(5);
  CNStageIntLLRInputS4xD(10)(1) <= VNStageIntLLROutputS3xD(109)(0);
  CNStageIntLLRInputS4xD(100)(1) <= VNStageIntLLROutputS3xD(109)(1);
  CNStageIntLLRInputS4xD(160)(1) <= VNStageIntLLROutputS3xD(109)(2);
  CNStageIntLLRInputS4xD(171)(1) <= VNStageIntLLROutputS3xD(109)(3);
  CNStageIntLLRInputS4xD(266)(1) <= VNStageIntLLROutputS3xD(109)(4);
  CNStageIntLLRInputS4xD(362)(1) <= VNStageIntLLROutputS3xD(109)(5);
  CNStageIntLLRInputS4xD(9)(1) <= VNStageIntLLROutputS3xD(110)(0);
  CNStageIntLLRInputS4xD(83)(1) <= VNStageIntLLROutputS3xD(110)(1);
  CNStageIntLLRInputS4xD(118)(1) <= VNStageIntLLROutputS3xD(110)(2);
  CNStageIntLLRInputS4xD(212)(1) <= VNStageIntLLROutputS3xD(110)(3);
  CNStageIntLLRInputS4xD(225)(1) <= VNStageIntLLROutputS3xD(110)(4);
  CNStageIntLLRInputS4xD(326)(1) <= VNStageIntLLROutputS3xD(110)(5);
  CNStageIntLLRInputS4xD(345)(1) <= VNStageIntLLROutputS3xD(110)(6);
  CNStageIntLLRInputS4xD(8)(1) <= VNStageIntLLROutputS3xD(111)(0);
  CNStageIntLLRInputS4xD(90)(1) <= VNStageIntLLROutputS3xD(111)(1);
  CNStageIntLLRInputS4xD(138)(1) <= VNStageIntLLROutputS3xD(111)(2);
  CNStageIntLLRInputS4xD(177)(1) <= VNStageIntLLROutputS3xD(111)(3);
  CNStageIntLLRInputS4xD(252)(1) <= VNStageIntLLROutputS3xD(111)(4);
  CNStageIntLLRInputS4xD(287)(1) <= VNStageIntLLROutputS3xD(111)(5);
  CNStageIntLLRInputS4xD(357)(1) <= VNStageIntLLROutputS3xD(111)(6);
  CNStageIntLLRInputS4xD(7)(1) <= VNStageIntLLROutputS3xD(112)(0);
  CNStageIntLLRInputS4xD(54)(1) <= VNStageIntLLROutputS3xD(112)(1);
  CNStageIntLLRInputS4xD(148)(1) <= VNStageIntLLROutputS3xD(112)(2);
  CNStageIntLLRInputS4xD(205)(1) <= VNStageIntLLROutputS3xD(112)(3);
  CNStageIntLLRInputS4xD(233)(1) <= VNStageIntLLROutputS3xD(112)(4);
  CNStageIntLLRInputS4xD(305)(1) <= VNStageIntLLROutputS3xD(112)(5);
  CNStageIntLLRInputS4xD(369)(1) <= VNStageIntLLROutputS3xD(112)(6);
  CNStageIntLLRInputS4xD(6)(1) <= VNStageIntLLROutputS3xD(113)(0);
  CNStageIntLLRInputS4xD(108)(1) <= VNStageIntLLROutputS3xD(113)(1);
  CNStageIntLLRInputS4xD(143)(1) <= VNStageIntLLROutputS3xD(113)(2);
  CNStageIntLLRInputS4xD(202)(1) <= VNStageIntLLROutputS3xD(113)(3);
  CNStageIntLLRInputS4xD(253)(1) <= VNStageIntLLROutputS3xD(113)(4);
  CNStageIntLLRInputS4xD(314)(1) <= VNStageIntLLROutputS3xD(113)(5);
  CNStageIntLLRInputS4xD(339)(1) <= VNStageIntLLROutputS3xD(113)(6);
  CNStageIntLLRInputS4xD(5)(1) <= VNStageIntLLROutputS3xD(114)(0);
  CNStageIntLLRInputS4xD(88)(1) <= VNStageIntLLROutputS3xD(114)(1);
  CNStageIntLLRInputS4xD(149)(1) <= VNStageIntLLROutputS3xD(114)(2);
  CNStageIntLLRInputS4xD(216)(1) <= VNStageIntLLROutputS3xD(114)(3);
  CNStageIntLLRInputS4xD(268)(1) <= VNStageIntLLROutputS3xD(114)(4);
  CNStageIntLLRInputS4xD(309)(1) <= VNStageIntLLROutputS3xD(114)(5);
  CNStageIntLLRInputS4xD(4)(1) <= VNStageIntLLROutputS3xD(115)(0);
  CNStageIntLLRInputS4xD(68)(1) <= VNStageIntLLROutputS3xD(115)(1);
  CNStageIntLLRInputS4xD(137)(1) <= VNStageIntLLROutputS3xD(115)(2);
  CNStageIntLLRInputS4xD(209)(1) <= VNStageIntLLROutputS3xD(115)(3);
  CNStageIntLLRInputS4xD(264)(1) <= VNStageIntLLROutputS3xD(115)(4);
  CNStageIntLLRInputS4xD(315)(1) <= VNStageIntLLROutputS3xD(115)(5);
  CNStageIntLLRInputS4xD(372)(1) <= VNStageIntLLROutputS3xD(115)(6);
  CNStageIntLLRInputS4xD(71)(1) <= VNStageIntLLROutputS3xD(116)(0);
  CNStageIntLLRInputS4xD(163)(1) <= VNStageIntLLROutputS3xD(116)(1);
  CNStageIntLLRInputS4xD(187)(1) <= VNStageIntLLROutputS3xD(116)(2);
  CNStageIntLLRInputS4xD(228)(1) <= VNStageIntLLROutputS3xD(116)(3);
  CNStageIntLLRInputS4xD(304)(1) <= VNStageIntLLROutputS3xD(116)(4);
  CNStageIntLLRInputS4xD(3)(1) <= VNStageIntLLROutputS3xD(117)(0);
  CNStageIntLLRInputS4xD(55)(1) <= VNStageIntLLROutputS3xD(117)(1);
  CNStageIntLLRInputS4xD(111)(1) <= VNStageIntLLROutputS3xD(117)(2);
  CNStageIntLLRInputS4xD(196)(1) <= VNStageIntLLROutputS3xD(117)(3);
  CNStageIntLLRInputS4xD(2)(1) <= VNStageIntLLROutputS3xD(118)(0);
  CNStageIntLLRInputS4xD(89)(1) <= VNStageIntLLROutputS3xD(118)(1);
  CNStageIntLLRInputS4xD(152)(1) <= VNStageIntLLROutputS3xD(118)(2);
  CNStageIntLLRInputS4xD(249)(1) <= VNStageIntLLROutputS3xD(118)(3);
  CNStageIntLLRInputS4xD(282)(1) <= VNStageIntLLROutputS3xD(118)(4);
  CNStageIntLLRInputS4xD(359)(1) <= VNStageIntLLROutputS3xD(118)(5);
  CNStageIntLLRInputS4xD(1)(1) <= VNStageIntLLROutputS3xD(119)(0);
  CNStageIntLLRInputS4xD(107)(1) <= VNStageIntLLROutputS3xD(119)(1);
  CNStageIntLLRInputS4xD(154)(1) <= VNStageIntLLROutputS3xD(119)(2);
  CNStageIntLLRInputS4xD(227)(1) <= VNStageIntLLROutputS3xD(119)(3);
  CNStageIntLLRInputS4xD(319)(1) <= VNStageIntLLROutputS3xD(119)(4);
  CNStageIntLLRInputS4xD(0)(1) <= VNStageIntLLROutputS3xD(120)(0);
  CNStageIntLLRInputS4xD(80)(1) <= VNStageIntLLROutputS3xD(120)(1);
  CNStageIntLLRInputS4xD(321)(1) <= VNStageIntLLROutputS3xD(120)(2);
  CNStageIntLLRInputS4xD(360)(1) <= VNStageIntLLROutputS3xD(120)(3);
  CNStageIntLLRInputS4xD(64)(1) <= VNStageIntLLROutputS3xD(121)(0);
  CNStageIntLLRInputS4xD(161)(1) <= VNStageIntLLROutputS3xD(121)(1);
  CNStageIntLLRInputS4xD(217)(1) <= VNStageIntLLROutputS3xD(121)(2);
  CNStageIntLLRInputS4xD(236)(1) <= VNStageIntLLROutputS3xD(121)(3);
  CNStageIntLLRInputS4xD(291)(1) <= VNStageIntLLROutputS3xD(121)(4);
  CNStageIntLLRInputS4xD(350)(1) <= VNStageIntLLROutputS3xD(121)(5);
  CNStageIntLLRInputS4xD(91)(1) <= VNStageIntLLROutputS3xD(122)(0);
  CNStageIntLLRInputS4xD(114)(1) <= VNStageIntLLROutputS3xD(122)(1);
  CNStageIntLLRInputS4xD(201)(1) <= VNStageIntLLROutputS3xD(122)(2);
  CNStageIntLLRInputS4xD(241)(1) <= VNStageIntLLROutputS3xD(122)(3);
  CNStageIntLLRInputS4xD(327)(1) <= VNStageIntLLROutputS3xD(122)(4);
  CNStageIntLLRInputS4xD(375)(1) <= VNStageIntLLROutputS3xD(122)(5);
  CNStageIntLLRInputS4xD(82)(1) <= VNStageIntLLROutputS3xD(123)(0);
  CNStageIntLLRInputS4xD(122)(1) <= VNStageIntLLROutputS3xD(123)(1);
  CNStageIntLLRInputS4xD(213)(1) <= VNStageIntLLROutputS3xD(123)(2);
  CNStageIntLLRInputS4xD(279)(1) <= VNStageIntLLROutputS3xD(123)(3);
  CNStageIntLLRInputS4xD(382)(1) <= VNStageIntLLROutputS3xD(123)(4);
  CNStageIntLLRInputS4xD(69)(1) <= VNStageIntLLROutputS3xD(124)(0);
  CNStageIntLLRInputS4xD(153)(1) <= VNStageIntLLROutputS3xD(124)(1);
  CNStageIntLLRInputS4xD(240)(1) <= VNStageIntLLROutputS3xD(124)(2);
  CNStageIntLLRInputS4xD(292)(1) <= VNStageIntLLROutputS3xD(124)(3);
  CNStageIntLLRInputS4xD(364)(1) <= VNStageIntLLROutputS3xD(124)(4);
  CNStageIntLLRInputS4xD(87)(1) <= VNStageIntLLROutputS3xD(125)(0);
  CNStageIntLLRInputS4xD(169)(1) <= VNStageIntLLROutputS3xD(125)(1);
  CNStageIntLLRInputS4xD(320)(1) <= VNStageIntLLROutputS3xD(125)(2);
  CNStageIntLLRInputS4xD(366)(1) <= VNStageIntLLROutputS3xD(125)(3);
  CNStageIntLLRInputS4xD(60)(1) <= VNStageIntLLROutputS3xD(126)(0);
  CNStageIntLLRInputS4xD(139)(1) <= VNStageIntLLROutputS3xD(126)(1);
  CNStageIntLLRInputS4xD(186)(1) <= VNStageIntLLROutputS3xD(126)(2);
  CNStageIntLLRInputS4xD(271)(1) <= VNStageIntLLROutputS3xD(126)(3);
  CNStageIntLLRInputS4xD(281)(1) <= VNStageIntLLROutputS3xD(126)(4);
  CNStageIntLLRInputS4xD(334)(1) <= VNStageIntLLROutputS3xD(126)(5);
  CNStageIntLLRInputS4xD(52)(1) <= VNStageIntLLROutputS3xD(127)(0);
  CNStageIntLLRInputS4xD(57)(1) <= VNStageIntLLROutputS3xD(127)(1);
  CNStageIntLLRInputS4xD(117)(1) <= VNStageIntLLROutputS3xD(127)(2);
  CNStageIntLLRInputS4xD(173)(1) <= VNStageIntLLROutputS3xD(127)(3);
  CNStageIntLLRInputS4xD(277)(1) <= VNStageIntLLROutputS3xD(127)(4);
  CNStageIntLLRInputS4xD(306)(1) <= VNStageIntLLROutputS3xD(127)(5);
  CNStageIntLLRInputS4xD(373)(1) <= VNStageIntLLROutputS3xD(127)(6);
  CNStageIntLLRInputS4xD(53)(2) <= VNStageIntLLROutputS3xD(128)(0);
  CNStageIntLLRInputS4xD(108)(2) <= VNStageIntLLROutputS3xD(128)(1);
  CNStageIntLLRInputS4xD(129)(2) <= VNStageIntLLROutputS3xD(128)(2);
  CNStageIntLLRInputS4xD(198)(2) <= VNStageIntLLROutputS3xD(128)(3);
  CNStageIntLLRInputS4xD(244)(2) <= VNStageIntLLROutputS3xD(128)(4);
  CNStageIntLLRInputS4xD(298)(2) <= VNStageIntLLROutputS3xD(128)(5);
  CNStageIntLLRInputS4xD(341)(2) <= VNStageIntLLROutputS3xD(128)(6);
  CNStageIntLLRInputS4xD(51)(2) <= VNStageIntLLROutputS3xD(129)(0);
  CNStageIntLLRInputS4xD(56)(2) <= VNStageIntLLROutputS3xD(129)(1);
  CNStageIntLLRInputS4xD(116)(2) <= VNStageIntLLROutputS3xD(129)(2);
  CNStageIntLLRInputS4xD(172)(2) <= VNStageIntLLROutputS3xD(129)(3);
  CNStageIntLLRInputS4xD(276)(2) <= VNStageIntLLROutputS3xD(129)(4);
  CNStageIntLLRInputS4xD(305)(2) <= VNStageIntLLROutputS3xD(129)(5);
  CNStageIntLLRInputS4xD(372)(2) <= VNStageIntLLROutputS3xD(129)(6);
  CNStageIntLLRInputS4xD(50)(2) <= VNStageIntLLROutputS3xD(130)(0);
  CNStageIntLLRInputS4xD(73)(2) <= VNStageIntLLROutputS3xD(130)(1);
  CNStageIntLLRInputS4xD(140)(2) <= VNStageIntLLROutputS3xD(130)(2);
  CNStageIntLLRInputS4xD(188)(2) <= VNStageIntLLROutputS3xD(130)(3);
  CNStageIntLLRInputS4xD(245)(2) <= VNStageIntLLROutputS3xD(130)(4);
  CNStageIntLLRInputS4xD(285)(2) <= VNStageIntLLROutputS3xD(130)(5);
  CNStageIntLLRInputS4xD(65)(2) <= VNStageIntLLROutputS3xD(131)(0);
  CNStageIntLLRInputS4xD(154)(2) <= VNStageIntLLROutputS3xD(131)(1);
  CNStageIntLLRInputS4xD(206)(2) <= VNStageIntLLROutputS3xD(131)(2);
  CNStageIntLLRInputS4xD(243)(2) <= VNStageIntLLROutputS3xD(131)(3);
  CNStageIntLLRInputS4xD(307)(2) <= VNStageIntLLROutputS3xD(131)(4);
  CNStageIntLLRInputS4xD(334)(2) <= VNStageIntLLROutputS3xD(131)(5);
  CNStageIntLLRInputS4xD(49)(2) <= VNStageIntLLROutputS3xD(132)(0);
  CNStageIntLLRInputS4xD(151)(2) <= VNStageIntLLROutputS3xD(132)(1);
  CNStageIntLLRInputS4xD(214)(2) <= VNStageIntLLROutputS3xD(132)(2);
  CNStageIntLLRInputS4xD(274)(2) <= VNStageIntLLROutputS3xD(132)(3);
  CNStageIntLLRInputS4xD(321)(2) <= VNStageIntLLROutputS3xD(132)(4);
  CNStageIntLLRInputS4xD(364)(2) <= VNStageIntLLROutputS3xD(132)(5);
  CNStageIntLLRInputS4xD(48)(2) <= VNStageIntLLROutputS3xD(133)(0);
  CNStageIntLLRInputS4xD(209)(2) <= VNStageIntLLROutputS3xD(133)(1);
  CNStageIntLLRInputS4xD(255)(2) <= VNStageIntLLROutputS3xD(133)(2);
  CNStageIntLLRInputS4xD(317)(2) <= VNStageIntLLROutputS3xD(133)(3);
  CNStageIntLLRInputS4xD(380)(2) <= VNStageIntLLROutputS3xD(133)(4);
  CNStageIntLLRInputS4xD(47)(2) <= VNStageIntLLROutputS3xD(134)(0);
  CNStageIntLLRInputS4xD(100)(2) <= VNStageIntLLROutputS3xD(134)(1);
  CNStageIntLLRInputS4xD(134)(2) <= VNStageIntLLROutputS3xD(134)(2);
  CNStageIntLLRInputS4xD(258)(2) <= VNStageIntLLROutputS3xD(134)(3);
  CNStageIntLLRInputS4xD(46)(2) <= VNStageIntLLROutputS3xD(135)(0);
  CNStageIntLLRInputS4xD(103)(2) <= VNStageIntLLROutputS3xD(135)(1);
  CNStageIntLLRInputS4xD(135)(2) <= VNStageIntLLROutputS3xD(135)(2);
  CNStageIntLLRInputS4xD(205)(2) <= VNStageIntLLROutputS3xD(135)(3);
  CNStageIntLLRInputS4xD(45)(2) <= VNStageIntLLROutputS3xD(136)(0);
  CNStageIntLLRInputS4xD(94)(2) <= VNStageIntLLROutputS3xD(136)(1);
  CNStageIntLLRInputS4xD(111)(2) <= VNStageIntLLROutputS3xD(136)(2);
  CNStageIntLLRInputS4xD(175)(2) <= VNStageIntLLROutputS3xD(136)(3);
  CNStageIntLLRInputS4xD(275)(2) <= VNStageIntLLROutputS3xD(136)(4);
  CNStageIntLLRInputS4xD(301)(2) <= VNStageIntLLROutputS3xD(136)(5);
  CNStageIntLLRInputS4xD(352)(2) <= VNStageIntLLROutputS3xD(136)(6);
  CNStageIntLLRInputS4xD(44)(2) <= VNStageIntLLROutputS3xD(137)(0);
  CNStageIntLLRInputS4xD(74)(2) <= VNStageIntLLROutputS3xD(137)(1);
  CNStageIntLLRInputS4xD(161)(2) <= VNStageIntLLROutputS3xD(137)(2);
  CNStageIntLLRInputS4xD(182)(2) <= VNStageIntLLROutputS3xD(137)(3);
  CNStageIntLLRInputS4xD(242)(2) <= VNStageIntLLROutputS3xD(137)(4);
  CNStageIntLLRInputS4xD(282)(2) <= VNStageIntLLROutputS3xD(137)(5);
  CNStageIntLLRInputS4xD(366)(2) <= VNStageIntLLROutputS3xD(137)(6);
  CNStageIntLLRInputS4xD(43)(2) <= VNStageIntLLROutputS3xD(138)(0);
  CNStageIntLLRInputS4xD(55)(2) <= VNStageIntLLROutputS3xD(138)(1);
  CNStageIntLLRInputS4xD(120)(2) <= VNStageIntLLROutputS3xD(138)(2);
  CNStageIntLLRInputS4xD(218)(2) <= VNStageIntLLROutputS3xD(138)(3);
  CNStageIntLLRInputS4xD(268)(2) <= VNStageIntLLROutputS3xD(138)(4);
  CNStageIntLLRInputS4xD(327)(2) <= VNStageIntLLROutputS3xD(138)(5);
  CNStageIntLLRInputS4xD(362)(2) <= VNStageIntLLROutputS3xD(138)(6);
  CNStageIntLLRInputS4xD(42)(2) <= VNStageIntLLROutputS3xD(139)(0);
  CNStageIntLLRInputS4xD(69)(2) <= VNStageIntLLROutputS3xD(139)(1);
  CNStageIntLLRInputS4xD(124)(2) <= VNStageIntLLROutputS3xD(139)(2);
  CNStageIntLLRInputS4xD(220)(2) <= VNStageIntLLROutputS3xD(139)(3);
  CNStageIntLLRInputS4xD(252)(2) <= VNStageIntLLROutputS3xD(139)(4);
  CNStageIntLLRInputS4xD(289)(2) <= VNStageIntLLROutputS3xD(139)(5);
  CNStageIntLLRInputS4xD(383)(2) <= VNStageIntLLROutputS3xD(139)(6);
  CNStageIntLLRInputS4xD(41)(2) <= VNStageIntLLROutputS3xD(140)(0);
  CNStageIntLLRInputS4xD(80)(2) <= VNStageIntLLROutputS3xD(140)(1);
  CNStageIntLLRInputS4xD(170)(2) <= VNStageIntLLROutputS3xD(140)(2);
  CNStageIntLLRInputS4xD(191)(2) <= VNStageIntLLROutputS3xD(140)(3);
  CNStageIntLLRInputS4xD(277)(2) <= VNStageIntLLROutputS3xD(140)(4);
  CNStageIntLLRInputS4xD(293)(2) <= VNStageIntLLROutputS3xD(140)(5);
  CNStageIntLLRInputS4xD(346)(2) <= VNStageIntLLROutputS3xD(140)(6);
  CNStageIntLLRInputS4xD(123)(2) <= VNStageIntLLROutputS3xD(141)(0);
  CNStageIntLLRInputS4xD(173)(2) <= VNStageIntLLROutputS3xD(141)(1);
  CNStageIntLLRInputS4xD(269)(2) <= VNStageIntLLROutputS3xD(141)(2);
  CNStageIntLLRInputS4xD(332)(2) <= VNStageIntLLROutputS3xD(141)(3);
  CNStageIntLLRInputS4xD(347)(2) <= VNStageIntLLROutputS3xD(141)(4);
  CNStageIntLLRInputS4xD(40)(2) <= VNStageIntLLROutputS3xD(142)(0);
  CNStageIntLLRInputS4xD(96)(2) <= VNStageIntLLROutputS3xD(142)(1);
  CNStageIntLLRInputS4xD(118)(2) <= VNStageIntLLROutputS3xD(142)(2);
  CNStageIntLLRInputS4xD(256)(2) <= VNStageIntLLROutputS3xD(142)(3);
  CNStageIntLLRInputS4xD(382)(2) <= VNStageIntLLROutputS3xD(142)(4);
  CNStageIntLLRInputS4xD(39)(2) <= VNStageIntLLROutputS3xD(143)(0);
  CNStageIntLLRInputS4xD(83)(2) <= VNStageIntLLROutputS3xD(143)(1);
  CNStageIntLLRInputS4xD(158)(2) <= VNStageIntLLROutputS3xD(143)(2);
  CNStageIntLLRInputS4xD(192)(2) <= VNStageIntLLROutputS3xD(143)(3);
  CNStageIntLLRInputS4xD(273)(2) <= VNStageIntLLROutputS3xD(143)(4);
  CNStageIntLLRInputS4xD(287)(2) <= VNStageIntLLROutputS3xD(143)(5);
  CNStageIntLLRInputS4xD(373)(2) <= VNStageIntLLROutputS3xD(143)(6);
  CNStageIntLLRInputS4xD(38)(2) <= VNStageIntLLROutputS3xD(144)(0);
  CNStageIntLLRInputS4xD(98)(2) <= VNStageIntLLROutputS3xD(144)(1);
  CNStageIntLLRInputS4xD(166)(2) <= VNStageIntLLROutputS3xD(144)(2);
  CNStageIntLLRInputS4xD(219)(2) <= VNStageIntLLROutputS3xD(144)(3);
  CNStageIntLLRInputS4xD(249)(2) <= VNStageIntLLROutputS3xD(144)(4);
  CNStageIntLLRInputS4xD(324)(2) <= VNStageIntLLROutputS3xD(144)(5);
  CNStageIntLLRInputS4xD(333)(2) <= VNStageIntLLROutputS3xD(144)(6);
  CNStageIntLLRInputS4xD(37)(2) <= VNStageIntLLROutputS3xD(145)(0);
  CNStageIntLLRInputS4xD(61)(2) <= VNStageIntLLROutputS3xD(145)(1);
  CNStageIntLLRInputS4xD(130)(2) <= VNStageIntLLROutputS3xD(145)(2);
  CNStageIntLLRInputS4xD(181)(2) <= VNStageIntLLROutputS3xD(145)(3);
  CNStageIntLLRInputS4xD(247)(2) <= VNStageIntLLROutputS3xD(145)(4);
  CNStageIntLLRInputS4xD(331)(2) <= VNStageIntLLROutputS3xD(145)(5);
  CNStageIntLLRInputS4xD(336)(2) <= VNStageIntLLROutputS3xD(145)(6);
  CNStageIntLLRInputS4xD(36)(2) <= VNStageIntLLROutputS3xD(146)(0);
  CNStageIntLLRInputS4xD(71)(2) <= VNStageIntLLROutputS3xD(146)(1);
  CNStageIntLLRInputS4xD(128)(2) <= VNStageIntLLROutputS3xD(146)(2);
  CNStageIntLLRInputS4xD(261)(2) <= VNStageIntLLROutputS3xD(146)(3);
  CNStageIntLLRInputS4xD(299)(2) <= VNStageIntLLROutputS3xD(146)(4);
  CNStageIntLLRInputS4xD(35)(2) <= VNStageIntLLROutputS3xD(147)(0);
  CNStageIntLLRInputS4xD(66)(2) <= VNStageIntLLROutputS3xD(147)(1);
  CNStageIntLLRInputS4xD(164)(2) <= VNStageIntLLROutputS3xD(147)(2);
  CNStageIntLLRInputS4xD(187)(2) <= VNStageIntLLROutputS3xD(147)(3);
  CNStageIntLLRInputS4xD(253)(2) <= VNStageIntLLROutputS3xD(147)(4);
  CNStageIntLLRInputS4xD(297)(2) <= VNStageIntLLROutputS3xD(147)(5);
  CNStageIntLLRInputS4xD(335)(2) <= VNStageIntLLROutputS3xD(147)(6);
  CNStageIntLLRInputS4xD(34)(2) <= VNStageIntLLROutputS3xD(148)(0);
  CNStageIntLLRInputS4xD(72)(2) <= VNStageIntLLROutputS3xD(148)(1);
  CNStageIntLLRInputS4xD(143)(2) <= VNStageIntLLROutputS3xD(148)(2);
  CNStageIntLLRInputS4xD(207)(2) <= VNStageIntLLROutputS3xD(148)(3);
  CNStageIntLLRInputS4xD(231)(2) <= VNStageIntLLROutputS3xD(148)(4);
  CNStageIntLLRInputS4xD(329)(2) <= VNStageIntLLROutputS3xD(148)(5);
  CNStageIntLLRInputS4xD(33)(2) <= VNStageIntLLROutputS3xD(149)(0);
  CNStageIntLLRInputS4xD(60)(2) <= VNStageIntLLROutputS3xD(149)(1);
  CNStageIntLLRInputS4xD(146)(2) <= VNStageIntLLROutputS3xD(149)(2);
  CNStageIntLLRInputS4xD(221)(2) <= VNStageIntLLROutputS3xD(149)(3);
  CNStageIntLLRInputS4xD(241)(2) <= VNStageIntLLROutputS3xD(149)(4);
  CNStageIntLLRInputS4xD(309)(2) <= VNStageIntLLROutputS3xD(149)(5);
  CNStageIntLLRInputS4xD(370)(2) <= VNStageIntLLROutputS3xD(149)(6);
  CNStageIntLLRInputS4xD(32)(2) <= VNStageIntLLROutputS3xD(150)(0);
  CNStageIntLLRInputS4xD(86)(2) <= VNStageIntLLROutputS3xD(150)(1);
  CNStageIntLLRInputS4xD(131)(2) <= VNStageIntLLROutputS3xD(150)(2);
  CNStageIntLLRInputS4xD(217)(2) <= VNStageIntLLROutputS3xD(150)(3);
  CNStageIntLLRInputS4xD(312)(2) <= VNStageIntLLROutputS3xD(150)(4);
  CNStageIntLLRInputS4xD(378)(2) <= VNStageIntLLROutputS3xD(150)(5);
  CNStageIntLLRInputS4xD(31)(2) <= VNStageIntLLROutputS3xD(151)(0);
  CNStageIntLLRInputS4xD(92)(2) <= VNStageIntLLROutputS3xD(151)(1);
  CNStageIntLLRInputS4xD(165)(2) <= VNStageIntLLROutputS3xD(151)(2);
  CNStageIntLLRInputS4xD(184)(2) <= VNStageIntLLROutputS3xD(151)(3);
  CNStageIntLLRInputS4xD(238)(2) <= VNStageIntLLROutputS3xD(151)(4);
  CNStageIntLLRInputS4xD(342)(2) <= VNStageIntLLROutputS3xD(151)(5);
  CNStageIntLLRInputS4xD(30)(2) <= VNStageIntLLROutputS3xD(152)(0);
  CNStageIntLLRInputS4xD(76)(2) <= VNStageIntLLROutputS3xD(152)(1);
  CNStageIntLLRInputS4xD(127)(2) <= VNStageIntLLROutputS3xD(152)(2);
  CNStageIntLLRInputS4xD(202)(2) <= VNStageIntLLROutputS3xD(152)(3);
  CNStageIntLLRInputS4xD(228)(2) <= VNStageIntLLROutputS3xD(152)(4);
  CNStageIntLLRInputS4xD(330)(2) <= VNStageIntLLROutputS3xD(152)(5);
  CNStageIntLLRInputS4xD(340)(2) <= VNStageIntLLROutputS3xD(152)(6);
  CNStageIntLLRInputS4xD(29)(2) <= VNStageIntLLROutputS3xD(153)(0);
  CNStageIntLLRInputS4xD(78)(2) <= VNStageIntLLROutputS3xD(153)(1);
  CNStageIntLLRInputS4xD(155)(2) <= VNStageIntLLROutputS3xD(153)(2);
  CNStageIntLLRInputS4xD(203)(2) <= VNStageIntLLROutputS3xD(153)(3);
  CNStageIntLLRInputS4xD(262)(2) <= VNStageIntLLROutputS3xD(153)(4);
  CNStageIntLLRInputS4xD(296)(2) <= VNStageIntLLROutputS3xD(153)(5);
  CNStageIntLLRInputS4xD(376)(2) <= VNStageIntLLROutputS3xD(153)(6);
  CNStageIntLLRInputS4xD(28)(2) <= VNStageIntLLROutputS3xD(154)(0);
  CNStageIntLLRInputS4xD(139)(2) <= VNStageIntLLROutputS3xD(154)(1);
  CNStageIntLLRInputS4xD(183)(2) <= VNStageIntLLROutputS3xD(154)(2);
  CNStageIntLLRInputS4xD(246)(2) <= VNStageIntLLROutputS3xD(154)(3);
  CNStageIntLLRInputS4xD(322)(2) <= VNStageIntLLROutputS3xD(154)(4);
  CNStageIntLLRInputS4xD(27)(2) <= VNStageIntLLROutputS3xD(155)(0);
  CNStageIntLLRInputS4xD(84)(2) <= VNStageIntLLROutputS3xD(155)(1);
  CNStageIntLLRInputS4xD(167)(2) <= VNStageIntLLROutputS3xD(155)(2);
  CNStageIntLLRInputS4xD(174)(2) <= VNStageIntLLROutputS3xD(155)(3);
  CNStageIntLLRInputS4xD(257)(2) <= VNStageIntLLROutputS3xD(155)(4);
  CNStageIntLLRInputS4xD(306)(2) <= VNStageIntLLROutputS3xD(155)(5);
  CNStageIntLLRInputS4xD(357)(2) <= VNStageIntLLROutputS3xD(155)(6);
  CNStageIntLLRInputS4xD(26)(2) <= VNStageIntLLROutputS3xD(156)(0);
  CNStageIntLLRInputS4xD(95)(2) <= VNStageIntLLROutputS3xD(156)(1);
  CNStageIntLLRInputS4xD(157)(2) <= VNStageIntLLROutputS3xD(156)(2);
  CNStageIntLLRInputS4xD(343)(2) <= VNStageIntLLROutputS3xD(156)(3);
  CNStageIntLLRInputS4xD(25)(2) <= VNStageIntLLROutputS3xD(157)(0);
  CNStageIntLLRInputS4xD(102)(2) <= VNStageIntLLROutputS3xD(157)(1);
  CNStageIntLLRInputS4xD(144)(2) <= VNStageIntLLROutputS3xD(157)(2);
  CNStageIntLLRInputS4xD(194)(2) <= VNStageIntLLROutputS3xD(157)(3);
  CNStageIntLLRInputS4xD(323)(2) <= VNStageIntLLROutputS3xD(157)(4);
  CNStageIntLLRInputS4xD(377)(2) <= VNStageIntLLROutputS3xD(157)(5);
  CNStageIntLLRInputS4xD(24)(2) <= VNStageIntLLROutputS3xD(158)(0);
  CNStageIntLLRInputS4xD(77)(2) <= VNStageIntLLROutputS3xD(158)(1);
  CNStageIntLLRInputS4xD(163)(2) <= VNStageIntLLROutputS3xD(158)(2);
  CNStageIntLLRInputS4xD(224)(2) <= VNStageIntLLROutputS3xD(158)(3);
  CNStageIntLLRInputS4xD(230)(2) <= VNStageIntLLROutputS3xD(158)(4);
  CNStageIntLLRInputS4xD(310)(2) <= VNStageIntLLROutputS3xD(158)(5);
  CNStageIntLLRInputS4xD(339)(2) <= VNStageIntLLROutputS3xD(158)(6);
  CNStageIntLLRInputS4xD(23)(2) <= VNStageIntLLROutputS3xD(159)(0);
  CNStageIntLLRInputS4xD(91)(2) <= VNStageIntLLROutputS3xD(159)(1);
  CNStageIntLLRInputS4xD(136)(2) <= VNStageIntLLROutputS3xD(159)(2);
  CNStageIntLLRInputS4xD(271)(2) <= VNStageIntLLROutputS3xD(159)(3);
  CNStageIntLLRInputS4xD(367)(2) <= VNStageIntLLROutputS3xD(159)(4);
  CNStageIntLLRInputS4xD(22)(2) <= VNStageIntLLROutputS3xD(160)(0);
  CNStageIntLLRInputS4xD(62)(2) <= VNStageIntLLROutputS3xD(160)(1);
  CNStageIntLLRInputS4xD(133)(2) <= VNStageIntLLROutputS3xD(160)(2);
  CNStageIntLLRInputS4xD(189)(2) <= VNStageIntLLROutputS3xD(160)(3);
  CNStageIntLLRInputS4xD(233)(2) <= VNStageIntLLROutputS3xD(160)(4);
  CNStageIntLLRInputS4xD(302)(2) <= VNStageIntLLROutputS3xD(160)(5);
  CNStageIntLLRInputS4xD(351)(2) <= VNStageIntLLROutputS3xD(160)(6);
  CNStageIntLLRInputS4xD(21)(2) <= VNStageIntLLROutputS3xD(161)(0);
  CNStageIntLLRInputS4xD(97)(2) <= VNStageIntLLROutputS3xD(161)(1);
  CNStageIntLLRInputS4xD(149)(2) <= VNStageIntLLROutputS3xD(161)(2);
  CNStageIntLLRInputS4xD(171)(2) <= VNStageIntLLROutputS3xD(161)(3);
  CNStageIntLLRInputS4xD(250)(2) <= VNStageIntLLROutputS3xD(161)(4);
  CNStageIntLLRInputS4xD(300)(2) <= VNStageIntLLROutputS3xD(161)(5);
  CNStageIntLLRInputS4xD(379)(2) <= VNStageIntLLROutputS3xD(161)(6);
  CNStageIntLLRInputS4xD(20)(2) <= VNStageIntLLROutputS3xD(162)(0);
  CNStageIntLLRInputS4xD(64)(2) <= VNStageIntLLROutputS3xD(162)(1);
  CNStageIntLLRInputS4xD(141)(2) <= VNStageIntLLROutputS3xD(162)(2);
  CNStageIntLLRInputS4xD(179)(2) <= VNStageIntLLROutputS3xD(162)(3);
  CNStageIntLLRInputS4xD(259)(2) <= VNStageIntLLROutputS3xD(162)(4);
  CNStageIntLLRInputS4xD(315)(2) <= VNStageIntLLROutputS3xD(162)(5);
  CNStageIntLLRInputS4xD(369)(2) <= VNStageIntLLROutputS3xD(162)(6);
  CNStageIntLLRInputS4xD(19)(2) <= VNStageIntLLROutputS3xD(163)(0);
  CNStageIntLLRInputS4xD(79)(2) <= VNStageIntLLROutputS3xD(163)(1);
  CNStageIntLLRInputS4xD(115)(2) <= VNStageIntLLROutputS3xD(163)(2);
  CNStageIntLLRInputS4xD(254)(2) <= VNStageIntLLROutputS3xD(163)(3);
  CNStageIntLLRInputS4xD(355)(2) <= VNStageIntLLROutputS3xD(163)(4);
  CNStageIntLLRInputS4xD(18)(2) <= VNStageIntLLROutputS3xD(164)(0);
  CNStageIntLLRInputS4xD(75)(2) <= VNStageIntLLROutputS3xD(164)(1);
  CNStageIntLLRInputS4xD(125)(2) <= VNStageIntLLROutputS3xD(164)(2);
  CNStageIntLLRInputS4xD(197)(2) <= VNStageIntLLROutputS3xD(164)(3);
  CNStageIntLLRInputS4xD(260)(2) <= VNStageIntLLROutputS3xD(164)(4);
  CNStageIntLLRInputS4xD(375)(2) <= VNStageIntLLROutputS3xD(164)(5);
  CNStageIntLLRInputS4xD(17)(2) <= VNStageIntLLROutputS3xD(165)(0);
  CNStageIntLLRInputS4xD(93)(2) <= VNStageIntLLROutputS3xD(165)(1);
  CNStageIntLLRInputS4xD(119)(2) <= VNStageIntLLROutputS3xD(165)(2);
  CNStageIntLLRInputS4xD(177)(2) <= VNStageIntLLROutputS3xD(165)(3);
  CNStageIntLLRInputS4xD(294)(2) <= VNStageIntLLROutputS3xD(165)(4);
  CNStageIntLLRInputS4xD(348)(2) <= VNStageIntLLROutputS3xD(165)(5);
  CNStageIntLLRInputS4xD(16)(2) <= VNStageIntLLROutputS3xD(166)(0);
  CNStageIntLLRInputS4xD(57)(2) <= VNStageIntLLROutputS3xD(166)(1);
  CNStageIntLLRInputS4xD(122)(2) <= VNStageIntLLROutputS3xD(166)(2);
  CNStageIntLLRInputS4xD(210)(2) <= VNStageIntLLROutputS3xD(166)(3);
  CNStageIntLLRInputS4xD(288)(2) <= VNStageIntLLROutputS3xD(166)(4);
  CNStageIntLLRInputS4xD(345)(2) <= VNStageIntLLROutputS3xD(166)(5);
  CNStageIntLLRInputS4xD(15)(2) <= VNStageIntLLROutputS3xD(167)(0);
  CNStageIntLLRInputS4xD(58)(2) <= VNStageIntLLROutputS3xD(167)(1);
  CNStageIntLLRInputS4xD(112)(2) <= VNStageIntLLROutputS3xD(167)(2);
  CNStageIntLLRInputS4xD(213)(2) <= VNStageIntLLROutputS3xD(167)(3);
  CNStageIntLLRInputS4xD(225)(2) <= VNStageIntLLROutputS3xD(167)(4);
  CNStageIntLLRInputS4xD(292)(2) <= VNStageIntLLROutputS3xD(167)(5);
  CNStageIntLLRInputS4xD(360)(2) <= VNStageIntLLROutputS3xD(167)(6);
  CNStageIntLLRInputS4xD(14)(2) <= VNStageIntLLROutputS3xD(168)(0);
  CNStageIntLLRInputS4xD(150)(2) <= VNStageIntLLROutputS3xD(168)(1);
  CNStageIntLLRInputS4xD(199)(2) <= VNStageIntLLROutputS3xD(168)(2);
  CNStageIntLLRInputS4xD(264)(2) <= VNStageIntLLROutputS3xD(168)(3);
  CNStageIntLLRInputS4xD(283)(2) <= VNStageIntLLROutputS3xD(168)(4);
  CNStageIntLLRInputS4xD(353)(2) <= VNStageIntLLROutputS3xD(168)(5);
  CNStageIntLLRInputS4xD(13)(2) <= VNStageIntLLROutputS3xD(169)(0);
  CNStageIntLLRInputS4xD(85)(2) <= VNStageIntLLROutputS3xD(169)(1);
  CNStageIntLLRInputS4xD(132)(2) <= VNStageIntLLROutputS3xD(169)(2);
  CNStageIntLLRInputS4xD(178)(2) <= VNStageIntLLROutputS3xD(169)(3);
  CNStageIntLLRInputS4xD(266)(2) <= VNStageIntLLROutputS3xD(169)(4);
  CNStageIntLLRInputS4xD(316)(2) <= VNStageIntLLROutputS3xD(169)(5);
  CNStageIntLLRInputS4xD(12)(2) <= VNStageIntLLROutputS3xD(170)(0);
  CNStageIntLLRInputS4xD(101)(2) <= VNStageIntLLROutputS3xD(170)(1);
  CNStageIntLLRInputS4xD(145)(2) <= VNStageIntLLROutputS3xD(170)(2);
  CNStageIntLLRInputS4xD(236)(2) <= VNStageIntLLROutputS3xD(170)(3);
  CNStageIntLLRInputS4xD(337)(2) <= VNStageIntLLROutputS3xD(170)(4);
  CNStageIntLLRInputS4xD(105)(2) <= VNStageIntLLROutputS3xD(171)(0);
  CNStageIntLLRInputS4xD(156)(2) <= VNStageIntLLROutputS3xD(171)(1);
  CNStageIntLLRInputS4xD(222)(2) <= VNStageIntLLROutputS3xD(171)(2);
  CNStageIntLLRInputS4xD(311)(2) <= VNStageIntLLROutputS3xD(171)(3);
  CNStageIntLLRInputS4xD(11)(2) <= VNStageIntLLROutputS3xD(172)(0);
  CNStageIntLLRInputS4xD(110)(2) <= VNStageIntLLROutputS3xD(172)(1);
  CNStageIntLLRInputS4xD(126)(2) <= VNStageIntLLROutputS3xD(172)(2);
  CNStageIntLLRInputS4xD(229)(2) <= VNStageIntLLROutputS3xD(172)(3);
  CNStageIntLLRInputS4xD(10)(2) <= VNStageIntLLROutputS3xD(173)(0);
  CNStageIntLLRInputS4xD(104)(2) <= VNStageIntLLROutputS3xD(173)(1);
  CNStageIntLLRInputS4xD(114)(2) <= VNStageIntLLROutputS3xD(173)(2);
  CNStageIntLLRInputS4xD(180)(2) <= VNStageIntLLROutputS3xD(173)(3);
  CNStageIntLLRInputS4xD(237)(2) <= VNStageIntLLROutputS3xD(173)(4);
  CNStageIntLLRInputS4xD(295)(2) <= VNStageIntLLROutputS3xD(173)(5);
  CNStageIntLLRInputS4xD(9)(2) <= VNStageIntLLROutputS3xD(174)(0);
  CNStageIntLLRInputS4xD(99)(2) <= VNStageIntLLROutputS3xD(174)(1);
  CNStageIntLLRInputS4xD(159)(2) <= VNStageIntLLROutputS3xD(174)(2);
  CNStageIntLLRInputS4xD(265)(2) <= VNStageIntLLROutputS3xD(174)(3);
  CNStageIntLLRInputS4xD(361)(2) <= VNStageIntLLROutputS3xD(174)(4);
  CNStageIntLLRInputS4xD(8)(2) <= VNStageIntLLROutputS3xD(175)(0);
  CNStageIntLLRInputS4xD(82)(2) <= VNStageIntLLROutputS3xD(175)(1);
  CNStageIntLLRInputS4xD(117)(2) <= VNStageIntLLROutputS3xD(175)(2);
  CNStageIntLLRInputS4xD(211)(2) <= VNStageIntLLROutputS3xD(175)(3);
  CNStageIntLLRInputS4xD(278)(2) <= VNStageIntLLROutputS3xD(175)(4);
  CNStageIntLLRInputS4xD(325)(2) <= VNStageIntLLROutputS3xD(175)(5);
  CNStageIntLLRInputS4xD(344)(2) <= VNStageIntLLROutputS3xD(175)(6);
  CNStageIntLLRInputS4xD(7)(2) <= VNStageIntLLROutputS3xD(176)(0);
  CNStageIntLLRInputS4xD(89)(2) <= VNStageIntLLROutputS3xD(176)(1);
  CNStageIntLLRInputS4xD(137)(2) <= VNStageIntLLROutputS3xD(176)(2);
  CNStageIntLLRInputS4xD(176)(2) <= VNStageIntLLROutputS3xD(176)(3);
  CNStageIntLLRInputS4xD(251)(2) <= VNStageIntLLROutputS3xD(176)(4);
  CNStageIntLLRInputS4xD(286)(2) <= VNStageIntLLROutputS3xD(176)(5);
  CNStageIntLLRInputS4xD(356)(2) <= VNStageIntLLROutputS3xD(176)(6);
  CNStageIntLLRInputS4xD(6)(2) <= VNStageIntLLROutputS3xD(177)(0);
  CNStageIntLLRInputS4xD(109)(2) <= VNStageIntLLROutputS3xD(177)(1);
  CNStageIntLLRInputS4xD(147)(2) <= VNStageIntLLROutputS3xD(177)(2);
  CNStageIntLLRInputS4xD(204)(2) <= VNStageIntLLROutputS3xD(177)(3);
  CNStageIntLLRInputS4xD(232)(2) <= VNStageIntLLROutputS3xD(177)(4);
  CNStageIntLLRInputS4xD(304)(2) <= VNStageIntLLROutputS3xD(177)(5);
  CNStageIntLLRInputS4xD(368)(2) <= VNStageIntLLROutputS3xD(177)(6);
  CNStageIntLLRInputS4xD(5)(2) <= VNStageIntLLROutputS3xD(178)(0);
  CNStageIntLLRInputS4xD(107)(2) <= VNStageIntLLROutputS3xD(178)(1);
  CNStageIntLLRInputS4xD(142)(2) <= VNStageIntLLROutputS3xD(178)(2);
  CNStageIntLLRInputS4xD(201)(2) <= VNStageIntLLROutputS3xD(178)(3);
  CNStageIntLLRInputS4xD(313)(2) <= VNStageIntLLROutputS3xD(178)(4);
  CNStageIntLLRInputS4xD(338)(2) <= VNStageIntLLROutputS3xD(178)(5);
  CNStageIntLLRInputS4xD(4)(2) <= VNStageIntLLROutputS3xD(179)(0);
  CNStageIntLLRInputS4xD(87)(2) <= VNStageIntLLROutputS3xD(179)(1);
  CNStageIntLLRInputS4xD(148)(2) <= VNStageIntLLROutputS3xD(179)(2);
  CNStageIntLLRInputS4xD(215)(2) <= VNStageIntLLROutputS3xD(179)(3);
  CNStageIntLLRInputS4xD(267)(2) <= VNStageIntLLROutputS3xD(179)(4);
  CNStageIntLLRInputS4xD(308)(2) <= VNStageIntLLROutputS3xD(179)(5);
  CNStageIntLLRInputS4xD(67)(2) <= VNStageIntLLROutputS3xD(180)(0);
  CNStageIntLLRInputS4xD(208)(2) <= VNStageIntLLROutputS3xD(180)(1);
  CNStageIntLLRInputS4xD(263)(2) <= VNStageIntLLROutputS3xD(180)(2);
  CNStageIntLLRInputS4xD(314)(2) <= VNStageIntLLROutputS3xD(180)(3);
  CNStageIntLLRInputS4xD(371)(2) <= VNStageIntLLROutputS3xD(180)(4);
  CNStageIntLLRInputS4xD(3)(2) <= VNStageIntLLROutputS3xD(181)(0);
  CNStageIntLLRInputS4xD(70)(2) <= VNStageIntLLROutputS3xD(181)(1);
  CNStageIntLLRInputS4xD(162)(2) <= VNStageIntLLROutputS3xD(181)(2);
  CNStageIntLLRInputS4xD(186)(2) <= VNStageIntLLROutputS3xD(181)(3);
  CNStageIntLLRInputS4xD(227)(2) <= VNStageIntLLROutputS3xD(181)(4);
  CNStageIntLLRInputS4xD(303)(2) <= VNStageIntLLROutputS3xD(181)(5);
  CNStageIntLLRInputS4xD(2)(2) <= VNStageIntLLROutputS3xD(182)(0);
  CNStageIntLLRInputS4xD(54)(2) <= VNStageIntLLROutputS3xD(182)(1);
  CNStageIntLLRInputS4xD(169)(2) <= VNStageIntLLROutputS3xD(182)(2);
  CNStageIntLLRInputS4xD(195)(2) <= VNStageIntLLROutputS3xD(182)(3);
  CNStageIntLLRInputS4xD(248)(2) <= VNStageIntLLROutputS3xD(182)(4);
  CNStageIntLLRInputS4xD(328)(2) <= VNStageIntLLROutputS3xD(182)(5);
  CNStageIntLLRInputS4xD(350)(2) <= VNStageIntLLROutputS3xD(182)(6);
  CNStageIntLLRInputS4xD(1)(2) <= VNStageIntLLROutputS3xD(183)(0);
  CNStageIntLLRInputS4xD(88)(2) <= VNStageIntLLROutputS3xD(183)(1);
  CNStageIntLLRInputS4xD(190)(2) <= VNStageIntLLROutputS3xD(183)(2);
  CNStageIntLLRInputS4xD(281)(2) <= VNStageIntLLROutputS3xD(183)(3);
  CNStageIntLLRInputS4xD(358)(2) <= VNStageIntLLROutputS3xD(183)(4);
  CNStageIntLLRInputS4xD(0)(2) <= VNStageIntLLROutputS3xD(184)(0);
  CNStageIntLLRInputS4xD(106)(2) <= VNStageIntLLROutputS3xD(184)(1);
  CNStageIntLLRInputS4xD(153)(2) <= VNStageIntLLROutputS3xD(184)(2);
  CNStageIntLLRInputS4xD(193)(2) <= VNStageIntLLROutputS3xD(184)(3);
  CNStageIntLLRInputS4xD(226)(2) <= VNStageIntLLROutputS3xD(184)(4);
  CNStageIntLLRInputS4xD(318)(2) <= VNStageIntLLROutputS3xD(184)(5);
  CNStageIntLLRInputS4xD(354)(2) <= VNStageIntLLROutputS3xD(184)(6);
  CNStageIntLLRInputS4xD(121)(2) <= VNStageIntLLROutputS3xD(185)(0);
  CNStageIntLLRInputS4xD(272)(2) <= VNStageIntLLROutputS3xD(185)(1);
  CNStageIntLLRInputS4xD(320)(2) <= VNStageIntLLROutputS3xD(185)(2);
  CNStageIntLLRInputS4xD(359)(2) <= VNStageIntLLROutputS3xD(185)(3);
  CNStageIntLLRInputS4xD(63)(2) <= VNStageIntLLROutputS3xD(186)(0);
  CNStageIntLLRInputS4xD(160)(2) <= VNStageIntLLROutputS3xD(186)(1);
  CNStageIntLLRInputS4xD(216)(2) <= VNStageIntLLROutputS3xD(186)(2);
  CNStageIntLLRInputS4xD(235)(2) <= VNStageIntLLROutputS3xD(186)(3);
  CNStageIntLLRInputS4xD(290)(2) <= VNStageIntLLROutputS3xD(186)(4);
  CNStageIntLLRInputS4xD(349)(2) <= VNStageIntLLROutputS3xD(186)(5);
  CNStageIntLLRInputS4xD(90)(2) <= VNStageIntLLROutputS3xD(187)(0);
  CNStageIntLLRInputS4xD(113)(2) <= VNStageIntLLROutputS3xD(187)(1);
  CNStageIntLLRInputS4xD(200)(2) <= VNStageIntLLROutputS3xD(187)(2);
  CNStageIntLLRInputS4xD(240)(2) <= VNStageIntLLROutputS3xD(187)(3);
  CNStageIntLLRInputS4xD(326)(2) <= VNStageIntLLROutputS3xD(187)(4);
  CNStageIntLLRInputS4xD(374)(2) <= VNStageIntLLROutputS3xD(187)(5);
  CNStageIntLLRInputS4xD(81)(2) <= VNStageIntLLROutputS3xD(188)(0);
  CNStageIntLLRInputS4xD(212)(2) <= VNStageIntLLROutputS3xD(188)(1);
  CNStageIntLLRInputS4xD(279)(2) <= VNStageIntLLROutputS3xD(188)(2);
  CNStageIntLLRInputS4xD(284)(2) <= VNStageIntLLROutputS3xD(188)(3);
  CNStageIntLLRInputS4xD(381)(2) <= VNStageIntLLROutputS3xD(188)(4);
  CNStageIntLLRInputS4xD(68)(2) <= VNStageIntLLROutputS3xD(189)(0);
  CNStageIntLLRInputS4xD(152)(2) <= VNStageIntLLROutputS3xD(189)(1);
  CNStageIntLLRInputS4xD(223)(2) <= VNStageIntLLROutputS3xD(189)(2);
  CNStageIntLLRInputS4xD(239)(2) <= VNStageIntLLROutputS3xD(189)(3);
  CNStageIntLLRInputS4xD(291)(2) <= VNStageIntLLROutputS3xD(189)(4);
  CNStageIntLLRInputS4xD(363)(2) <= VNStageIntLLROutputS3xD(189)(5);
  CNStageIntLLRInputS4xD(168)(2) <= VNStageIntLLROutputS3xD(190)(0);
  CNStageIntLLRInputS4xD(196)(2) <= VNStageIntLLROutputS3xD(190)(1);
  CNStageIntLLRInputS4xD(234)(2) <= VNStageIntLLROutputS3xD(190)(2);
  CNStageIntLLRInputS4xD(319)(2) <= VNStageIntLLROutputS3xD(190)(3);
  CNStageIntLLRInputS4xD(365)(2) <= VNStageIntLLROutputS3xD(190)(4);
  CNStageIntLLRInputS4xD(52)(2) <= VNStageIntLLROutputS3xD(191)(0);
  CNStageIntLLRInputS4xD(59)(2) <= VNStageIntLLROutputS3xD(191)(1);
  CNStageIntLLRInputS4xD(138)(2) <= VNStageIntLLROutputS3xD(191)(2);
  CNStageIntLLRInputS4xD(185)(2) <= VNStageIntLLROutputS3xD(191)(3);
  CNStageIntLLRInputS4xD(270)(2) <= VNStageIntLLROutputS3xD(191)(4);
  CNStageIntLLRInputS4xD(280)(2) <= VNStageIntLLROutputS3xD(191)(5);
  CNStageIntLLRInputS4xD(53)(3) <= VNStageIntLLROutputS3xD(192)(0);
  CNStageIntLLRInputS4xD(107)(3) <= VNStageIntLLROutputS3xD(192)(1);
  CNStageIntLLRInputS4xD(128)(3) <= VNStageIntLLROutputS3xD(192)(2);
  CNStageIntLLRInputS4xD(197)(3) <= VNStageIntLLROutputS3xD(192)(3);
  CNStageIntLLRInputS4xD(243)(3) <= VNStageIntLLROutputS3xD(192)(4);
  CNStageIntLLRInputS4xD(297)(3) <= VNStageIntLLROutputS3xD(192)(5);
  CNStageIntLLRInputS4xD(340)(3) <= VNStageIntLLROutputS3xD(192)(6);
  CNStageIntLLRInputS4xD(51)(3) <= VNStageIntLLROutputS3xD(193)(0);
  CNStageIntLLRInputS4xD(58)(3) <= VNStageIntLLROutputS3xD(193)(1);
  CNStageIntLLRInputS4xD(137)(3) <= VNStageIntLLROutputS3xD(193)(2);
  CNStageIntLLRInputS4xD(269)(3) <= VNStageIntLLROutputS3xD(193)(3);
  CNStageIntLLRInputS4xD(333)(3) <= VNStageIntLLROutputS3xD(193)(4);
  CNStageIntLLRInputS4xD(50)(3) <= VNStageIntLLROutputS3xD(194)(0);
  CNStageIntLLRInputS4xD(55)(3) <= VNStageIntLLROutputS3xD(194)(1);
  CNStageIntLLRInputS4xD(115)(3) <= VNStageIntLLROutputS3xD(194)(2);
  CNStageIntLLRInputS4xD(171)(3) <= VNStageIntLLROutputS3xD(194)(3);
  CNStageIntLLRInputS4xD(275)(3) <= VNStageIntLLROutputS3xD(194)(4);
  CNStageIntLLRInputS4xD(304)(3) <= VNStageIntLLROutputS3xD(194)(5);
  CNStageIntLLRInputS4xD(371)(3) <= VNStageIntLLROutputS3xD(194)(6);
  CNStageIntLLRInputS4xD(72)(3) <= VNStageIntLLROutputS3xD(195)(0);
  CNStageIntLLRInputS4xD(139)(3) <= VNStageIntLLROutputS3xD(195)(1);
  CNStageIntLLRInputS4xD(187)(3) <= VNStageIntLLROutputS3xD(195)(2);
  CNStageIntLLRInputS4xD(244)(3) <= VNStageIntLLROutputS3xD(195)(3);
  CNStageIntLLRInputS4xD(49)(3) <= VNStageIntLLROutputS3xD(196)(0);
  CNStageIntLLRInputS4xD(64)(3) <= VNStageIntLLROutputS3xD(196)(1);
  CNStageIntLLRInputS4xD(153)(3) <= VNStageIntLLROutputS3xD(196)(2);
  CNStageIntLLRInputS4xD(205)(3) <= VNStageIntLLROutputS3xD(196)(3);
  CNStageIntLLRInputS4xD(242)(3) <= VNStageIntLLROutputS3xD(196)(4);
  CNStageIntLLRInputS4xD(306)(3) <= VNStageIntLLROutputS3xD(196)(5);
  CNStageIntLLRInputS4xD(48)(3) <= VNStageIntLLROutputS3xD(197)(0);
  CNStageIntLLRInputS4xD(96)(3) <= VNStageIntLLROutputS3xD(197)(1);
  CNStageIntLLRInputS4xD(150)(3) <= VNStageIntLLROutputS3xD(197)(2);
  CNStageIntLLRInputS4xD(213)(3) <= VNStageIntLLROutputS3xD(197)(3);
  CNStageIntLLRInputS4xD(273)(3) <= VNStageIntLLROutputS3xD(197)(4);
  CNStageIntLLRInputS4xD(320)(3) <= VNStageIntLLROutputS3xD(197)(5);
  CNStageIntLLRInputS4xD(363)(3) <= VNStageIntLLROutputS3xD(197)(6);
  CNStageIntLLRInputS4xD(47)(3) <= VNStageIntLLROutputS3xD(198)(0);
  CNStageIntLLRInputS4xD(105)(3) <= VNStageIntLLROutputS3xD(198)(1);
  CNStageIntLLRInputS4xD(111)(3) <= VNStageIntLLROutputS3xD(198)(2);
  CNStageIntLLRInputS4xD(208)(3) <= VNStageIntLLROutputS3xD(198)(3);
  CNStageIntLLRInputS4xD(254)(3) <= VNStageIntLLROutputS3xD(198)(4);
  CNStageIntLLRInputS4xD(316)(3) <= VNStageIntLLROutputS3xD(198)(5);
  CNStageIntLLRInputS4xD(379)(3) <= VNStageIntLLROutputS3xD(198)(6);
  CNStageIntLLRInputS4xD(46)(3) <= VNStageIntLLROutputS3xD(199)(0);
  CNStageIntLLRInputS4xD(99)(3) <= VNStageIntLLROutputS3xD(199)(1);
  CNStageIntLLRInputS4xD(133)(3) <= VNStageIntLLROutputS3xD(199)(2);
  CNStageIntLLRInputS4xD(214)(3) <= VNStageIntLLROutputS3xD(199)(3);
  CNStageIntLLRInputS4xD(257)(3) <= VNStageIntLLROutputS3xD(199)(4);
  CNStageIntLLRInputS4xD(282)(3) <= VNStageIntLLROutputS3xD(199)(5);
  CNStageIntLLRInputS4xD(350)(3) <= VNStageIntLLROutputS3xD(199)(6);
  CNStageIntLLRInputS4xD(45)(3) <= VNStageIntLLROutputS3xD(200)(0);
  CNStageIntLLRInputS4xD(102)(3) <= VNStageIntLLROutputS3xD(200)(1);
  CNStageIntLLRInputS4xD(134)(3) <= VNStageIntLLROutputS3xD(200)(2);
  CNStageIntLLRInputS4xD(204)(3) <= VNStageIntLLROutputS3xD(200)(3);
  CNStageIntLLRInputS4xD(245)(3) <= VNStageIntLLROutputS3xD(200)(4);
  CNStageIntLLRInputS4xD(300)(3) <= VNStageIntLLROutputS3xD(200)(5);
  CNStageIntLLRInputS4xD(44)(3) <= VNStageIntLLROutputS3xD(201)(0);
  CNStageIntLLRInputS4xD(93)(3) <= VNStageIntLLROutputS3xD(201)(1);
  CNStageIntLLRInputS4xD(169)(3) <= VNStageIntLLROutputS3xD(201)(2);
  CNStageIntLLRInputS4xD(174)(3) <= VNStageIntLLROutputS3xD(201)(3);
  CNStageIntLLRInputS4xD(274)(3) <= VNStageIntLLROutputS3xD(201)(4);
  CNStageIntLLRInputS4xD(351)(3) <= VNStageIntLLROutputS3xD(201)(5);
  CNStageIntLLRInputS4xD(43)(3) <= VNStageIntLLROutputS3xD(202)(0);
  CNStageIntLLRInputS4xD(73)(3) <= VNStageIntLLROutputS3xD(202)(1);
  CNStageIntLLRInputS4xD(160)(3) <= VNStageIntLLROutputS3xD(202)(2);
  CNStageIntLLRInputS4xD(181)(3) <= VNStageIntLLROutputS3xD(202)(3);
  CNStageIntLLRInputS4xD(281)(3) <= VNStageIntLLROutputS3xD(202)(4);
  CNStageIntLLRInputS4xD(365)(3) <= VNStageIntLLROutputS3xD(202)(5);
  CNStageIntLLRInputS4xD(42)(3) <= VNStageIntLLROutputS3xD(203)(0);
  CNStageIntLLRInputS4xD(54)(3) <= VNStageIntLLROutputS3xD(203)(1);
  CNStageIntLLRInputS4xD(119)(3) <= VNStageIntLLROutputS3xD(203)(2);
  CNStageIntLLRInputS4xD(217)(3) <= VNStageIntLLROutputS3xD(203)(3);
  CNStageIntLLRInputS4xD(267)(3) <= VNStageIntLLROutputS3xD(203)(4);
  CNStageIntLLRInputS4xD(326)(3) <= VNStageIntLLROutputS3xD(203)(5);
  CNStageIntLLRInputS4xD(361)(3) <= VNStageIntLLROutputS3xD(203)(6);
  CNStageIntLLRInputS4xD(41)(3) <= VNStageIntLLROutputS3xD(204)(0);
  CNStageIntLLRInputS4xD(68)(3) <= VNStageIntLLROutputS3xD(204)(1);
  CNStageIntLLRInputS4xD(123)(3) <= VNStageIntLLROutputS3xD(204)(2);
  CNStageIntLLRInputS4xD(219)(3) <= VNStageIntLLROutputS3xD(204)(3);
  CNStageIntLLRInputS4xD(251)(3) <= VNStageIntLLROutputS3xD(204)(4);
  CNStageIntLLRInputS4xD(288)(3) <= VNStageIntLLROutputS3xD(204)(5);
  CNStageIntLLRInputS4xD(382)(3) <= VNStageIntLLROutputS3xD(204)(6);
  CNStageIntLLRInputS4xD(170)(3) <= VNStageIntLLROutputS3xD(205)(0);
  CNStageIntLLRInputS4xD(276)(3) <= VNStageIntLLROutputS3xD(205)(1);
  CNStageIntLLRInputS4xD(345)(3) <= VNStageIntLLROutputS3xD(205)(2);
  CNStageIntLLRInputS4xD(40)(3) <= VNStageIntLLROutputS3xD(206)(0);
  CNStageIntLLRInputS4xD(122)(3) <= VNStageIntLLROutputS3xD(206)(1);
  CNStageIntLLRInputS4xD(172)(3) <= VNStageIntLLROutputS3xD(206)(2);
  CNStageIntLLRInputS4xD(332)(3) <= VNStageIntLLROutputS3xD(206)(3);
  CNStageIntLLRInputS4xD(346)(3) <= VNStageIntLLROutputS3xD(206)(4);
  CNStageIntLLRInputS4xD(39)(3) <= VNStageIntLLROutputS3xD(207)(0);
  CNStageIntLLRInputS4xD(95)(3) <= VNStageIntLLROutputS3xD(207)(1);
  CNStageIntLLRInputS4xD(117)(3) <= VNStageIntLLROutputS3xD(207)(2);
  CNStageIntLLRInputS4xD(255)(3) <= VNStageIntLLROutputS3xD(207)(3);
  CNStageIntLLRInputS4xD(292)(3) <= VNStageIntLLROutputS3xD(207)(4);
  CNStageIntLLRInputS4xD(381)(3) <= VNStageIntLLROutputS3xD(207)(5);
  CNStageIntLLRInputS4xD(38)(3) <= VNStageIntLLROutputS3xD(208)(0);
  CNStageIntLLRInputS4xD(82)(3) <= VNStageIntLLROutputS3xD(208)(1);
  CNStageIntLLRInputS4xD(157)(3) <= VNStageIntLLROutputS3xD(208)(2);
  CNStageIntLLRInputS4xD(191)(3) <= VNStageIntLLROutputS3xD(208)(3);
  CNStageIntLLRInputS4xD(286)(3) <= VNStageIntLLROutputS3xD(208)(4);
  CNStageIntLLRInputS4xD(372)(3) <= VNStageIntLLROutputS3xD(208)(5);
  CNStageIntLLRInputS4xD(37)(3) <= VNStageIntLLROutputS3xD(209)(0);
  CNStageIntLLRInputS4xD(97)(3) <= VNStageIntLLROutputS3xD(209)(1);
  CNStageIntLLRInputS4xD(165)(3) <= VNStageIntLLROutputS3xD(209)(2);
  CNStageIntLLRInputS4xD(218)(3) <= VNStageIntLLROutputS3xD(209)(3);
  CNStageIntLLRInputS4xD(323)(3) <= VNStageIntLLROutputS3xD(209)(4);
  CNStageIntLLRInputS4xD(36)(3) <= VNStageIntLLROutputS3xD(210)(0);
  CNStageIntLLRInputS4xD(60)(3) <= VNStageIntLLROutputS3xD(210)(1);
  CNStageIntLLRInputS4xD(129)(3) <= VNStageIntLLROutputS3xD(210)(2);
  CNStageIntLLRInputS4xD(180)(3) <= VNStageIntLLROutputS3xD(210)(3);
  CNStageIntLLRInputS4xD(246)(3) <= VNStageIntLLROutputS3xD(210)(4);
  CNStageIntLLRInputS4xD(330)(3) <= VNStageIntLLROutputS3xD(210)(5);
  CNStageIntLLRInputS4xD(335)(3) <= VNStageIntLLROutputS3xD(210)(6);
  CNStageIntLLRInputS4xD(35)(3) <= VNStageIntLLROutputS3xD(211)(0);
  CNStageIntLLRInputS4xD(70)(3) <= VNStageIntLLROutputS3xD(211)(1);
  CNStageIntLLRInputS4xD(127)(3) <= VNStageIntLLROutputS3xD(211)(2);
  CNStageIntLLRInputS4xD(206)(3) <= VNStageIntLLROutputS3xD(211)(3);
  CNStageIntLLRInputS4xD(260)(3) <= VNStageIntLLROutputS3xD(211)(4);
  CNStageIntLLRInputS4xD(298)(3) <= VNStageIntLLROutputS3xD(211)(5);
  CNStageIntLLRInputS4xD(34)(3) <= VNStageIntLLROutputS3xD(212)(0);
  CNStageIntLLRInputS4xD(65)(3) <= VNStageIntLLROutputS3xD(212)(1);
  CNStageIntLLRInputS4xD(163)(3) <= VNStageIntLLROutputS3xD(212)(2);
  CNStageIntLLRInputS4xD(186)(3) <= VNStageIntLLROutputS3xD(212)(3);
  CNStageIntLLRInputS4xD(296)(3) <= VNStageIntLLROutputS3xD(212)(4);
  CNStageIntLLRInputS4xD(33)(3) <= VNStageIntLLROutputS3xD(213)(0);
  CNStageIntLLRInputS4xD(71)(3) <= VNStageIntLLROutputS3xD(213)(1);
  CNStageIntLLRInputS4xD(142)(3) <= VNStageIntLLROutputS3xD(213)(2);
  CNStageIntLLRInputS4xD(230)(3) <= VNStageIntLLROutputS3xD(213)(3);
  CNStageIntLLRInputS4xD(32)(3) <= VNStageIntLLROutputS3xD(214)(0);
  CNStageIntLLRInputS4xD(59)(3) <= VNStageIntLLROutputS3xD(214)(1);
  CNStageIntLLRInputS4xD(145)(3) <= VNStageIntLLROutputS3xD(214)(2);
  CNStageIntLLRInputS4xD(220)(3) <= VNStageIntLLROutputS3xD(214)(3);
  CNStageIntLLRInputS4xD(240)(3) <= VNStageIntLLROutputS3xD(214)(4);
  CNStageIntLLRInputS4xD(308)(3) <= VNStageIntLLROutputS3xD(214)(5);
  CNStageIntLLRInputS4xD(369)(3) <= VNStageIntLLROutputS3xD(214)(6);
  CNStageIntLLRInputS4xD(31)(3) <= VNStageIntLLROutputS3xD(215)(0);
  CNStageIntLLRInputS4xD(85)(3) <= VNStageIntLLROutputS3xD(215)(1);
  CNStageIntLLRInputS4xD(130)(3) <= VNStageIntLLROutputS3xD(215)(2);
  CNStageIntLLRInputS4xD(216)(3) <= VNStageIntLLROutputS3xD(215)(3);
  CNStageIntLLRInputS4xD(234)(3) <= VNStageIntLLROutputS3xD(215)(4);
  CNStageIntLLRInputS4xD(311)(3) <= VNStageIntLLROutputS3xD(215)(5);
  CNStageIntLLRInputS4xD(377)(3) <= VNStageIntLLROutputS3xD(215)(6);
  CNStageIntLLRInputS4xD(30)(3) <= VNStageIntLLROutputS3xD(216)(0);
  CNStageIntLLRInputS4xD(91)(3) <= VNStageIntLLROutputS3xD(216)(1);
  CNStageIntLLRInputS4xD(164)(3) <= VNStageIntLLROutputS3xD(216)(2);
  CNStageIntLLRInputS4xD(183)(3) <= VNStageIntLLROutputS3xD(216)(3);
  CNStageIntLLRInputS4xD(237)(3) <= VNStageIntLLROutputS3xD(216)(4);
  CNStageIntLLRInputS4xD(299)(3) <= VNStageIntLLROutputS3xD(216)(5);
  CNStageIntLLRInputS4xD(341)(3) <= VNStageIntLLROutputS3xD(216)(6);
  CNStageIntLLRInputS4xD(29)(3) <= VNStageIntLLROutputS3xD(217)(0);
  CNStageIntLLRInputS4xD(75)(3) <= VNStageIntLLROutputS3xD(217)(1);
  CNStageIntLLRInputS4xD(126)(3) <= VNStageIntLLROutputS3xD(217)(2);
  CNStageIntLLRInputS4xD(201)(3) <= VNStageIntLLROutputS3xD(217)(3);
  CNStageIntLLRInputS4xD(227)(3) <= VNStageIntLLROutputS3xD(217)(4);
  CNStageIntLLRInputS4xD(329)(3) <= VNStageIntLLROutputS3xD(217)(5);
  CNStageIntLLRInputS4xD(339)(3) <= VNStageIntLLROutputS3xD(217)(6);
  CNStageIntLLRInputS4xD(28)(3) <= VNStageIntLLROutputS3xD(218)(0);
  CNStageIntLLRInputS4xD(77)(3) <= VNStageIntLLROutputS3xD(218)(1);
  CNStageIntLLRInputS4xD(154)(3) <= VNStageIntLLROutputS3xD(218)(2);
  CNStageIntLLRInputS4xD(202)(3) <= VNStageIntLLROutputS3xD(218)(3);
  CNStageIntLLRInputS4xD(261)(3) <= VNStageIntLLROutputS3xD(218)(4);
  CNStageIntLLRInputS4xD(295)(3) <= VNStageIntLLROutputS3xD(218)(5);
  CNStageIntLLRInputS4xD(375)(3) <= VNStageIntLLROutputS3xD(218)(6);
  CNStageIntLLRInputS4xD(27)(3) <= VNStageIntLLROutputS3xD(219)(0);
  CNStageIntLLRInputS4xD(101)(3) <= VNStageIntLLROutputS3xD(219)(1);
  CNStageIntLLRInputS4xD(138)(3) <= VNStageIntLLROutputS3xD(219)(2);
  CNStageIntLLRInputS4xD(182)(3) <= VNStageIntLLROutputS3xD(219)(3);
  CNStageIntLLRInputS4xD(321)(3) <= VNStageIntLLROutputS3xD(219)(4);
  CNStageIntLLRInputS4xD(354)(3) <= VNStageIntLLROutputS3xD(219)(5);
  CNStageIntLLRInputS4xD(26)(3) <= VNStageIntLLROutputS3xD(220)(0);
  CNStageIntLLRInputS4xD(83)(3) <= VNStageIntLLROutputS3xD(220)(1);
  CNStageIntLLRInputS4xD(166)(3) <= VNStageIntLLROutputS3xD(220)(2);
  CNStageIntLLRInputS4xD(173)(3) <= VNStageIntLLROutputS3xD(220)(3);
  CNStageIntLLRInputS4xD(256)(3) <= VNStageIntLLROutputS3xD(220)(4);
  CNStageIntLLRInputS4xD(305)(3) <= VNStageIntLLROutputS3xD(220)(5);
  CNStageIntLLRInputS4xD(356)(3) <= VNStageIntLLROutputS3xD(220)(6);
  CNStageIntLLRInputS4xD(25)(3) <= VNStageIntLLROutputS3xD(221)(0);
  CNStageIntLLRInputS4xD(94)(3) <= VNStageIntLLROutputS3xD(221)(1);
  CNStageIntLLRInputS4xD(156)(3) <= VNStageIntLLROutputS3xD(221)(2);
  CNStageIntLLRInputS4xD(190)(3) <= VNStageIntLLROutputS3xD(221)(3);
  CNStageIntLLRInputS4xD(268)(3) <= VNStageIntLLROutputS3xD(221)(4);
  CNStageIntLLRInputS4xD(331)(3) <= VNStageIntLLROutputS3xD(221)(5);
  CNStageIntLLRInputS4xD(342)(3) <= VNStageIntLLROutputS3xD(221)(6);
  CNStageIntLLRInputS4xD(24)(3) <= VNStageIntLLROutputS3xD(222)(0);
  CNStageIntLLRInputS4xD(143)(3) <= VNStageIntLLROutputS3xD(222)(1);
  CNStageIntLLRInputS4xD(241)(3) <= VNStageIntLLROutputS3xD(222)(2);
  CNStageIntLLRInputS4xD(376)(3) <= VNStageIntLLROutputS3xD(222)(3);
  CNStageIntLLRInputS4xD(23)(3) <= VNStageIntLLROutputS3xD(223)(0);
  CNStageIntLLRInputS4xD(76)(3) <= VNStageIntLLROutputS3xD(223)(1);
  CNStageIntLLRInputS4xD(162)(3) <= VNStageIntLLROutputS3xD(223)(2);
  CNStageIntLLRInputS4xD(224)(3) <= VNStageIntLLROutputS3xD(223)(3);
  CNStageIntLLRInputS4xD(229)(3) <= VNStageIntLLROutputS3xD(223)(4);
  CNStageIntLLRInputS4xD(309)(3) <= VNStageIntLLROutputS3xD(223)(5);
  CNStageIntLLRInputS4xD(338)(3) <= VNStageIntLLROutputS3xD(223)(6);
  CNStageIntLLRInputS4xD(22)(3) <= VNStageIntLLROutputS3xD(224)(0);
  CNStageIntLLRInputS4xD(90)(3) <= VNStageIntLLROutputS3xD(224)(1);
  CNStageIntLLRInputS4xD(135)(3) <= VNStageIntLLROutputS3xD(224)(2);
  CNStageIntLLRInputS4xD(193)(3) <= VNStageIntLLROutputS3xD(224)(3);
  CNStageIntLLRInputS4xD(270)(3) <= VNStageIntLLROutputS3xD(224)(4);
  CNStageIntLLRInputS4xD(328)(3) <= VNStageIntLLROutputS3xD(224)(5);
  CNStageIntLLRInputS4xD(366)(3) <= VNStageIntLLROutputS3xD(224)(6);
  CNStageIntLLRInputS4xD(21)(3) <= VNStageIntLLROutputS3xD(225)(0);
  CNStageIntLLRInputS4xD(61)(3) <= VNStageIntLLROutputS3xD(225)(1);
  CNStageIntLLRInputS4xD(132)(3) <= VNStageIntLLROutputS3xD(225)(2);
  CNStageIntLLRInputS4xD(188)(3) <= VNStageIntLLROutputS3xD(225)(3);
  CNStageIntLLRInputS4xD(232)(3) <= VNStageIntLLROutputS3xD(225)(4);
  CNStageIntLLRInputS4xD(301)(3) <= VNStageIntLLROutputS3xD(225)(5);
  CNStageIntLLRInputS4xD(20)(3) <= VNStageIntLLROutputS3xD(226)(0);
  CNStageIntLLRInputS4xD(148)(3) <= VNStageIntLLROutputS3xD(226)(1);
  CNStageIntLLRInputS4xD(378)(3) <= VNStageIntLLROutputS3xD(226)(2);
  CNStageIntLLRInputS4xD(19)(3) <= VNStageIntLLROutputS3xD(227)(0);
  CNStageIntLLRInputS4xD(63)(3) <= VNStageIntLLROutputS3xD(227)(1);
  CNStageIntLLRInputS4xD(140)(3) <= VNStageIntLLROutputS3xD(227)(2);
  CNStageIntLLRInputS4xD(178)(3) <= VNStageIntLLROutputS3xD(227)(3);
  CNStageIntLLRInputS4xD(258)(3) <= VNStageIntLLROutputS3xD(227)(4);
  CNStageIntLLRInputS4xD(314)(3) <= VNStageIntLLROutputS3xD(227)(5);
  CNStageIntLLRInputS4xD(368)(3) <= VNStageIntLLROutputS3xD(227)(6);
  CNStageIntLLRInputS4xD(18)(3) <= VNStageIntLLROutputS3xD(228)(0);
  CNStageIntLLRInputS4xD(78)(3) <= VNStageIntLLROutputS3xD(228)(1);
  CNStageIntLLRInputS4xD(114)(3) <= VNStageIntLLROutputS3xD(228)(2);
  CNStageIntLLRInputS4xD(198)(3) <= VNStageIntLLROutputS3xD(228)(3);
  CNStageIntLLRInputS4xD(253)(3) <= VNStageIntLLROutputS3xD(228)(4);
  CNStageIntLLRInputS4xD(307)(3) <= VNStageIntLLROutputS3xD(228)(5);
  CNStageIntLLRInputS4xD(17)(3) <= VNStageIntLLROutputS3xD(229)(0);
  CNStageIntLLRInputS4xD(74)(3) <= VNStageIntLLROutputS3xD(229)(1);
  CNStageIntLLRInputS4xD(124)(3) <= VNStageIntLLROutputS3xD(229)(2);
  CNStageIntLLRInputS4xD(259)(3) <= VNStageIntLLROutputS3xD(229)(3);
  CNStageIntLLRInputS4xD(374)(3) <= VNStageIntLLROutputS3xD(229)(4);
  CNStageIntLLRInputS4xD(16)(3) <= VNStageIntLLROutputS3xD(230)(0);
  CNStageIntLLRInputS4xD(118)(3) <= VNStageIntLLROutputS3xD(230)(1);
  CNStageIntLLRInputS4xD(176)(3) <= VNStageIntLLROutputS3xD(230)(2);
  CNStageIntLLRInputS4xD(249)(3) <= VNStageIntLLROutputS3xD(230)(3);
  CNStageIntLLRInputS4xD(293)(3) <= VNStageIntLLROutputS3xD(230)(4);
  CNStageIntLLRInputS4xD(347)(3) <= VNStageIntLLROutputS3xD(230)(5);
  CNStageIntLLRInputS4xD(15)(3) <= VNStageIntLLROutputS3xD(231)(0);
  CNStageIntLLRInputS4xD(56)(3) <= VNStageIntLLROutputS3xD(231)(1);
  CNStageIntLLRInputS4xD(209)(3) <= VNStageIntLLROutputS3xD(231)(2);
  CNStageIntLLRInputS4xD(272)(3) <= VNStageIntLLROutputS3xD(231)(3);
  CNStageIntLLRInputS4xD(287)(3) <= VNStageIntLLROutputS3xD(231)(4);
  CNStageIntLLRInputS4xD(344)(3) <= VNStageIntLLROutputS3xD(231)(5);
  CNStageIntLLRInputS4xD(14)(3) <= VNStageIntLLROutputS3xD(232)(0);
  CNStageIntLLRInputS4xD(57)(3) <= VNStageIntLLROutputS3xD(232)(1);
  CNStageIntLLRInputS4xD(212)(3) <= VNStageIntLLROutputS3xD(232)(2);
  CNStageIntLLRInputS4xD(278)(3) <= VNStageIntLLROutputS3xD(232)(3);
  CNStageIntLLRInputS4xD(291)(3) <= VNStageIntLLROutputS3xD(232)(4);
  CNStageIntLLRInputS4xD(359)(3) <= VNStageIntLLROutputS3xD(232)(5);
  CNStageIntLLRInputS4xD(13)(3) <= VNStageIntLLROutputS3xD(233)(0);
  CNStageIntLLRInputS4xD(92)(3) <= VNStageIntLLROutputS3xD(233)(1);
  CNStageIntLLRInputS4xD(149)(3) <= VNStageIntLLROutputS3xD(233)(2);
  CNStageIntLLRInputS4xD(263)(3) <= VNStageIntLLROutputS3xD(233)(3);
  CNStageIntLLRInputS4xD(352)(3) <= VNStageIntLLROutputS3xD(233)(4);
  CNStageIntLLRInputS4xD(12)(3) <= VNStageIntLLROutputS3xD(234)(0);
  CNStageIntLLRInputS4xD(84)(3) <= VNStageIntLLROutputS3xD(234)(1);
  CNStageIntLLRInputS4xD(131)(3) <= VNStageIntLLROutputS3xD(234)(2);
  CNStageIntLLRInputS4xD(177)(3) <= VNStageIntLLROutputS3xD(234)(3);
  CNStageIntLLRInputS4xD(265)(3) <= VNStageIntLLROutputS3xD(234)(4);
  CNStageIntLLRInputS4xD(315)(3) <= VNStageIntLLROutputS3xD(234)(5);
  CNStageIntLLRInputS4xD(100)(3) <= VNStageIntLLROutputS3xD(235)(0);
  CNStageIntLLRInputS4xD(144)(3) <= VNStageIntLLROutputS3xD(235)(1);
  CNStageIntLLRInputS4xD(196)(3) <= VNStageIntLLROutputS3xD(235)(2);
  CNStageIntLLRInputS4xD(235)(3) <= VNStageIntLLROutputS3xD(235)(3);
  CNStageIntLLRInputS4xD(336)(3) <= VNStageIntLLROutputS3xD(235)(4);
  CNStageIntLLRInputS4xD(11)(3) <= VNStageIntLLROutputS3xD(236)(0);
  CNStageIntLLRInputS4xD(104)(3) <= VNStageIntLLROutputS3xD(236)(1);
  CNStageIntLLRInputS4xD(155)(3) <= VNStageIntLLROutputS3xD(236)(2);
  CNStageIntLLRInputS4xD(221)(3) <= VNStageIntLLROutputS3xD(236)(3);
  CNStageIntLLRInputS4xD(271)(3) <= VNStageIntLLROutputS3xD(236)(4);
  CNStageIntLLRInputS4xD(310)(3) <= VNStageIntLLROutputS3xD(236)(5);
  CNStageIntLLRInputS4xD(10)(3) <= VNStageIntLLROutputS3xD(237)(0);
  CNStageIntLLRInputS4xD(110)(3) <= VNStageIntLLROutputS3xD(237)(1);
  CNStageIntLLRInputS4xD(125)(3) <= VNStageIntLLROutputS3xD(237)(2);
  CNStageIntLLRInputS4xD(228)(3) <= VNStageIntLLROutputS3xD(237)(3);
  CNStageIntLLRInputS4xD(322)(3) <= VNStageIntLLROutputS3xD(237)(4);
  CNStageIntLLRInputS4xD(334)(3) <= VNStageIntLLROutputS3xD(237)(5);
  CNStageIntLLRInputS4xD(9)(3) <= VNStageIntLLROutputS3xD(238)(0);
  CNStageIntLLRInputS4xD(103)(3) <= VNStageIntLLROutputS3xD(238)(1);
  CNStageIntLLRInputS4xD(113)(3) <= VNStageIntLLROutputS3xD(238)(2);
  CNStageIntLLRInputS4xD(179)(3) <= VNStageIntLLROutputS3xD(238)(3);
  CNStageIntLLRInputS4xD(236)(3) <= VNStageIntLLROutputS3xD(238)(4);
  CNStageIntLLRInputS4xD(294)(3) <= VNStageIntLLROutputS3xD(238)(5);
  CNStageIntLLRInputS4xD(383)(3) <= VNStageIntLLROutputS3xD(238)(6);
  CNStageIntLLRInputS4xD(8)(3) <= VNStageIntLLROutputS3xD(239)(0);
  CNStageIntLLRInputS4xD(98)(3) <= VNStageIntLLROutputS3xD(239)(1);
  CNStageIntLLRInputS4xD(158)(3) <= VNStageIntLLROutputS3xD(239)(2);
  CNStageIntLLRInputS4xD(223)(3) <= VNStageIntLLROutputS3xD(239)(3);
  CNStageIntLLRInputS4xD(264)(3) <= VNStageIntLLROutputS3xD(239)(4);
  CNStageIntLLRInputS4xD(284)(3) <= VNStageIntLLROutputS3xD(239)(5);
  CNStageIntLLRInputS4xD(360)(3) <= VNStageIntLLROutputS3xD(239)(6);
  CNStageIntLLRInputS4xD(7)(3) <= VNStageIntLLROutputS3xD(240)(0);
  CNStageIntLLRInputS4xD(81)(3) <= VNStageIntLLROutputS3xD(240)(1);
  CNStageIntLLRInputS4xD(116)(3) <= VNStageIntLLROutputS3xD(240)(2);
  CNStageIntLLRInputS4xD(210)(3) <= VNStageIntLLROutputS3xD(240)(3);
  CNStageIntLLRInputS4xD(277)(3) <= VNStageIntLLROutputS3xD(240)(4);
  CNStageIntLLRInputS4xD(324)(3) <= VNStageIntLLROutputS3xD(240)(5);
  CNStageIntLLRInputS4xD(343)(3) <= VNStageIntLLROutputS3xD(240)(6);
  CNStageIntLLRInputS4xD(6)(3) <= VNStageIntLLROutputS3xD(241)(0);
  CNStageIntLLRInputS4xD(88)(3) <= VNStageIntLLROutputS3xD(241)(1);
  CNStageIntLLRInputS4xD(175)(3) <= VNStageIntLLROutputS3xD(241)(2);
  CNStageIntLLRInputS4xD(250)(3) <= VNStageIntLLROutputS3xD(241)(3);
  CNStageIntLLRInputS4xD(285)(3) <= VNStageIntLLROutputS3xD(241)(4);
  CNStageIntLLRInputS4xD(355)(3) <= VNStageIntLLROutputS3xD(241)(5);
  CNStageIntLLRInputS4xD(5)(3) <= VNStageIntLLROutputS3xD(242)(0);
  CNStageIntLLRInputS4xD(108)(3) <= VNStageIntLLROutputS3xD(242)(1);
  CNStageIntLLRInputS4xD(146)(3) <= VNStageIntLLROutputS3xD(242)(2);
  CNStageIntLLRInputS4xD(203)(3) <= VNStageIntLLROutputS3xD(242)(3);
  CNStageIntLLRInputS4xD(231)(3) <= VNStageIntLLROutputS3xD(242)(4);
  CNStageIntLLRInputS4xD(303)(3) <= VNStageIntLLROutputS3xD(242)(5);
  CNStageIntLLRInputS4xD(367)(3) <= VNStageIntLLROutputS3xD(242)(6);
  CNStageIntLLRInputS4xD(4)(3) <= VNStageIntLLROutputS3xD(243)(0);
  CNStageIntLLRInputS4xD(106)(3) <= VNStageIntLLROutputS3xD(243)(1);
  CNStageIntLLRInputS4xD(141)(3) <= VNStageIntLLROutputS3xD(243)(2);
  CNStageIntLLRInputS4xD(200)(3) <= VNStageIntLLROutputS3xD(243)(3);
  CNStageIntLLRInputS4xD(252)(3) <= VNStageIntLLROutputS3xD(243)(4);
  CNStageIntLLRInputS4xD(312)(3) <= VNStageIntLLROutputS3xD(243)(5);
  CNStageIntLLRInputS4xD(337)(3) <= VNStageIntLLROutputS3xD(243)(6);
  CNStageIntLLRInputS4xD(147)(3) <= VNStageIntLLROutputS3xD(244)(0);
  CNStageIntLLRInputS4xD(266)(3) <= VNStageIntLLROutputS3xD(244)(1);
  CNStageIntLLRInputS4xD(3)(3) <= VNStageIntLLROutputS3xD(245)(0);
  CNStageIntLLRInputS4xD(66)(3) <= VNStageIntLLROutputS3xD(245)(1);
  CNStageIntLLRInputS4xD(136)(3) <= VNStageIntLLROutputS3xD(245)(2);
  CNStageIntLLRInputS4xD(207)(3) <= VNStageIntLLROutputS3xD(245)(3);
  CNStageIntLLRInputS4xD(262)(3) <= VNStageIntLLROutputS3xD(245)(4);
  CNStageIntLLRInputS4xD(313)(3) <= VNStageIntLLROutputS3xD(245)(5);
  CNStageIntLLRInputS4xD(370)(3) <= VNStageIntLLROutputS3xD(245)(6);
  CNStageIntLLRInputS4xD(2)(3) <= VNStageIntLLROutputS3xD(246)(0);
  CNStageIntLLRInputS4xD(69)(3) <= VNStageIntLLROutputS3xD(246)(1);
  CNStageIntLLRInputS4xD(161)(3) <= VNStageIntLLROutputS3xD(246)(2);
  CNStageIntLLRInputS4xD(185)(3) <= VNStageIntLLROutputS3xD(246)(3);
  CNStageIntLLRInputS4xD(226)(3) <= VNStageIntLLROutputS3xD(246)(4);
  CNStageIntLLRInputS4xD(302)(3) <= VNStageIntLLROutputS3xD(246)(5);
  CNStageIntLLRInputS4xD(1)(3) <= VNStageIntLLROutputS3xD(247)(0);
  CNStageIntLLRInputS4xD(109)(3) <= VNStageIntLLROutputS3xD(247)(1);
  CNStageIntLLRInputS4xD(168)(3) <= VNStageIntLLROutputS3xD(247)(2);
  CNStageIntLLRInputS4xD(194)(3) <= VNStageIntLLROutputS3xD(247)(3);
  CNStageIntLLRInputS4xD(247)(3) <= VNStageIntLLROutputS3xD(247)(4);
  CNStageIntLLRInputS4xD(327)(3) <= VNStageIntLLROutputS3xD(247)(5);
  CNStageIntLLRInputS4xD(349)(3) <= VNStageIntLLROutputS3xD(247)(6);
  CNStageIntLLRInputS4xD(0)(3) <= VNStageIntLLROutputS3xD(248)(0);
  CNStageIntLLRInputS4xD(87)(3) <= VNStageIntLLROutputS3xD(248)(1);
  CNStageIntLLRInputS4xD(151)(3) <= VNStageIntLLROutputS3xD(248)(2);
  CNStageIntLLRInputS4xD(189)(3) <= VNStageIntLLROutputS3xD(248)(3);
  CNStageIntLLRInputS4xD(248)(3) <= VNStageIntLLROutputS3xD(248)(4);
  CNStageIntLLRInputS4xD(280)(3) <= VNStageIntLLROutputS3xD(248)(5);
  CNStageIntLLRInputS4xD(357)(3) <= VNStageIntLLROutputS3xD(248)(6);
  CNStageIntLLRInputS4xD(152)(3) <= VNStageIntLLROutputS3xD(249)(0);
  CNStageIntLLRInputS4xD(192)(3) <= VNStageIntLLROutputS3xD(249)(1);
  CNStageIntLLRInputS4xD(225)(3) <= VNStageIntLLROutputS3xD(249)(2);
  CNStageIntLLRInputS4xD(317)(3) <= VNStageIntLLROutputS3xD(249)(3);
  CNStageIntLLRInputS4xD(353)(3) <= VNStageIntLLROutputS3xD(249)(4);
  CNStageIntLLRInputS4xD(79)(3) <= VNStageIntLLROutputS3xD(250)(0);
  CNStageIntLLRInputS4xD(120)(3) <= VNStageIntLLROutputS3xD(250)(1);
  CNStageIntLLRInputS4xD(184)(3) <= VNStageIntLLROutputS3xD(250)(2);
  CNStageIntLLRInputS4xD(319)(3) <= VNStageIntLLROutputS3xD(250)(3);
  CNStageIntLLRInputS4xD(358)(3) <= VNStageIntLLROutputS3xD(250)(4);
  CNStageIntLLRInputS4xD(62)(3) <= VNStageIntLLROutputS3xD(251)(0);
  CNStageIntLLRInputS4xD(159)(3) <= VNStageIntLLROutputS3xD(251)(1);
  CNStageIntLLRInputS4xD(215)(3) <= VNStageIntLLROutputS3xD(251)(2);
  CNStageIntLLRInputS4xD(289)(3) <= VNStageIntLLROutputS3xD(251)(3);
  CNStageIntLLRInputS4xD(348)(3) <= VNStageIntLLROutputS3xD(251)(4);
  CNStageIntLLRInputS4xD(89)(3) <= VNStageIntLLROutputS3xD(252)(0);
  CNStageIntLLRInputS4xD(112)(3) <= VNStageIntLLROutputS3xD(252)(1);
  CNStageIntLLRInputS4xD(199)(3) <= VNStageIntLLROutputS3xD(252)(2);
  CNStageIntLLRInputS4xD(239)(3) <= VNStageIntLLROutputS3xD(252)(3);
  CNStageIntLLRInputS4xD(325)(3) <= VNStageIntLLROutputS3xD(252)(4);
  CNStageIntLLRInputS4xD(373)(3) <= VNStageIntLLROutputS3xD(252)(5);
  CNStageIntLLRInputS4xD(80)(3) <= VNStageIntLLROutputS3xD(253)(0);
  CNStageIntLLRInputS4xD(121)(3) <= VNStageIntLLROutputS3xD(253)(1);
  CNStageIntLLRInputS4xD(211)(3) <= VNStageIntLLROutputS3xD(253)(2);
  CNStageIntLLRInputS4xD(279)(3) <= VNStageIntLLROutputS3xD(253)(3);
  CNStageIntLLRInputS4xD(283)(3) <= VNStageIntLLROutputS3xD(253)(4);
  CNStageIntLLRInputS4xD(380)(3) <= VNStageIntLLROutputS3xD(253)(5);
  CNStageIntLLRInputS4xD(67)(3) <= VNStageIntLLROutputS3xD(254)(0);
  CNStageIntLLRInputS4xD(222)(3) <= VNStageIntLLROutputS3xD(254)(1);
  CNStageIntLLRInputS4xD(238)(3) <= VNStageIntLLROutputS3xD(254)(2);
  CNStageIntLLRInputS4xD(290)(3) <= VNStageIntLLROutputS3xD(254)(3);
  CNStageIntLLRInputS4xD(362)(3) <= VNStageIntLLROutputS3xD(254)(4);
  CNStageIntLLRInputS4xD(52)(3) <= VNStageIntLLROutputS3xD(255)(0);
  CNStageIntLLRInputS4xD(86)(3) <= VNStageIntLLROutputS3xD(255)(1);
  CNStageIntLLRInputS4xD(167)(3) <= VNStageIntLLROutputS3xD(255)(2);
  CNStageIntLLRInputS4xD(195)(3) <= VNStageIntLLROutputS3xD(255)(3);
  CNStageIntLLRInputS4xD(233)(3) <= VNStageIntLLROutputS3xD(255)(4);
  CNStageIntLLRInputS4xD(318)(3) <= VNStageIntLLROutputS3xD(255)(5);
  CNStageIntLLRInputS4xD(364)(3) <= VNStageIntLLROutputS3xD(255)(6);
  CNStageIntLLRInputS4xD(53)(4) <= VNStageIntLLROutputS3xD(256)(0);
  CNStageIntLLRInputS4xD(106)(4) <= VNStageIntLLROutputS3xD(256)(1);
  CNStageIntLLRInputS4xD(127)(4) <= VNStageIntLLROutputS3xD(256)(2);
  CNStageIntLLRInputS4xD(242)(4) <= VNStageIntLLROutputS3xD(256)(3);
  CNStageIntLLRInputS4xD(296)(4) <= VNStageIntLLROutputS3xD(256)(4);
  CNStageIntLLRInputS4xD(339)(4) <= VNStageIntLLROutputS3xD(256)(5);
  CNStageIntLLRInputS4xD(51)(4) <= VNStageIntLLROutputS3xD(257)(0);
  CNStageIntLLRInputS4xD(85)(4) <= VNStageIntLLROutputS3xD(257)(1);
  CNStageIntLLRInputS4xD(166)(4) <= VNStageIntLLROutputS3xD(257)(2);
  CNStageIntLLRInputS4xD(194)(4) <= VNStageIntLLROutputS3xD(257)(3);
  CNStageIntLLRInputS4xD(232)(4) <= VNStageIntLLROutputS3xD(257)(4);
  CNStageIntLLRInputS4xD(317)(4) <= VNStageIntLLROutputS3xD(257)(5);
  CNStageIntLLRInputS4xD(363)(4) <= VNStageIntLLROutputS3xD(257)(6);
  CNStageIntLLRInputS4xD(50)(4) <= VNStageIntLLROutputS3xD(258)(0);
  CNStageIntLLRInputS4xD(57)(4) <= VNStageIntLLROutputS3xD(258)(1);
  CNStageIntLLRInputS4xD(331)(4) <= VNStageIntLLROutputS3xD(258)(2);
  CNStageIntLLRInputS4xD(54)(4) <= VNStageIntLLROutputS3xD(259)(0);
  CNStageIntLLRInputS4xD(114)(4) <= VNStageIntLLROutputS3xD(259)(1);
  CNStageIntLLRInputS4xD(274)(4) <= VNStageIntLLROutputS3xD(259)(2);
  CNStageIntLLRInputS4xD(303)(4) <= VNStageIntLLROutputS3xD(259)(3);
  CNStageIntLLRInputS4xD(370)(4) <= VNStageIntLLROutputS3xD(259)(4);
  CNStageIntLLRInputS4xD(49)(4) <= VNStageIntLLROutputS3xD(260)(0);
  CNStageIntLLRInputS4xD(71)(4) <= VNStageIntLLROutputS3xD(260)(1);
  CNStageIntLLRInputS4xD(138)(4) <= VNStageIntLLROutputS3xD(260)(2);
  CNStageIntLLRInputS4xD(186)(4) <= VNStageIntLLROutputS3xD(260)(3);
  CNStageIntLLRInputS4xD(243)(4) <= VNStageIntLLROutputS3xD(260)(4);
  CNStageIntLLRInputS4xD(383)(4) <= VNStageIntLLROutputS3xD(260)(5);
  CNStageIntLLRInputS4xD(48)(4) <= VNStageIntLLROutputS3xD(261)(0);
  CNStageIntLLRInputS4xD(63)(4) <= VNStageIntLLROutputS3xD(261)(1);
  CNStageIntLLRInputS4xD(152)(4) <= VNStageIntLLROutputS3xD(261)(2);
  CNStageIntLLRInputS4xD(204)(4) <= VNStageIntLLROutputS3xD(261)(3);
  CNStageIntLLRInputS4xD(305)(4) <= VNStageIntLLROutputS3xD(261)(4);
  CNStageIntLLRInputS4xD(333)(4) <= VNStageIntLLROutputS3xD(261)(5);
  CNStageIntLLRInputS4xD(47)(4) <= VNStageIntLLROutputS3xD(262)(0);
  CNStageIntLLRInputS4xD(95)(4) <= VNStageIntLLROutputS3xD(262)(1);
  CNStageIntLLRInputS4xD(149)(4) <= VNStageIntLLROutputS3xD(262)(2);
  CNStageIntLLRInputS4xD(212)(4) <= VNStageIntLLROutputS3xD(262)(3);
  CNStageIntLLRInputS4xD(319)(4) <= VNStageIntLLROutputS3xD(262)(4);
  CNStageIntLLRInputS4xD(362)(4) <= VNStageIntLLROutputS3xD(262)(5);
  CNStageIntLLRInputS4xD(46)(4) <= VNStageIntLLROutputS3xD(263)(0);
  CNStageIntLLRInputS4xD(104)(4) <= VNStageIntLLROutputS3xD(263)(1);
  CNStageIntLLRInputS4xD(169)(4) <= VNStageIntLLROutputS3xD(263)(2);
  CNStageIntLLRInputS4xD(207)(4) <= VNStageIntLLROutputS3xD(263)(3);
  CNStageIntLLRInputS4xD(253)(4) <= VNStageIntLLROutputS3xD(263)(4);
  CNStageIntLLRInputS4xD(315)(4) <= VNStageIntLLROutputS3xD(263)(5);
  CNStageIntLLRInputS4xD(378)(4) <= VNStageIntLLROutputS3xD(263)(6);
  CNStageIntLLRInputS4xD(45)(4) <= VNStageIntLLROutputS3xD(264)(0);
  CNStageIntLLRInputS4xD(98)(4) <= VNStageIntLLROutputS3xD(264)(1);
  CNStageIntLLRInputS4xD(132)(4) <= VNStageIntLLROutputS3xD(264)(2);
  CNStageIntLLRInputS4xD(213)(4) <= VNStageIntLLROutputS3xD(264)(3);
  CNStageIntLLRInputS4xD(256)(4) <= VNStageIntLLROutputS3xD(264)(4);
  CNStageIntLLRInputS4xD(281)(4) <= VNStageIntLLROutputS3xD(264)(5);
  CNStageIntLLRInputS4xD(349)(4) <= VNStageIntLLROutputS3xD(264)(6);
  CNStageIntLLRInputS4xD(44)(4) <= VNStageIntLLROutputS3xD(265)(0);
  CNStageIntLLRInputS4xD(133)(4) <= VNStageIntLLROutputS3xD(265)(1);
  CNStageIntLLRInputS4xD(203)(4) <= VNStageIntLLROutputS3xD(265)(2);
  CNStageIntLLRInputS4xD(244)(4) <= VNStageIntLLROutputS3xD(265)(3);
  CNStageIntLLRInputS4xD(43)(4) <= VNStageIntLLROutputS3xD(266)(0);
  CNStageIntLLRInputS4xD(168)(4) <= VNStageIntLLROutputS3xD(266)(1);
  CNStageIntLLRInputS4xD(173)(4) <= VNStageIntLLROutputS3xD(266)(2);
  CNStageIntLLRInputS4xD(273)(4) <= VNStageIntLLROutputS3xD(266)(3);
  CNStageIntLLRInputS4xD(300)(4) <= VNStageIntLLROutputS3xD(266)(4);
  CNStageIntLLRInputS4xD(42)(4) <= VNStageIntLLROutputS3xD(267)(0);
  CNStageIntLLRInputS4xD(72)(4) <= VNStageIntLLROutputS3xD(267)(1);
  CNStageIntLLRInputS4xD(159)(4) <= VNStageIntLLROutputS3xD(267)(2);
  CNStageIntLLRInputS4xD(180)(4) <= VNStageIntLLROutputS3xD(267)(3);
  CNStageIntLLRInputS4xD(241)(4) <= VNStageIntLLROutputS3xD(267)(4);
  CNStageIntLLRInputS4xD(280)(4) <= VNStageIntLLROutputS3xD(267)(5);
  CNStageIntLLRInputS4xD(364)(4) <= VNStageIntLLROutputS3xD(267)(6);
  CNStageIntLLRInputS4xD(41)(4) <= VNStageIntLLROutputS3xD(268)(0);
  CNStageIntLLRInputS4xD(109)(4) <= VNStageIntLLROutputS3xD(268)(1);
  CNStageIntLLRInputS4xD(118)(4) <= VNStageIntLLROutputS3xD(268)(2);
  CNStageIntLLRInputS4xD(216)(4) <= VNStageIntLLROutputS3xD(268)(3);
  CNStageIntLLRInputS4xD(266)(4) <= VNStageIntLLROutputS3xD(268)(4);
  CNStageIntLLRInputS4xD(325)(4) <= VNStageIntLLROutputS3xD(268)(5);
  CNStageIntLLRInputS4xD(360)(4) <= VNStageIntLLROutputS3xD(268)(6);
  CNStageIntLLRInputS4xD(67)(4) <= VNStageIntLLROutputS3xD(269)(0);
  CNStageIntLLRInputS4xD(122)(4) <= VNStageIntLLROutputS3xD(269)(1);
  CNStageIntLLRInputS4xD(218)(4) <= VNStageIntLLROutputS3xD(269)(2);
  CNStageIntLLRInputS4xD(250)(4) <= VNStageIntLLROutputS3xD(269)(3);
  CNStageIntLLRInputS4xD(287)(4) <= VNStageIntLLROutputS3xD(269)(4);
  CNStageIntLLRInputS4xD(381)(4) <= VNStageIntLLROutputS3xD(269)(5);
  CNStageIntLLRInputS4xD(40)(4) <= VNStageIntLLROutputS3xD(270)(0);
  CNStageIntLLRInputS4xD(79)(4) <= VNStageIntLLROutputS3xD(270)(1);
  CNStageIntLLRInputS4xD(170)(4) <= VNStageIntLLROutputS3xD(270)(2);
  CNStageIntLLRInputS4xD(190)(4) <= VNStageIntLLROutputS3xD(270)(3);
  CNStageIntLLRInputS4xD(275)(4) <= VNStageIntLLROutputS3xD(270)(4);
  CNStageIntLLRInputS4xD(292)(4) <= VNStageIntLLROutputS3xD(270)(5);
  CNStageIntLLRInputS4xD(344)(4) <= VNStageIntLLROutputS3xD(270)(6);
  CNStageIntLLRInputS4xD(39)(4) <= VNStageIntLLROutputS3xD(271)(0);
  CNStageIntLLRInputS4xD(105)(4) <= VNStageIntLLROutputS3xD(271)(1);
  CNStageIntLLRInputS4xD(171)(4) <= VNStageIntLLROutputS3xD(271)(2);
  CNStageIntLLRInputS4xD(268)(4) <= VNStageIntLLROutputS3xD(271)(3);
  CNStageIntLLRInputS4xD(332)(4) <= VNStageIntLLROutputS3xD(271)(4);
  CNStageIntLLRInputS4xD(345)(4) <= VNStageIntLLROutputS3xD(271)(5);
  CNStageIntLLRInputS4xD(38)(4) <= VNStageIntLLROutputS3xD(272)(0);
  CNStageIntLLRInputS4xD(94)(4) <= VNStageIntLLROutputS3xD(272)(1);
  CNStageIntLLRInputS4xD(116)(4) <= VNStageIntLLROutputS3xD(272)(2);
  CNStageIntLLRInputS4xD(184)(4) <= VNStageIntLLROutputS3xD(272)(3);
  CNStageIntLLRInputS4xD(254)(4) <= VNStageIntLLROutputS3xD(272)(4);
  CNStageIntLLRInputS4xD(291)(4) <= VNStageIntLLROutputS3xD(272)(5);
  CNStageIntLLRInputS4xD(380)(4) <= VNStageIntLLROutputS3xD(272)(6);
  CNStageIntLLRInputS4xD(37)(4) <= VNStageIntLLROutputS3xD(273)(0);
  CNStageIntLLRInputS4xD(81)(4) <= VNStageIntLLROutputS3xD(273)(1);
  CNStageIntLLRInputS4xD(156)(4) <= VNStageIntLLROutputS3xD(273)(2);
  CNStageIntLLRInputS4xD(272)(4) <= VNStageIntLLROutputS3xD(273)(3);
  CNStageIntLLRInputS4xD(285)(4) <= VNStageIntLLROutputS3xD(273)(4);
  CNStageIntLLRInputS4xD(371)(4) <= VNStageIntLLROutputS3xD(273)(5);
  CNStageIntLLRInputS4xD(36)(4) <= VNStageIntLLROutputS3xD(274)(0);
  CNStageIntLLRInputS4xD(164)(4) <= VNStageIntLLROutputS3xD(274)(1);
  CNStageIntLLRInputS4xD(217)(4) <= VNStageIntLLROutputS3xD(274)(2);
  CNStageIntLLRInputS4xD(248)(4) <= VNStageIntLLROutputS3xD(274)(3);
  CNStageIntLLRInputS4xD(35)(4) <= VNStageIntLLROutputS3xD(275)(0);
  CNStageIntLLRInputS4xD(59)(4) <= VNStageIntLLROutputS3xD(275)(1);
  CNStageIntLLRInputS4xD(128)(4) <= VNStageIntLLROutputS3xD(275)(2);
  CNStageIntLLRInputS4xD(179)(4) <= VNStageIntLLROutputS3xD(275)(3);
  CNStageIntLLRInputS4xD(329)(4) <= VNStageIntLLROutputS3xD(275)(4);
  CNStageIntLLRInputS4xD(34)(4) <= VNStageIntLLROutputS3xD(276)(0);
  CNStageIntLLRInputS4xD(69)(4) <= VNStageIntLLROutputS3xD(276)(1);
  CNStageIntLLRInputS4xD(126)(4) <= VNStageIntLLROutputS3xD(276)(2);
  CNStageIntLLRInputS4xD(205)(4) <= VNStageIntLLROutputS3xD(276)(3);
  CNStageIntLLRInputS4xD(259)(4) <= VNStageIntLLROutputS3xD(276)(4);
  CNStageIntLLRInputS4xD(297)(4) <= VNStageIntLLROutputS3xD(276)(5);
  CNStageIntLLRInputS4xD(33)(4) <= VNStageIntLLROutputS3xD(277)(0);
  CNStageIntLLRInputS4xD(64)(4) <= VNStageIntLLROutputS3xD(277)(1);
  CNStageIntLLRInputS4xD(162)(4) <= VNStageIntLLROutputS3xD(277)(2);
  CNStageIntLLRInputS4xD(185)(4) <= VNStageIntLLROutputS3xD(277)(3);
  CNStageIntLLRInputS4xD(252)(4) <= VNStageIntLLROutputS3xD(277)(4);
  CNStageIntLLRInputS4xD(295)(4) <= VNStageIntLLROutputS3xD(277)(5);
  CNStageIntLLRInputS4xD(334)(4) <= VNStageIntLLROutputS3xD(277)(6);
  CNStageIntLLRInputS4xD(32)(4) <= VNStageIntLLROutputS3xD(278)(0);
  CNStageIntLLRInputS4xD(70)(4) <= VNStageIntLLROutputS3xD(278)(1);
  CNStageIntLLRInputS4xD(141)(4) <= VNStageIntLLROutputS3xD(278)(2);
  CNStageIntLLRInputS4xD(229)(4) <= VNStageIntLLROutputS3xD(278)(3);
  CNStageIntLLRInputS4xD(328)(4) <= VNStageIntLLROutputS3xD(278)(4);
  CNStageIntLLRInputS4xD(31)(4) <= VNStageIntLLROutputS3xD(279)(0);
  CNStageIntLLRInputS4xD(58)(4) <= VNStageIntLLROutputS3xD(279)(1);
  CNStageIntLLRInputS4xD(144)(4) <= VNStageIntLLROutputS3xD(279)(2);
  CNStageIntLLRInputS4xD(219)(4) <= VNStageIntLLROutputS3xD(279)(3);
  CNStageIntLLRInputS4xD(239)(4) <= VNStageIntLLROutputS3xD(279)(4);
  CNStageIntLLRInputS4xD(368)(4) <= VNStageIntLLROutputS3xD(279)(5);
  CNStageIntLLRInputS4xD(30)(4) <= VNStageIntLLROutputS3xD(280)(0);
  CNStageIntLLRInputS4xD(84)(4) <= VNStageIntLLROutputS3xD(280)(1);
  CNStageIntLLRInputS4xD(129)(4) <= VNStageIntLLROutputS3xD(280)(2);
  CNStageIntLLRInputS4xD(215)(4) <= VNStageIntLLROutputS3xD(280)(3);
  CNStageIntLLRInputS4xD(233)(4) <= VNStageIntLLROutputS3xD(280)(4);
  CNStageIntLLRInputS4xD(310)(4) <= VNStageIntLLROutputS3xD(280)(5);
  CNStageIntLLRInputS4xD(376)(4) <= VNStageIntLLROutputS3xD(280)(6);
  CNStageIntLLRInputS4xD(29)(4) <= VNStageIntLLROutputS3xD(281)(0);
  CNStageIntLLRInputS4xD(90)(4) <= VNStageIntLLROutputS3xD(281)(1);
  CNStageIntLLRInputS4xD(163)(4) <= VNStageIntLLROutputS3xD(281)(2);
  CNStageIntLLRInputS4xD(182)(4) <= VNStageIntLLROutputS3xD(281)(3);
  CNStageIntLLRInputS4xD(236)(4) <= VNStageIntLLROutputS3xD(281)(4);
  CNStageIntLLRInputS4xD(298)(4) <= VNStageIntLLROutputS3xD(281)(5);
  CNStageIntLLRInputS4xD(340)(4) <= VNStageIntLLROutputS3xD(281)(6);
  CNStageIntLLRInputS4xD(28)(4) <= VNStageIntLLROutputS3xD(282)(0);
  CNStageIntLLRInputS4xD(74)(4) <= VNStageIntLLROutputS3xD(282)(1);
  CNStageIntLLRInputS4xD(125)(4) <= VNStageIntLLROutputS3xD(282)(2);
  CNStageIntLLRInputS4xD(200)(4) <= VNStageIntLLROutputS3xD(282)(3);
  CNStageIntLLRInputS4xD(226)(4) <= VNStageIntLLROutputS3xD(282)(4);
  CNStageIntLLRInputS4xD(338)(4) <= VNStageIntLLROutputS3xD(282)(5);
  CNStageIntLLRInputS4xD(27)(4) <= VNStageIntLLROutputS3xD(283)(0);
  CNStageIntLLRInputS4xD(76)(4) <= VNStageIntLLROutputS3xD(283)(1);
  CNStageIntLLRInputS4xD(153)(4) <= VNStageIntLLROutputS3xD(283)(2);
  CNStageIntLLRInputS4xD(201)(4) <= VNStageIntLLROutputS3xD(283)(3);
  CNStageIntLLRInputS4xD(260)(4) <= VNStageIntLLROutputS3xD(283)(4);
  CNStageIntLLRInputS4xD(294)(4) <= VNStageIntLLROutputS3xD(283)(5);
  CNStageIntLLRInputS4xD(374)(4) <= VNStageIntLLROutputS3xD(283)(6);
  CNStageIntLLRInputS4xD(26)(4) <= VNStageIntLLROutputS3xD(284)(0);
  CNStageIntLLRInputS4xD(100)(4) <= VNStageIntLLROutputS3xD(284)(1);
  CNStageIntLLRInputS4xD(137)(4) <= VNStageIntLLROutputS3xD(284)(2);
  CNStageIntLLRInputS4xD(181)(4) <= VNStageIntLLROutputS3xD(284)(3);
  CNStageIntLLRInputS4xD(245)(4) <= VNStageIntLLROutputS3xD(284)(4);
  CNStageIntLLRInputS4xD(320)(4) <= VNStageIntLLROutputS3xD(284)(5);
  CNStageIntLLRInputS4xD(353)(4) <= VNStageIntLLROutputS3xD(284)(6);
  CNStageIntLLRInputS4xD(25)(4) <= VNStageIntLLROutputS3xD(285)(0);
  CNStageIntLLRInputS4xD(82)(4) <= VNStageIntLLROutputS3xD(285)(1);
  CNStageIntLLRInputS4xD(165)(4) <= VNStageIntLLROutputS3xD(285)(2);
  CNStageIntLLRInputS4xD(172)(4) <= VNStageIntLLROutputS3xD(285)(3);
  CNStageIntLLRInputS4xD(255)(4) <= VNStageIntLLROutputS3xD(285)(4);
  CNStageIntLLRInputS4xD(304)(4) <= VNStageIntLLROutputS3xD(285)(5);
  CNStageIntLLRInputS4xD(355)(4) <= VNStageIntLLROutputS3xD(285)(6);
  CNStageIntLLRInputS4xD(24)(4) <= VNStageIntLLROutputS3xD(286)(0);
  CNStageIntLLRInputS4xD(93)(4) <= VNStageIntLLROutputS3xD(286)(1);
  CNStageIntLLRInputS4xD(155)(4) <= VNStageIntLLROutputS3xD(286)(2);
  CNStageIntLLRInputS4xD(189)(4) <= VNStageIntLLROutputS3xD(286)(3);
  CNStageIntLLRInputS4xD(267)(4) <= VNStageIntLLROutputS3xD(286)(4);
  CNStageIntLLRInputS4xD(330)(4) <= VNStageIntLLROutputS3xD(286)(5);
  CNStageIntLLRInputS4xD(341)(4) <= VNStageIntLLROutputS3xD(286)(6);
  CNStageIntLLRInputS4xD(23)(4) <= VNStageIntLLROutputS3xD(287)(0);
  CNStageIntLLRInputS4xD(101)(4) <= VNStageIntLLROutputS3xD(287)(1);
  CNStageIntLLRInputS4xD(142)(4) <= VNStageIntLLROutputS3xD(287)(2);
  CNStageIntLLRInputS4xD(193)(4) <= VNStageIntLLROutputS3xD(287)(3);
  CNStageIntLLRInputS4xD(240)(4) <= VNStageIntLLROutputS3xD(287)(4);
  CNStageIntLLRInputS4xD(322)(4) <= VNStageIntLLROutputS3xD(287)(5);
  CNStageIntLLRInputS4xD(375)(4) <= VNStageIntLLROutputS3xD(287)(6);
  CNStageIntLLRInputS4xD(22)(4) <= VNStageIntLLROutputS3xD(288)(0);
  CNStageIntLLRInputS4xD(75)(4) <= VNStageIntLLROutputS3xD(288)(1);
  CNStageIntLLRInputS4xD(161)(4) <= VNStageIntLLROutputS3xD(288)(2);
  CNStageIntLLRInputS4xD(224)(4) <= VNStageIntLLROutputS3xD(288)(3);
  CNStageIntLLRInputS4xD(228)(4) <= VNStageIntLLROutputS3xD(288)(4);
  CNStageIntLLRInputS4xD(308)(4) <= VNStageIntLLROutputS3xD(288)(5);
  CNStageIntLLRInputS4xD(337)(4) <= VNStageIntLLROutputS3xD(288)(6);
  CNStageIntLLRInputS4xD(21)(4) <= VNStageIntLLROutputS3xD(289)(0);
  CNStageIntLLRInputS4xD(89)(4) <= VNStageIntLLROutputS3xD(289)(1);
  CNStageIntLLRInputS4xD(134)(4) <= VNStageIntLLROutputS3xD(289)(2);
  CNStageIntLLRInputS4xD(192)(4) <= VNStageIntLLROutputS3xD(289)(3);
  CNStageIntLLRInputS4xD(269)(4) <= VNStageIntLLROutputS3xD(289)(4);
  CNStageIntLLRInputS4xD(327)(4) <= VNStageIntLLROutputS3xD(289)(5);
  CNStageIntLLRInputS4xD(365)(4) <= VNStageIntLLROutputS3xD(289)(6);
  CNStageIntLLRInputS4xD(20)(4) <= VNStageIntLLROutputS3xD(290)(0);
  CNStageIntLLRInputS4xD(60)(4) <= VNStageIntLLROutputS3xD(290)(1);
  CNStageIntLLRInputS4xD(131)(4) <= VNStageIntLLROutputS3xD(290)(2);
  CNStageIntLLRInputS4xD(187)(4) <= VNStageIntLLROutputS3xD(290)(3);
  CNStageIntLLRInputS4xD(231)(4) <= VNStageIntLLROutputS3xD(290)(4);
  CNStageIntLLRInputS4xD(350)(4) <= VNStageIntLLROutputS3xD(290)(5);
  CNStageIntLLRInputS4xD(19)(4) <= VNStageIntLLROutputS3xD(291)(0);
  CNStageIntLLRInputS4xD(96)(4) <= VNStageIntLLROutputS3xD(291)(1);
  CNStageIntLLRInputS4xD(147)(4) <= VNStageIntLLROutputS3xD(291)(2);
  CNStageIntLLRInputS4xD(223)(4) <= VNStageIntLLROutputS3xD(291)(3);
  CNStageIntLLRInputS4xD(249)(4) <= VNStageIntLLROutputS3xD(291)(4);
  CNStageIntLLRInputS4xD(377)(4) <= VNStageIntLLROutputS3xD(291)(5);
  CNStageIntLLRInputS4xD(18)(4) <= VNStageIntLLROutputS3xD(292)(0);
  CNStageIntLLRInputS4xD(62)(4) <= VNStageIntLLROutputS3xD(292)(1);
  CNStageIntLLRInputS4xD(139)(4) <= VNStageIntLLROutputS3xD(292)(2);
  CNStageIntLLRInputS4xD(177)(4) <= VNStageIntLLROutputS3xD(292)(3);
  CNStageIntLLRInputS4xD(257)(4) <= VNStageIntLLROutputS3xD(292)(4);
  CNStageIntLLRInputS4xD(313)(4) <= VNStageIntLLROutputS3xD(292)(5);
  CNStageIntLLRInputS4xD(367)(4) <= VNStageIntLLROutputS3xD(292)(6);
  CNStageIntLLRInputS4xD(17)(4) <= VNStageIntLLROutputS3xD(293)(0);
  CNStageIntLLRInputS4xD(77)(4) <= VNStageIntLLROutputS3xD(293)(1);
  CNStageIntLLRInputS4xD(113)(4) <= VNStageIntLLROutputS3xD(293)(2);
  CNStageIntLLRInputS4xD(197)(4) <= VNStageIntLLROutputS3xD(293)(3);
  CNStageIntLLRInputS4xD(306)(4) <= VNStageIntLLROutputS3xD(293)(4);
  CNStageIntLLRInputS4xD(354)(4) <= VNStageIntLLROutputS3xD(293)(5);
  CNStageIntLLRInputS4xD(16)(4) <= VNStageIntLLROutputS3xD(294)(0);
  CNStageIntLLRInputS4xD(73)(4) <= VNStageIntLLROutputS3xD(294)(1);
  CNStageIntLLRInputS4xD(123)(4) <= VNStageIntLLROutputS3xD(294)(2);
  CNStageIntLLRInputS4xD(196)(4) <= VNStageIntLLROutputS3xD(294)(3);
  CNStageIntLLRInputS4xD(258)(4) <= VNStageIntLLROutputS3xD(294)(4);
  CNStageIntLLRInputS4xD(284)(4) <= VNStageIntLLROutputS3xD(294)(5);
  CNStageIntLLRInputS4xD(373)(4) <= VNStageIntLLROutputS3xD(294)(6);
  CNStageIntLLRInputS4xD(15)(4) <= VNStageIntLLROutputS3xD(295)(0);
  CNStageIntLLRInputS4xD(92)(4) <= VNStageIntLLROutputS3xD(295)(1);
  CNStageIntLLRInputS4xD(117)(4) <= VNStageIntLLROutputS3xD(295)(2);
  CNStageIntLLRInputS4xD(175)(4) <= VNStageIntLLROutputS3xD(295)(3);
  CNStageIntLLRInputS4xD(346)(4) <= VNStageIntLLROutputS3xD(295)(4);
  CNStageIntLLRInputS4xD(14)(4) <= VNStageIntLLROutputS3xD(296)(0);
  CNStageIntLLRInputS4xD(55)(4) <= VNStageIntLLROutputS3xD(296)(1);
  CNStageIntLLRInputS4xD(121)(4) <= VNStageIntLLROutputS3xD(296)(2);
  CNStageIntLLRInputS4xD(208)(4) <= VNStageIntLLROutputS3xD(296)(3);
  CNStageIntLLRInputS4xD(286)(4) <= VNStageIntLLROutputS3xD(296)(4);
  CNStageIntLLRInputS4xD(343)(4) <= VNStageIntLLROutputS3xD(296)(5);
  CNStageIntLLRInputS4xD(13)(4) <= VNStageIntLLROutputS3xD(297)(0);
  CNStageIntLLRInputS4xD(56)(4) <= VNStageIntLLROutputS3xD(297)(1);
  CNStageIntLLRInputS4xD(111)(4) <= VNStageIntLLROutputS3xD(297)(2);
  CNStageIntLLRInputS4xD(211)(4) <= VNStageIntLLROutputS3xD(297)(3);
  CNStageIntLLRInputS4xD(277)(4) <= VNStageIntLLROutputS3xD(297)(4);
  CNStageIntLLRInputS4xD(290)(4) <= VNStageIntLLROutputS3xD(297)(5);
  CNStageIntLLRInputS4xD(358)(4) <= VNStageIntLLROutputS3xD(297)(6);
  CNStageIntLLRInputS4xD(12)(4) <= VNStageIntLLROutputS3xD(298)(0);
  CNStageIntLLRInputS4xD(91)(4) <= VNStageIntLLROutputS3xD(298)(1);
  CNStageIntLLRInputS4xD(148)(4) <= VNStageIntLLROutputS3xD(298)(2);
  CNStageIntLLRInputS4xD(198)(4) <= VNStageIntLLROutputS3xD(298)(3);
  CNStageIntLLRInputS4xD(262)(4) <= VNStageIntLLROutputS3xD(298)(4);
  CNStageIntLLRInputS4xD(282)(4) <= VNStageIntLLROutputS3xD(298)(5);
  CNStageIntLLRInputS4xD(351)(4) <= VNStageIntLLROutputS3xD(298)(6);
  CNStageIntLLRInputS4xD(83)(4) <= VNStageIntLLROutputS3xD(299)(0);
  CNStageIntLLRInputS4xD(130)(4) <= VNStageIntLLROutputS3xD(299)(1);
  CNStageIntLLRInputS4xD(176)(4) <= VNStageIntLLROutputS3xD(299)(2);
  CNStageIntLLRInputS4xD(264)(4) <= VNStageIntLLROutputS3xD(299)(3);
  CNStageIntLLRInputS4xD(314)(4) <= VNStageIntLLROutputS3xD(299)(4);
  CNStageIntLLRInputS4xD(11)(4) <= VNStageIntLLROutputS3xD(300)(0);
  CNStageIntLLRInputS4xD(99)(4) <= VNStageIntLLROutputS3xD(300)(1);
  CNStageIntLLRInputS4xD(143)(4) <= VNStageIntLLROutputS3xD(300)(2);
  CNStageIntLLRInputS4xD(195)(4) <= VNStageIntLLROutputS3xD(300)(3);
  CNStageIntLLRInputS4xD(299)(4) <= VNStageIntLLROutputS3xD(300)(4);
  CNStageIntLLRInputS4xD(335)(4) <= VNStageIntLLROutputS3xD(300)(5);
  CNStageIntLLRInputS4xD(10)(4) <= VNStageIntLLROutputS3xD(301)(0);
  CNStageIntLLRInputS4xD(103)(4) <= VNStageIntLLROutputS3xD(301)(1);
  CNStageIntLLRInputS4xD(154)(4) <= VNStageIntLLROutputS3xD(301)(2);
  CNStageIntLLRInputS4xD(220)(4) <= VNStageIntLLROutputS3xD(301)(3);
  CNStageIntLLRInputS4xD(270)(4) <= VNStageIntLLROutputS3xD(301)(4);
  CNStageIntLLRInputS4xD(309)(4) <= VNStageIntLLROutputS3xD(301)(5);
  CNStageIntLLRInputS4xD(9)(4) <= VNStageIntLLROutputS3xD(302)(0);
  CNStageIntLLRInputS4xD(110)(4) <= VNStageIntLLROutputS3xD(302)(1);
  CNStageIntLLRInputS4xD(124)(4) <= VNStageIntLLROutputS3xD(302)(2);
  CNStageIntLLRInputS4xD(206)(4) <= VNStageIntLLROutputS3xD(302)(3);
  CNStageIntLLRInputS4xD(227)(4) <= VNStageIntLLROutputS3xD(302)(4);
  CNStageIntLLRInputS4xD(321)(4) <= VNStageIntLLROutputS3xD(302)(5);
  CNStageIntLLRInputS4xD(8)(4) <= VNStageIntLLROutputS3xD(303)(0);
  CNStageIntLLRInputS4xD(102)(4) <= VNStageIntLLROutputS3xD(303)(1);
  CNStageIntLLRInputS4xD(112)(4) <= VNStageIntLLROutputS3xD(303)(2);
  CNStageIntLLRInputS4xD(178)(4) <= VNStageIntLLROutputS3xD(303)(3);
  CNStageIntLLRInputS4xD(235)(4) <= VNStageIntLLROutputS3xD(303)(4);
  CNStageIntLLRInputS4xD(293)(4) <= VNStageIntLLROutputS3xD(303)(5);
  CNStageIntLLRInputS4xD(382)(4) <= VNStageIntLLROutputS3xD(303)(6);
  CNStageIntLLRInputS4xD(7)(4) <= VNStageIntLLROutputS3xD(304)(0);
  CNStageIntLLRInputS4xD(97)(4) <= VNStageIntLLROutputS3xD(304)(1);
  CNStageIntLLRInputS4xD(157)(4) <= VNStageIntLLROutputS3xD(304)(2);
  CNStageIntLLRInputS4xD(222)(4) <= VNStageIntLLROutputS3xD(304)(3);
  CNStageIntLLRInputS4xD(263)(4) <= VNStageIntLLROutputS3xD(304)(4);
  CNStageIntLLRInputS4xD(283)(4) <= VNStageIntLLROutputS3xD(304)(5);
  CNStageIntLLRInputS4xD(359)(4) <= VNStageIntLLROutputS3xD(304)(6);
  CNStageIntLLRInputS4xD(6)(4) <= VNStageIntLLROutputS3xD(305)(0);
  CNStageIntLLRInputS4xD(80)(4) <= VNStageIntLLROutputS3xD(305)(1);
  CNStageIntLLRInputS4xD(115)(4) <= VNStageIntLLROutputS3xD(305)(2);
  CNStageIntLLRInputS4xD(209)(4) <= VNStageIntLLROutputS3xD(305)(3);
  CNStageIntLLRInputS4xD(276)(4) <= VNStageIntLLROutputS3xD(305)(4);
  CNStageIntLLRInputS4xD(323)(4) <= VNStageIntLLROutputS3xD(305)(5);
  CNStageIntLLRInputS4xD(342)(4) <= VNStageIntLLROutputS3xD(305)(6);
  CNStageIntLLRInputS4xD(5)(4) <= VNStageIntLLROutputS3xD(306)(0);
  CNStageIntLLRInputS4xD(87)(4) <= VNStageIntLLROutputS3xD(306)(1);
  CNStageIntLLRInputS4xD(136)(4) <= VNStageIntLLROutputS3xD(306)(2);
  CNStageIntLLRInputS4xD(174)(4) <= VNStageIntLLROutputS3xD(306)(3);
  CNStageIntLLRInputS4xD(4)(4) <= VNStageIntLLROutputS3xD(307)(0);
  CNStageIntLLRInputS4xD(107)(4) <= VNStageIntLLROutputS3xD(307)(1);
  CNStageIntLLRInputS4xD(145)(4) <= VNStageIntLLROutputS3xD(307)(2);
  CNStageIntLLRInputS4xD(202)(4) <= VNStageIntLLROutputS3xD(307)(3);
  CNStageIntLLRInputS4xD(230)(4) <= VNStageIntLLROutputS3xD(307)(4);
  CNStageIntLLRInputS4xD(302)(4) <= VNStageIntLLROutputS3xD(307)(5);
  CNStageIntLLRInputS4xD(366)(4) <= VNStageIntLLROutputS3xD(307)(6);
  CNStageIntLLRInputS4xD(140)(4) <= VNStageIntLLROutputS3xD(308)(0);
  CNStageIntLLRInputS4xD(199)(4) <= VNStageIntLLROutputS3xD(308)(1);
  CNStageIntLLRInputS4xD(251)(4) <= VNStageIntLLROutputS3xD(308)(2);
  CNStageIntLLRInputS4xD(311)(4) <= VNStageIntLLROutputS3xD(308)(3);
  CNStageIntLLRInputS4xD(336)(4) <= VNStageIntLLROutputS3xD(308)(4);
  CNStageIntLLRInputS4xD(3)(4) <= VNStageIntLLROutputS3xD(309)(0);
  CNStageIntLLRInputS4xD(86)(4) <= VNStageIntLLROutputS3xD(309)(1);
  CNStageIntLLRInputS4xD(146)(4) <= VNStageIntLLROutputS3xD(309)(2);
  CNStageIntLLRInputS4xD(214)(4) <= VNStageIntLLROutputS3xD(309)(3);
  CNStageIntLLRInputS4xD(265)(4) <= VNStageIntLLROutputS3xD(309)(4);
  CNStageIntLLRInputS4xD(307)(4) <= VNStageIntLLROutputS3xD(309)(5);
  CNStageIntLLRInputS4xD(2)(4) <= VNStageIntLLROutputS3xD(310)(0);
  CNStageIntLLRInputS4xD(65)(4) <= VNStageIntLLROutputS3xD(310)(1);
  CNStageIntLLRInputS4xD(135)(4) <= VNStageIntLLROutputS3xD(310)(2);
  CNStageIntLLRInputS4xD(261)(4) <= VNStageIntLLROutputS3xD(310)(3);
  CNStageIntLLRInputS4xD(312)(4) <= VNStageIntLLROutputS3xD(310)(4);
  CNStageIntLLRInputS4xD(369)(4) <= VNStageIntLLROutputS3xD(310)(5);
  CNStageIntLLRInputS4xD(1)(4) <= VNStageIntLLROutputS3xD(311)(0);
  CNStageIntLLRInputS4xD(68)(4) <= VNStageIntLLROutputS3xD(311)(1);
  CNStageIntLLRInputS4xD(160)(4) <= VNStageIntLLROutputS3xD(311)(2);
  CNStageIntLLRInputS4xD(225)(4) <= VNStageIntLLROutputS3xD(311)(3);
  CNStageIntLLRInputS4xD(301)(4) <= VNStageIntLLROutputS3xD(311)(4);
  CNStageIntLLRInputS4xD(0)(4) <= VNStageIntLLROutputS3xD(312)(0);
  CNStageIntLLRInputS4xD(108)(4) <= VNStageIntLLROutputS3xD(312)(1);
  CNStageIntLLRInputS4xD(167)(4) <= VNStageIntLLROutputS3xD(312)(2);
  CNStageIntLLRInputS4xD(246)(4) <= VNStageIntLLROutputS3xD(312)(3);
  CNStageIntLLRInputS4xD(326)(4) <= VNStageIntLLROutputS3xD(312)(4);
  CNStageIntLLRInputS4xD(348)(4) <= VNStageIntLLROutputS3xD(312)(5);
  CNStageIntLLRInputS4xD(150)(4) <= VNStageIntLLROutputS3xD(313)(0);
  CNStageIntLLRInputS4xD(188)(4) <= VNStageIntLLROutputS3xD(313)(1);
  CNStageIntLLRInputS4xD(247)(4) <= VNStageIntLLROutputS3xD(313)(2);
  CNStageIntLLRInputS4xD(356)(4) <= VNStageIntLLROutputS3xD(313)(3);
  CNStageIntLLRInputS4xD(191)(4) <= VNStageIntLLROutputS3xD(314)(0);
  CNStageIntLLRInputS4xD(278)(4) <= VNStageIntLLROutputS3xD(314)(1);
  CNStageIntLLRInputS4xD(316)(4) <= VNStageIntLLROutputS3xD(314)(2);
  CNStageIntLLRInputS4xD(352)(4) <= VNStageIntLLROutputS3xD(314)(3);
  CNStageIntLLRInputS4xD(78)(4) <= VNStageIntLLROutputS3xD(315)(0);
  CNStageIntLLRInputS4xD(119)(4) <= VNStageIntLLROutputS3xD(315)(1);
  CNStageIntLLRInputS4xD(183)(4) <= VNStageIntLLROutputS3xD(315)(2);
  CNStageIntLLRInputS4xD(271)(4) <= VNStageIntLLROutputS3xD(315)(3);
  CNStageIntLLRInputS4xD(318)(4) <= VNStageIntLLROutputS3xD(315)(4);
  CNStageIntLLRInputS4xD(357)(4) <= VNStageIntLLROutputS3xD(315)(5);
  CNStageIntLLRInputS4xD(61)(4) <= VNStageIntLLROutputS3xD(316)(0);
  CNStageIntLLRInputS4xD(158)(4) <= VNStageIntLLROutputS3xD(316)(1);
  CNStageIntLLRInputS4xD(234)(4) <= VNStageIntLLROutputS3xD(316)(2);
  CNStageIntLLRInputS4xD(288)(4) <= VNStageIntLLROutputS3xD(316)(3);
  CNStageIntLLRInputS4xD(347)(4) <= VNStageIntLLROutputS3xD(316)(4);
  CNStageIntLLRInputS4xD(88)(4) <= VNStageIntLLROutputS3xD(317)(0);
  CNStageIntLLRInputS4xD(238)(4) <= VNStageIntLLROutputS3xD(317)(1);
  CNStageIntLLRInputS4xD(324)(4) <= VNStageIntLLROutputS3xD(317)(2);
  CNStageIntLLRInputS4xD(372)(4) <= VNStageIntLLROutputS3xD(317)(3);
  CNStageIntLLRInputS4xD(120)(4) <= VNStageIntLLROutputS3xD(318)(0);
  CNStageIntLLRInputS4xD(210)(4) <= VNStageIntLLROutputS3xD(318)(1);
  CNStageIntLLRInputS4xD(279)(4) <= VNStageIntLLROutputS3xD(318)(2);
  CNStageIntLLRInputS4xD(379)(4) <= VNStageIntLLROutputS3xD(318)(3);
  CNStageIntLLRInputS4xD(52)(4) <= VNStageIntLLROutputS3xD(319)(0);
  CNStageIntLLRInputS4xD(66)(4) <= VNStageIntLLROutputS3xD(319)(1);
  CNStageIntLLRInputS4xD(151)(4) <= VNStageIntLLROutputS3xD(319)(2);
  CNStageIntLLRInputS4xD(221)(4) <= VNStageIntLLROutputS3xD(319)(3);
  CNStageIntLLRInputS4xD(237)(4) <= VNStageIntLLROutputS3xD(319)(4);
  CNStageIntLLRInputS4xD(289)(4) <= VNStageIntLLROutputS3xD(319)(5);
  CNStageIntLLRInputS4xD(361)(4) <= VNStageIntLLROutputS3xD(319)(6);
  CNStageIntLLRInputS4xD(53)(5) <= VNStageIntLLROutputS3xD(320)(0);
  CNStageIntLLRInputS4xD(126)(5) <= VNStageIntLLROutputS3xD(320)(1);
  CNStageIntLLRInputS4xD(196)(5) <= VNStageIntLLROutputS3xD(320)(2);
  CNStageIntLLRInputS4xD(295)(5) <= VNStageIntLLROutputS3xD(320)(3);
  CNStageIntLLRInputS4xD(338)(5) <= VNStageIntLLROutputS3xD(320)(4);
  CNStageIntLLRInputS4xD(51)(5) <= VNStageIntLLROutputS3xD(321)(0);
  CNStageIntLLRInputS4xD(65)(5) <= VNStageIntLLROutputS3xD(321)(1);
  CNStageIntLLRInputS4xD(150)(5) <= VNStageIntLLROutputS3xD(321)(2);
  CNStageIntLLRInputS4xD(220)(5) <= VNStageIntLLROutputS3xD(321)(3);
  CNStageIntLLRInputS4xD(236)(5) <= VNStageIntLLROutputS3xD(321)(4);
  CNStageIntLLRInputS4xD(288)(5) <= VNStageIntLLROutputS3xD(321)(5);
  CNStageIntLLRInputS4xD(360)(5) <= VNStageIntLLROutputS3xD(321)(6);
  CNStageIntLLRInputS4xD(50)(5) <= VNStageIntLLROutputS3xD(322)(0);
  CNStageIntLLRInputS4xD(84)(5) <= VNStageIntLLROutputS3xD(322)(1);
  CNStageIntLLRInputS4xD(165)(5) <= VNStageIntLLROutputS3xD(322)(2);
  CNStageIntLLRInputS4xD(231)(5) <= VNStageIntLLROutputS3xD(322)(3);
  CNStageIntLLRInputS4xD(316)(5) <= VNStageIntLLROutputS3xD(322)(4);
  CNStageIntLLRInputS4xD(362)(5) <= VNStageIntLLROutputS3xD(322)(5);
  CNStageIntLLRInputS4xD(56)(5) <= VNStageIntLLROutputS3xD(323)(0);
  CNStageIntLLRInputS4xD(136)(5) <= VNStageIntLLROutputS3xD(323)(1);
  CNStageIntLLRInputS4xD(184)(5) <= VNStageIntLLROutputS3xD(323)(2);
  CNStageIntLLRInputS4xD(268)(5) <= VNStageIntLLROutputS3xD(323)(3);
  CNStageIntLLRInputS4xD(330)(5) <= VNStageIntLLROutputS3xD(323)(4);
  CNStageIntLLRInputS4xD(49)(5) <= VNStageIntLLROutputS3xD(324)(0);
  CNStageIntLLRInputS4xD(109)(5) <= VNStageIntLLROutputS3xD(324)(1);
  CNStageIntLLRInputS4xD(113)(5) <= VNStageIntLLROutputS3xD(324)(2);
  CNStageIntLLRInputS4xD(223)(5) <= VNStageIntLLROutputS3xD(324)(3);
  CNStageIntLLRInputS4xD(273)(5) <= VNStageIntLLROutputS3xD(324)(4);
  CNStageIntLLRInputS4xD(302)(5) <= VNStageIntLLROutputS3xD(324)(5);
  CNStageIntLLRInputS4xD(369)(5) <= VNStageIntLLROutputS3xD(324)(6);
  CNStageIntLLRInputS4xD(48)(5) <= VNStageIntLLROutputS3xD(325)(0);
  CNStageIntLLRInputS4xD(70)(5) <= VNStageIntLLROutputS3xD(325)(1);
  CNStageIntLLRInputS4xD(137)(5) <= VNStageIntLLROutputS3xD(325)(2);
  CNStageIntLLRInputS4xD(185)(5) <= VNStageIntLLROutputS3xD(325)(3);
  CNStageIntLLRInputS4xD(242)(5) <= VNStageIntLLROutputS3xD(325)(4);
  CNStageIntLLRInputS4xD(284)(5) <= VNStageIntLLROutputS3xD(325)(5);
  CNStageIntLLRInputS4xD(382)(5) <= VNStageIntLLROutputS3xD(325)(6);
  CNStageIntLLRInputS4xD(47)(5) <= VNStageIntLLROutputS3xD(326)(0);
  CNStageIntLLRInputS4xD(62)(5) <= VNStageIntLLROutputS3xD(326)(1);
  CNStageIntLLRInputS4xD(203)(5) <= VNStageIntLLROutputS3xD(326)(2);
  CNStageIntLLRInputS4xD(241)(5) <= VNStageIntLLROutputS3xD(326)(3);
  CNStageIntLLRInputS4xD(304)(5) <= VNStageIntLLROutputS3xD(326)(4);
  CNStageIntLLRInputS4xD(46)(5) <= VNStageIntLLROutputS3xD(327)(0);
  CNStageIntLLRInputS4xD(94)(5) <= VNStageIntLLROutputS3xD(327)(1);
  CNStageIntLLRInputS4xD(148)(5) <= VNStageIntLLROutputS3xD(327)(2);
  CNStageIntLLRInputS4xD(211)(5) <= VNStageIntLLROutputS3xD(327)(3);
  CNStageIntLLRInputS4xD(272)(5) <= VNStageIntLLROutputS3xD(327)(4);
  CNStageIntLLRInputS4xD(318)(5) <= VNStageIntLLROutputS3xD(327)(5);
  CNStageIntLLRInputS4xD(361)(5) <= VNStageIntLLROutputS3xD(327)(6);
  CNStageIntLLRInputS4xD(45)(5) <= VNStageIntLLROutputS3xD(328)(0);
  CNStageIntLLRInputS4xD(103)(5) <= VNStageIntLLROutputS3xD(328)(1);
  CNStageIntLLRInputS4xD(168)(5) <= VNStageIntLLROutputS3xD(328)(2);
  CNStageIntLLRInputS4xD(314)(5) <= VNStageIntLLROutputS3xD(328)(3);
  CNStageIntLLRInputS4xD(377)(5) <= VNStageIntLLROutputS3xD(328)(4);
  CNStageIntLLRInputS4xD(44)(5) <= VNStageIntLLROutputS3xD(329)(0);
  CNStageIntLLRInputS4xD(97)(5) <= VNStageIntLLROutputS3xD(329)(1);
  CNStageIntLLRInputS4xD(131)(5) <= VNStageIntLLROutputS3xD(329)(2);
  CNStageIntLLRInputS4xD(212)(5) <= VNStageIntLLROutputS3xD(329)(3);
  CNStageIntLLRInputS4xD(255)(5) <= VNStageIntLLROutputS3xD(329)(4);
  CNStageIntLLRInputS4xD(280)(5) <= VNStageIntLLROutputS3xD(329)(5);
  CNStageIntLLRInputS4xD(348)(5) <= VNStageIntLLROutputS3xD(329)(6);
  CNStageIntLLRInputS4xD(43)(5) <= VNStageIntLLROutputS3xD(330)(0);
  CNStageIntLLRInputS4xD(101)(5) <= VNStageIntLLROutputS3xD(330)(1);
  CNStageIntLLRInputS4xD(132)(5) <= VNStageIntLLROutputS3xD(330)(2);
  CNStageIntLLRInputS4xD(202)(5) <= VNStageIntLLROutputS3xD(330)(3);
  CNStageIntLLRInputS4xD(243)(5) <= VNStageIntLLROutputS3xD(330)(4);
  CNStageIntLLRInputS4xD(42)(5) <= VNStageIntLLROutputS3xD(331)(0);
  CNStageIntLLRInputS4xD(92)(5) <= VNStageIntLLROutputS3xD(331)(1);
  CNStageIntLLRInputS4xD(167)(5) <= VNStageIntLLROutputS3xD(331)(2);
  CNStageIntLLRInputS4xD(172)(5) <= VNStageIntLLROutputS3xD(331)(3);
  CNStageIntLLRInputS4xD(350)(5) <= VNStageIntLLROutputS3xD(331)(4);
  CNStageIntLLRInputS4xD(41)(5) <= VNStageIntLLROutputS3xD(332)(0);
  CNStageIntLLRInputS4xD(71)(5) <= VNStageIntLLROutputS3xD(332)(1);
  CNStageIntLLRInputS4xD(158)(5) <= VNStageIntLLROutputS3xD(332)(2);
  CNStageIntLLRInputS4xD(179)(5) <= VNStageIntLLROutputS3xD(332)(3);
  CNStageIntLLRInputS4xD(240)(5) <= VNStageIntLLROutputS3xD(332)(4);
  CNStageIntLLRInputS4xD(363)(5) <= VNStageIntLLROutputS3xD(332)(5);
  CNStageIntLLRInputS4xD(108)(5) <= VNStageIntLLROutputS3xD(333)(0);
  CNStageIntLLRInputS4xD(117)(5) <= VNStageIntLLROutputS3xD(333)(1);
  CNStageIntLLRInputS4xD(215)(5) <= VNStageIntLLROutputS3xD(333)(2);
  CNStageIntLLRInputS4xD(265)(5) <= VNStageIntLLROutputS3xD(333)(3);
  CNStageIntLLRInputS4xD(324)(5) <= VNStageIntLLROutputS3xD(333)(4);
  CNStageIntLLRInputS4xD(359)(5) <= VNStageIntLLROutputS3xD(333)(5);
  CNStageIntLLRInputS4xD(40)(5) <= VNStageIntLLROutputS3xD(334)(0);
  CNStageIntLLRInputS4xD(66)(5) <= VNStageIntLLROutputS3xD(334)(1);
  CNStageIntLLRInputS4xD(217)(5) <= VNStageIntLLROutputS3xD(334)(2);
  CNStageIntLLRInputS4xD(286)(5) <= VNStageIntLLROutputS3xD(334)(3);
  CNStageIntLLRInputS4xD(380)(5) <= VNStageIntLLROutputS3xD(334)(4);
  CNStageIntLLRInputS4xD(39)(5) <= VNStageIntLLROutputS3xD(335)(0);
  CNStageIntLLRInputS4xD(78)(5) <= VNStageIntLLROutputS3xD(335)(1);
  CNStageIntLLRInputS4xD(170)(5) <= VNStageIntLLROutputS3xD(335)(2);
  CNStageIntLLRInputS4xD(189)(5) <= VNStageIntLLROutputS3xD(335)(3);
  CNStageIntLLRInputS4xD(274)(5) <= VNStageIntLLROutputS3xD(335)(4);
  CNStageIntLLRInputS4xD(291)(5) <= VNStageIntLLROutputS3xD(335)(5);
  CNStageIntLLRInputS4xD(343)(5) <= VNStageIntLLROutputS3xD(335)(6);
  CNStageIntLLRInputS4xD(38)(5) <= VNStageIntLLROutputS3xD(336)(0);
  CNStageIntLLRInputS4xD(104)(5) <= VNStageIntLLROutputS3xD(336)(1);
  CNStageIntLLRInputS4xD(121)(5) <= VNStageIntLLROutputS3xD(336)(2);
  CNStageIntLLRInputS4xD(267)(5) <= VNStageIntLLROutputS3xD(336)(3);
  CNStageIntLLRInputS4xD(332)(5) <= VNStageIntLLROutputS3xD(336)(4);
  CNStageIntLLRInputS4xD(344)(5) <= VNStageIntLLROutputS3xD(336)(5);
  CNStageIntLLRInputS4xD(37)(5) <= VNStageIntLLROutputS3xD(337)(0);
  CNStageIntLLRInputS4xD(93)(5) <= VNStageIntLLROutputS3xD(337)(1);
  CNStageIntLLRInputS4xD(115)(5) <= VNStageIntLLROutputS3xD(337)(2);
  CNStageIntLLRInputS4xD(183)(5) <= VNStageIntLLROutputS3xD(337)(3);
  CNStageIntLLRInputS4xD(253)(5) <= VNStageIntLLROutputS3xD(337)(4);
  CNStageIntLLRInputS4xD(290)(5) <= VNStageIntLLROutputS3xD(337)(5);
  CNStageIntLLRInputS4xD(379)(5) <= VNStageIntLLROutputS3xD(337)(6);
  CNStageIntLLRInputS4xD(36)(5) <= VNStageIntLLROutputS3xD(338)(0);
  CNStageIntLLRInputS4xD(80)(5) <= VNStageIntLLROutputS3xD(338)(1);
  CNStageIntLLRInputS4xD(155)(5) <= VNStageIntLLROutputS3xD(338)(2);
  CNStageIntLLRInputS4xD(190)(5) <= VNStageIntLLROutputS3xD(338)(3);
  CNStageIntLLRInputS4xD(370)(5) <= VNStageIntLLROutputS3xD(338)(4);
  CNStageIntLLRInputS4xD(35)(5) <= VNStageIntLLROutputS3xD(339)(0);
  CNStageIntLLRInputS4xD(96)(5) <= VNStageIntLLROutputS3xD(339)(1);
  CNStageIntLLRInputS4xD(163)(5) <= VNStageIntLLROutputS3xD(339)(2);
  CNStageIntLLRInputS4xD(216)(5) <= VNStageIntLLROutputS3xD(339)(3);
  CNStageIntLLRInputS4xD(247)(5) <= VNStageIntLLROutputS3xD(339)(4);
  CNStageIntLLRInputS4xD(322)(5) <= VNStageIntLLROutputS3xD(339)(5);
  CNStageIntLLRInputS4xD(34)(5) <= VNStageIntLLROutputS3xD(340)(0);
  CNStageIntLLRInputS4xD(58)(5) <= VNStageIntLLROutputS3xD(340)(1);
  CNStageIntLLRInputS4xD(127)(5) <= VNStageIntLLROutputS3xD(340)(2);
  CNStageIntLLRInputS4xD(178)(5) <= VNStageIntLLROutputS3xD(340)(3);
  CNStageIntLLRInputS4xD(245)(5) <= VNStageIntLLROutputS3xD(340)(4);
  CNStageIntLLRInputS4xD(334)(5) <= VNStageIntLLROutputS3xD(340)(5);
  CNStageIntLLRInputS4xD(33)(5) <= VNStageIntLLROutputS3xD(341)(0);
  CNStageIntLLRInputS4xD(68)(5) <= VNStageIntLLROutputS3xD(341)(1);
  CNStageIntLLRInputS4xD(125)(5) <= VNStageIntLLROutputS3xD(341)(2);
  CNStageIntLLRInputS4xD(204)(5) <= VNStageIntLLROutputS3xD(341)(3);
  CNStageIntLLRInputS4xD(258)(5) <= VNStageIntLLROutputS3xD(341)(4);
  CNStageIntLLRInputS4xD(296)(5) <= VNStageIntLLROutputS3xD(341)(5);
  CNStageIntLLRInputS4xD(32)(5) <= VNStageIntLLROutputS3xD(342)(0);
  CNStageIntLLRInputS4xD(63)(5) <= VNStageIntLLROutputS3xD(342)(1);
  CNStageIntLLRInputS4xD(161)(5) <= VNStageIntLLROutputS3xD(342)(2);
  CNStageIntLLRInputS4xD(251)(5) <= VNStageIntLLROutputS3xD(342)(3);
  CNStageIntLLRInputS4xD(294)(5) <= VNStageIntLLROutputS3xD(342)(4);
  CNStageIntLLRInputS4xD(31)(5) <= VNStageIntLLROutputS3xD(343)(0);
  CNStageIntLLRInputS4xD(69)(5) <= VNStageIntLLROutputS3xD(343)(1);
  CNStageIntLLRInputS4xD(140)(5) <= VNStageIntLLROutputS3xD(343)(2);
  CNStageIntLLRInputS4xD(206)(5) <= VNStageIntLLROutputS3xD(343)(3);
  CNStageIntLLRInputS4xD(228)(5) <= VNStageIntLLROutputS3xD(343)(4);
  CNStageIntLLRInputS4xD(327)(5) <= VNStageIntLLROutputS3xD(343)(5);
  CNStageIntLLRInputS4xD(30)(5) <= VNStageIntLLROutputS3xD(344)(0);
  CNStageIntLLRInputS4xD(57)(5) <= VNStageIntLLROutputS3xD(344)(1);
  CNStageIntLLRInputS4xD(143)(5) <= VNStageIntLLROutputS3xD(344)(2);
  CNStageIntLLRInputS4xD(218)(5) <= VNStageIntLLROutputS3xD(344)(3);
  CNStageIntLLRInputS4xD(238)(5) <= VNStageIntLLROutputS3xD(344)(4);
  CNStageIntLLRInputS4xD(307)(5) <= VNStageIntLLROutputS3xD(344)(5);
  CNStageIntLLRInputS4xD(367)(5) <= VNStageIntLLROutputS3xD(344)(6);
  CNStageIntLLRInputS4xD(29)(5) <= VNStageIntLLROutputS3xD(345)(0);
  CNStageIntLLRInputS4xD(83)(5) <= VNStageIntLLROutputS3xD(345)(1);
  CNStageIntLLRInputS4xD(128)(5) <= VNStageIntLLROutputS3xD(345)(2);
  CNStageIntLLRInputS4xD(232)(5) <= VNStageIntLLROutputS3xD(345)(3);
  CNStageIntLLRInputS4xD(309)(5) <= VNStageIntLLROutputS3xD(345)(4);
  CNStageIntLLRInputS4xD(375)(5) <= VNStageIntLLROutputS3xD(345)(5);
  CNStageIntLLRInputS4xD(28)(5) <= VNStageIntLLROutputS3xD(346)(0);
  CNStageIntLLRInputS4xD(89)(5) <= VNStageIntLLROutputS3xD(346)(1);
  CNStageIntLLRInputS4xD(162)(5) <= VNStageIntLLROutputS3xD(346)(2);
  CNStageIntLLRInputS4xD(181)(5) <= VNStageIntLLROutputS3xD(346)(3);
  CNStageIntLLRInputS4xD(235)(5) <= VNStageIntLLROutputS3xD(346)(4);
  CNStageIntLLRInputS4xD(297)(5) <= VNStageIntLLROutputS3xD(346)(5);
  CNStageIntLLRInputS4xD(339)(5) <= VNStageIntLLROutputS3xD(346)(6);
  CNStageIntLLRInputS4xD(27)(5) <= VNStageIntLLROutputS3xD(347)(0);
  CNStageIntLLRInputS4xD(73)(5) <= VNStageIntLLROutputS3xD(347)(1);
  CNStageIntLLRInputS4xD(124)(5) <= VNStageIntLLROutputS3xD(347)(2);
  CNStageIntLLRInputS4xD(199)(5) <= VNStageIntLLROutputS3xD(347)(3);
  CNStageIntLLRInputS4xD(225)(5) <= VNStageIntLLROutputS3xD(347)(4);
  CNStageIntLLRInputS4xD(328)(5) <= VNStageIntLLROutputS3xD(347)(5);
  CNStageIntLLRInputS4xD(337)(5) <= VNStageIntLLROutputS3xD(347)(6);
  CNStageIntLLRInputS4xD(26)(5) <= VNStageIntLLROutputS3xD(348)(0);
  CNStageIntLLRInputS4xD(75)(5) <= VNStageIntLLROutputS3xD(348)(1);
  CNStageIntLLRInputS4xD(152)(5) <= VNStageIntLLROutputS3xD(348)(2);
  CNStageIntLLRInputS4xD(200)(5) <= VNStageIntLLROutputS3xD(348)(3);
  CNStageIntLLRInputS4xD(259)(5) <= VNStageIntLLROutputS3xD(348)(4);
  CNStageIntLLRInputS4xD(293)(5) <= VNStageIntLLROutputS3xD(348)(5);
  CNStageIntLLRInputS4xD(373)(5) <= VNStageIntLLROutputS3xD(348)(6);
  CNStageIntLLRInputS4xD(25)(5) <= VNStageIntLLROutputS3xD(349)(0);
  CNStageIntLLRInputS4xD(99)(5) <= VNStageIntLLROutputS3xD(349)(1);
  CNStageIntLLRInputS4xD(180)(5) <= VNStageIntLLROutputS3xD(349)(2);
  CNStageIntLLRInputS4xD(244)(5) <= VNStageIntLLROutputS3xD(349)(3);
  CNStageIntLLRInputS4xD(319)(5) <= VNStageIntLLROutputS3xD(349)(4);
  CNStageIntLLRInputS4xD(352)(5) <= VNStageIntLLROutputS3xD(349)(5);
  CNStageIntLLRInputS4xD(24)(5) <= VNStageIntLLROutputS3xD(350)(0);
  CNStageIntLLRInputS4xD(81)(5) <= VNStageIntLLROutputS3xD(350)(1);
  CNStageIntLLRInputS4xD(164)(5) <= VNStageIntLLROutputS3xD(350)(2);
  CNStageIntLLRInputS4xD(171)(5) <= VNStageIntLLROutputS3xD(350)(3);
  CNStageIntLLRInputS4xD(254)(5) <= VNStageIntLLROutputS3xD(350)(4);
  CNStageIntLLRInputS4xD(303)(5) <= VNStageIntLLROutputS3xD(350)(5);
  CNStageIntLLRInputS4xD(23)(5) <= VNStageIntLLROutputS3xD(351)(0);
  CNStageIntLLRInputS4xD(154)(5) <= VNStageIntLLROutputS3xD(351)(1);
  CNStageIntLLRInputS4xD(188)(5) <= VNStageIntLLROutputS3xD(351)(2);
  CNStageIntLLRInputS4xD(266)(5) <= VNStageIntLLROutputS3xD(351)(3);
  CNStageIntLLRInputS4xD(329)(5) <= VNStageIntLLROutputS3xD(351)(4);
  CNStageIntLLRInputS4xD(340)(5) <= VNStageIntLLROutputS3xD(351)(5);
  CNStageIntLLRInputS4xD(22)(5) <= VNStageIntLLROutputS3xD(352)(0);
  CNStageIntLLRInputS4xD(100)(5) <= VNStageIntLLROutputS3xD(352)(1);
  CNStageIntLLRInputS4xD(141)(5) <= VNStageIntLLROutputS3xD(352)(2);
  CNStageIntLLRInputS4xD(192)(5) <= VNStageIntLLROutputS3xD(352)(3);
  CNStageIntLLRInputS4xD(239)(5) <= VNStageIntLLROutputS3xD(352)(4);
  CNStageIntLLRInputS4xD(321)(5) <= VNStageIntLLROutputS3xD(352)(5);
  CNStageIntLLRInputS4xD(374)(5) <= VNStageIntLLROutputS3xD(352)(6);
  CNStageIntLLRInputS4xD(21)(5) <= VNStageIntLLROutputS3xD(353)(0);
  CNStageIntLLRInputS4xD(74)(5) <= VNStageIntLLROutputS3xD(353)(1);
  CNStageIntLLRInputS4xD(160)(5) <= VNStageIntLLROutputS3xD(353)(2);
  CNStageIntLLRInputS4xD(224)(5) <= VNStageIntLLROutputS3xD(353)(3);
  CNStageIntLLRInputS4xD(227)(5) <= VNStageIntLLROutputS3xD(353)(4);
  CNStageIntLLRInputS4xD(336)(5) <= VNStageIntLLROutputS3xD(353)(5);
  CNStageIntLLRInputS4xD(20)(5) <= VNStageIntLLROutputS3xD(354)(0);
  CNStageIntLLRInputS4xD(88)(5) <= VNStageIntLLROutputS3xD(354)(1);
  CNStageIntLLRInputS4xD(133)(5) <= VNStageIntLLROutputS3xD(354)(2);
  CNStageIntLLRInputS4xD(191)(5) <= VNStageIntLLROutputS3xD(354)(3);
  CNStageIntLLRInputS4xD(326)(5) <= VNStageIntLLROutputS3xD(354)(4);
  CNStageIntLLRInputS4xD(364)(5) <= VNStageIntLLROutputS3xD(354)(5);
  CNStageIntLLRInputS4xD(19)(5) <= VNStageIntLLROutputS3xD(355)(0);
  CNStageIntLLRInputS4xD(59)(5) <= VNStageIntLLROutputS3xD(355)(1);
  CNStageIntLLRInputS4xD(130)(5) <= VNStageIntLLROutputS3xD(355)(2);
  CNStageIntLLRInputS4xD(186)(5) <= VNStageIntLLROutputS3xD(355)(3);
  CNStageIntLLRInputS4xD(230)(5) <= VNStageIntLLROutputS3xD(355)(4);
  CNStageIntLLRInputS4xD(300)(5) <= VNStageIntLLROutputS3xD(355)(5);
  CNStageIntLLRInputS4xD(349)(5) <= VNStageIntLLROutputS3xD(355)(6);
  CNStageIntLLRInputS4xD(18)(5) <= VNStageIntLLROutputS3xD(356)(0);
  CNStageIntLLRInputS4xD(95)(5) <= VNStageIntLLROutputS3xD(356)(1);
  CNStageIntLLRInputS4xD(146)(5) <= VNStageIntLLROutputS3xD(356)(2);
  CNStageIntLLRInputS4xD(222)(5) <= VNStageIntLLROutputS3xD(356)(3);
  CNStageIntLLRInputS4xD(299)(5) <= VNStageIntLLROutputS3xD(356)(4);
  CNStageIntLLRInputS4xD(376)(5) <= VNStageIntLLROutputS3xD(356)(5);
  CNStageIntLLRInputS4xD(17)(5) <= VNStageIntLLROutputS3xD(357)(0);
  CNStageIntLLRInputS4xD(61)(5) <= VNStageIntLLROutputS3xD(357)(1);
  CNStageIntLLRInputS4xD(138)(5) <= VNStageIntLLROutputS3xD(357)(2);
  CNStageIntLLRInputS4xD(176)(5) <= VNStageIntLLROutputS3xD(357)(3);
  CNStageIntLLRInputS4xD(256)(5) <= VNStageIntLLROutputS3xD(357)(4);
  CNStageIntLLRInputS4xD(312)(5) <= VNStageIntLLROutputS3xD(357)(5);
  CNStageIntLLRInputS4xD(366)(5) <= VNStageIntLLROutputS3xD(357)(6);
  CNStageIntLLRInputS4xD(16)(5) <= VNStageIntLLROutputS3xD(358)(0);
  CNStageIntLLRInputS4xD(76)(5) <= VNStageIntLLROutputS3xD(358)(1);
  CNStageIntLLRInputS4xD(112)(5) <= VNStageIntLLROutputS3xD(358)(2);
  CNStageIntLLRInputS4xD(252)(5) <= VNStageIntLLROutputS3xD(358)(3);
  CNStageIntLLRInputS4xD(305)(5) <= VNStageIntLLROutputS3xD(358)(4);
  CNStageIntLLRInputS4xD(353)(5) <= VNStageIntLLROutputS3xD(358)(5);
  CNStageIntLLRInputS4xD(15)(5) <= VNStageIntLLROutputS3xD(359)(0);
  CNStageIntLLRInputS4xD(72)(5) <= VNStageIntLLROutputS3xD(359)(1);
  CNStageIntLLRInputS4xD(122)(5) <= VNStageIntLLROutputS3xD(359)(2);
  CNStageIntLLRInputS4xD(195)(5) <= VNStageIntLLROutputS3xD(359)(3);
  CNStageIntLLRInputS4xD(257)(5) <= VNStageIntLLROutputS3xD(359)(4);
  CNStageIntLLRInputS4xD(283)(5) <= VNStageIntLLROutputS3xD(359)(5);
  CNStageIntLLRInputS4xD(372)(5) <= VNStageIntLLROutputS3xD(359)(6);
  CNStageIntLLRInputS4xD(14)(5) <= VNStageIntLLROutputS3xD(360)(0);
  CNStageIntLLRInputS4xD(91)(5) <= VNStageIntLLROutputS3xD(360)(1);
  CNStageIntLLRInputS4xD(116)(5) <= VNStageIntLLROutputS3xD(360)(2);
  CNStageIntLLRInputS4xD(174)(5) <= VNStageIntLLROutputS3xD(360)(3);
  CNStageIntLLRInputS4xD(248)(5) <= VNStageIntLLROutputS3xD(360)(4);
  CNStageIntLLRInputS4xD(292)(5) <= VNStageIntLLROutputS3xD(360)(5);
  CNStageIntLLRInputS4xD(345)(5) <= VNStageIntLLROutputS3xD(360)(6);
  CNStageIntLLRInputS4xD(13)(5) <= VNStageIntLLROutputS3xD(361)(0);
  CNStageIntLLRInputS4xD(54)(5) <= VNStageIntLLROutputS3xD(361)(1);
  CNStageIntLLRInputS4xD(120)(5) <= VNStageIntLLROutputS3xD(361)(2);
  CNStageIntLLRInputS4xD(207)(5) <= VNStageIntLLROutputS3xD(361)(3);
  CNStageIntLLRInputS4xD(271)(5) <= VNStageIntLLROutputS3xD(361)(4);
  CNStageIntLLRInputS4xD(285)(5) <= VNStageIntLLROutputS3xD(361)(5);
  CNStageIntLLRInputS4xD(342)(5) <= VNStageIntLLROutputS3xD(361)(6);
  CNStageIntLLRInputS4xD(12)(5) <= VNStageIntLLROutputS3xD(362)(0);
  CNStageIntLLRInputS4xD(55)(5) <= VNStageIntLLROutputS3xD(362)(1);
  CNStageIntLLRInputS4xD(169)(5) <= VNStageIntLLROutputS3xD(362)(2);
  CNStageIntLLRInputS4xD(210)(5) <= VNStageIntLLROutputS3xD(362)(3);
  CNStageIntLLRInputS4xD(276)(5) <= VNStageIntLLROutputS3xD(362)(4);
  CNStageIntLLRInputS4xD(289)(5) <= VNStageIntLLROutputS3xD(362)(5);
  CNStageIntLLRInputS4xD(357)(5) <= VNStageIntLLROutputS3xD(362)(6);
  CNStageIntLLRInputS4xD(90)(5) <= VNStageIntLLROutputS3xD(363)(0);
  CNStageIntLLRInputS4xD(147)(5) <= VNStageIntLLROutputS3xD(363)(1);
  CNStageIntLLRInputS4xD(197)(5) <= VNStageIntLLROutputS3xD(363)(2);
  CNStageIntLLRInputS4xD(261)(5) <= VNStageIntLLROutputS3xD(363)(3);
  CNStageIntLLRInputS4xD(281)(5) <= VNStageIntLLROutputS3xD(363)(4);
  CNStageIntLLRInputS4xD(11)(5) <= VNStageIntLLROutputS3xD(364)(0);
  CNStageIntLLRInputS4xD(82)(5) <= VNStageIntLLROutputS3xD(364)(1);
  CNStageIntLLRInputS4xD(129)(5) <= VNStageIntLLROutputS3xD(364)(2);
  CNStageIntLLRInputS4xD(175)(5) <= VNStageIntLLROutputS3xD(364)(3);
  CNStageIntLLRInputS4xD(263)(5) <= VNStageIntLLROutputS3xD(364)(4);
  CNStageIntLLRInputS4xD(313)(5) <= VNStageIntLLROutputS3xD(364)(5);
  CNStageIntLLRInputS4xD(10)(5) <= VNStageIntLLROutputS3xD(365)(0);
  CNStageIntLLRInputS4xD(98)(5) <= VNStageIntLLROutputS3xD(365)(1);
  CNStageIntLLRInputS4xD(142)(5) <= VNStageIntLLROutputS3xD(365)(2);
  CNStageIntLLRInputS4xD(194)(5) <= VNStageIntLLROutputS3xD(365)(3);
  CNStageIntLLRInputS4xD(234)(5) <= VNStageIntLLROutputS3xD(365)(4);
  CNStageIntLLRInputS4xD(298)(5) <= VNStageIntLLROutputS3xD(365)(5);
  CNStageIntLLRInputS4xD(9)(5) <= VNStageIntLLROutputS3xD(366)(0);
  CNStageIntLLRInputS4xD(102)(5) <= VNStageIntLLROutputS3xD(366)(1);
  CNStageIntLLRInputS4xD(153)(5) <= VNStageIntLLROutputS3xD(366)(2);
  CNStageIntLLRInputS4xD(219)(5) <= VNStageIntLLROutputS3xD(366)(3);
  CNStageIntLLRInputS4xD(269)(5) <= VNStageIntLLROutputS3xD(366)(4);
  CNStageIntLLRInputS4xD(308)(5) <= VNStageIntLLROutputS3xD(366)(5);
  CNStageIntLLRInputS4xD(8)(5) <= VNStageIntLLROutputS3xD(367)(0);
  CNStageIntLLRInputS4xD(110)(5) <= VNStageIntLLROutputS3xD(367)(1);
  CNStageIntLLRInputS4xD(123)(5) <= VNStageIntLLROutputS3xD(367)(2);
  CNStageIntLLRInputS4xD(205)(5) <= VNStageIntLLROutputS3xD(367)(3);
  CNStageIntLLRInputS4xD(226)(5) <= VNStageIntLLROutputS3xD(367)(4);
  CNStageIntLLRInputS4xD(320)(5) <= VNStageIntLLROutputS3xD(367)(5);
  CNStageIntLLRInputS4xD(333)(5) <= VNStageIntLLROutputS3xD(367)(6);
  CNStageIntLLRInputS4xD(7)(5) <= VNStageIntLLROutputS3xD(368)(0);
  CNStageIntLLRInputS4xD(177)(5) <= VNStageIntLLROutputS3xD(368)(1);
  CNStageIntLLRInputS4xD(381)(5) <= VNStageIntLLROutputS3xD(368)(2);
  CNStageIntLLRInputS4xD(6)(5) <= VNStageIntLLROutputS3xD(369)(0);
  CNStageIntLLRInputS4xD(156)(5) <= VNStageIntLLROutputS3xD(369)(1);
  CNStageIntLLRInputS4xD(221)(5) <= VNStageIntLLROutputS3xD(369)(2);
  CNStageIntLLRInputS4xD(262)(5) <= VNStageIntLLROutputS3xD(369)(3);
  CNStageIntLLRInputS4xD(358)(5) <= VNStageIntLLROutputS3xD(369)(4);
  CNStageIntLLRInputS4xD(5)(5) <= VNStageIntLLROutputS3xD(370)(0);
  CNStageIntLLRInputS4xD(114)(5) <= VNStageIntLLROutputS3xD(370)(1);
  CNStageIntLLRInputS4xD(208)(5) <= VNStageIntLLROutputS3xD(370)(2);
  CNStageIntLLRInputS4xD(275)(5) <= VNStageIntLLROutputS3xD(370)(3);
  CNStageIntLLRInputS4xD(341)(5) <= VNStageIntLLROutputS3xD(370)(4);
  CNStageIntLLRInputS4xD(4)(5) <= VNStageIntLLROutputS3xD(371)(0);
  CNStageIntLLRInputS4xD(135)(5) <= VNStageIntLLROutputS3xD(371)(1);
  CNStageIntLLRInputS4xD(173)(5) <= VNStageIntLLROutputS3xD(371)(2);
  CNStageIntLLRInputS4xD(249)(5) <= VNStageIntLLROutputS3xD(371)(3);
  CNStageIntLLRInputS4xD(354)(5) <= VNStageIntLLROutputS3xD(371)(4);
  CNStageIntLLRInputS4xD(106)(5) <= VNStageIntLLROutputS3xD(372)(0);
  CNStageIntLLRInputS4xD(144)(5) <= VNStageIntLLROutputS3xD(372)(1);
  CNStageIntLLRInputS4xD(201)(5) <= VNStageIntLLROutputS3xD(372)(2);
  CNStageIntLLRInputS4xD(229)(5) <= VNStageIntLLROutputS3xD(372)(3);
  CNStageIntLLRInputS4xD(301)(5) <= VNStageIntLLROutputS3xD(372)(4);
  CNStageIntLLRInputS4xD(365)(5) <= VNStageIntLLROutputS3xD(372)(5);
  CNStageIntLLRInputS4xD(3)(5) <= VNStageIntLLROutputS3xD(373)(0);
  CNStageIntLLRInputS4xD(139)(5) <= VNStageIntLLROutputS3xD(373)(1);
  CNStageIntLLRInputS4xD(250)(5) <= VNStageIntLLROutputS3xD(373)(2);
  CNStageIntLLRInputS4xD(310)(5) <= VNStageIntLLROutputS3xD(373)(3);
  CNStageIntLLRInputS4xD(335)(5) <= VNStageIntLLROutputS3xD(373)(4);
  CNStageIntLLRInputS4xD(2)(5) <= VNStageIntLLROutputS3xD(374)(0);
  CNStageIntLLRInputS4xD(85)(5) <= VNStageIntLLROutputS3xD(374)(1);
  CNStageIntLLRInputS4xD(145)(5) <= VNStageIntLLROutputS3xD(374)(2);
  CNStageIntLLRInputS4xD(213)(5) <= VNStageIntLLROutputS3xD(374)(3);
  CNStageIntLLRInputS4xD(264)(5) <= VNStageIntLLROutputS3xD(374)(4);
  CNStageIntLLRInputS4xD(306)(5) <= VNStageIntLLROutputS3xD(374)(5);
  CNStageIntLLRInputS4xD(383)(5) <= VNStageIntLLROutputS3xD(374)(6);
  CNStageIntLLRInputS4xD(1)(5) <= VNStageIntLLROutputS3xD(375)(0);
  CNStageIntLLRInputS4xD(64)(5) <= VNStageIntLLROutputS3xD(375)(1);
  CNStageIntLLRInputS4xD(134)(5) <= VNStageIntLLROutputS3xD(375)(2);
  CNStageIntLLRInputS4xD(260)(5) <= VNStageIntLLROutputS3xD(375)(3);
  CNStageIntLLRInputS4xD(311)(5) <= VNStageIntLLROutputS3xD(375)(4);
  CNStageIntLLRInputS4xD(368)(5) <= VNStageIntLLROutputS3xD(375)(5);
  CNStageIntLLRInputS4xD(0)(5) <= VNStageIntLLROutputS3xD(376)(0);
  CNStageIntLLRInputS4xD(67)(5) <= VNStageIntLLROutputS3xD(376)(1);
  CNStageIntLLRInputS4xD(159)(5) <= VNStageIntLLROutputS3xD(376)(2);
  CNStageIntLLRInputS4xD(278)(5) <= VNStageIntLLROutputS3xD(376)(3);
  CNStageIntLLRInputS4xD(107)(5) <= VNStageIntLLROutputS3xD(377)(0);
  CNStageIntLLRInputS4xD(166)(5) <= VNStageIntLLROutputS3xD(377)(1);
  CNStageIntLLRInputS4xD(193)(5) <= VNStageIntLLROutputS3xD(377)(2);
  CNStageIntLLRInputS4xD(325)(5) <= VNStageIntLLROutputS3xD(377)(3);
  CNStageIntLLRInputS4xD(347)(5) <= VNStageIntLLROutputS3xD(377)(4);
  CNStageIntLLRInputS4xD(86)(5) <= VNStageIntLLROutputS3xD(378)(0);
  CNStageIntLLRInputS4xD(149)(5) <= VNStageIntLLROutputS3xD(378)(1);
  CNStageIntLLRInputS4xD(187)(5) <= VNStageIntLLROutputS3xD(378)(2);
  CNStageIntLLRInputS4xD(246)(5) <= VNStageIntLLROutputS3xD(378)(3);
  CNStageIntLLRInputS4xD(331)(5) <= VNStageIntLLROutputS3xD(378)(4);
  CNStageIntLLRInputS4xD(355)(5) <= VNStageIntLLROutputS3xD(378)(5);
  CNStageIntLLRInputS4xD(105)(5) <= VNStageIntLLROutputS3xD(379)(0);
  CNStageIntLLRInputS4xD(151)(5) <= VNStageIntLLROutputS3xD(379)(1);
  CNStageIntLLRInputS4xD(277)(5) <= VNStageIntLLROutputS3xD(379)(2);
  CNStageIntLLRInputS4xD(315)(5) <= VNStageIntLLROutputS3xD(379)(3);
  CNStageIntLLRInputS4xD(351)(5) <= VNStageIntLLROutputS3xD(379)(4);
  CNStageIntLLRInputS4xD(77)(5) <= VNStageIntLLROutputS3xD(380)(0);
  CNStageIntLLRInputS4xD(118)(5) <= VNStageIntLLROutputS3xD(380)(1);
  CNStageIntLLRInputS4xD(182)(5) <= VNStageIntLLROutputS3xD(380)(2);
  CNStageIntLLRInputS4xD(270)(5) <= VNStageIntLLROutputS3xD(380)(3);
  CNStageIntLLRInputS4xD(317)(5) <= VNStageIntLLROutputS3xD(380)(4);
  CNStageIntLLRInputS4xD(356)(5) <= VNStageIntLLROutputS3xD(380)(5);
  CNStageIntLLRInputS4xD(60)(5) <= VNStageIntLLROutputS3xD(381)(0);
  CNStageIntLLRInputS4xD(157)(5) <= VNStageIntLLROutputS3xD(381)(1);
  CNStageIntLLRInputS4xD(214)(5) <= VNStageIntLLROutputS3xD(381)(2);
  CNStageIntLLRInputS4xD(233)(5) <= VNStageIntLLROutputS3xD(381)(3);
  CNStageIntLLRInputS4xD(287)(5) <= VNStageIntLLROutputS3xD(381)(4);
  CNStageIntLLRInputS4xD(346)(5) <= VNStageIntLLROutputS3xD(381)(5);
  CNStageIntLLRInputS4xD(87)(5) <= VNStageIntLLROutputS3xD(382)(0);
  CNStageIntLLRInputS4xD(111)(5) <= VNStageIntLLROutputS3xD(382)(1);
  CNStageIntLLRInputS4xD(198)(5) <= VNStageIntLLROutputS3xD(382)(2);
  CNStageIntLLRInputS4xD(237)(5) <= VNStageIntLLROutputS3xD(382)(3);
  CNStageIntLLRInputS4xD(323)(5) <= VNStageIntLLROutputS3xD(382)(4);
  CNStageIntLLRInputS4xD(371)(5) <= VNStageIntLLROutputS3xD(382)(5);
  CNStageIntLLRInputS4xD(52)(5) <= VNStageIntLLROutputS3xD(383)(0);
  CNStageIntLLRInputS4xD(79)(5) <= VNStageIntLLROutputS3xD(383)(1);
  CNStageIntLLRInputS4xD(119)(5) <= VNStageIntLLROutputS3xD(383)(2);
  CNStageIntLLRInputS4xD(209)(5) <= VNStageIntLLROutputS3xD(383)(3);
  CNStageIntLLRInputS4xD(279)(5) <= VNStageIntLLROutputS3xD(383)(4);
  CNStageIntLLRInputS4xD(282)(5) <= VNStageIntLLROutputS3xD(383)(5);
  CNStageIntLLRInputS4xD(378)(5) <= VNStageIntLLROutputS3xD(383)(6);

  -- Variable Nodes (Iteration 4)
  VNStageIntLLRInputS4xD(56)(0) <= CNStageIntLLROutputS4xD(0)(0);
  VNStageIntLLRInputS4xD(120)(0) <= CNStageIntLLROutputS4xD(0)(1);
  VNStageIntLLRInputS4xD(184)(0) <= CNStageIntLLROutputS4xD(0)(2);
  VNStageIntLLRInputS4xD(248)(0) <= CNStageIntLLROutputS4xD(0)(3);
  VNStageIntLLRInputS4xD(312)(0) <= CNStageIntLLROutputS4xD(0)(4);
  VNStageIntLLRInputS4xD(376)(0) <= CNStageIntLLROutputS4xD(0)(5);
  VNStageIntLLRInputS4xD(55)(0) <= CNStageIntLLROutputS4xD(1)(0);
  VNStageIntLLRInputS4xD(119)(0) <= CNStageIntLLROutputS4xD(1)(1);
  VNStageIntLLRInputS4xD(183)(0) <= CNStageIntLLROutputS4xD(1)(2);
  VNStageIntLLRInputS4xD(247)(0) <= CNStageIntLLROutputS4xD(1)(3);
  VNStageIntLLRInputS4xD(311)(0) <= CNStageIntLLROutputS4xD(1)(4);
  VNStageIntLLRInputS4xD(375)(0) <= CNStageIntLLROutputS4xD(1)(5);
  VNStageIntLLRInputS4xD(54)(0) <= CNStageIntLLROutputS4xD(2)(0);
  VNStageIntLLRInputS4xD(118)(0) <= CNStageIntLLROutputS4xD(2)(1);
  VNStageIntLLRInputS4xD(182)(0) <= CNStageIntLLROutputS4xD(2)(2);
  VNStageIntLLRInputS4xD(246)(0) <= CNStageIntLLROutputS4xD(2)(3);
  VNStageIntLLRInputS4xD(310)(0) <= CNStageIntLLROutputS4xD(2)(4);
  VNStageIntLLRInputS4xD(374)(0) <= CNStageIntLLROutputS4xD(2)(5);
  VNStageIntLLRInputS4xD(53)(0) <= CNStageIntLLROutputS4xD(3)(0);
  VNStageIntLLRInputS4xD(117)(0) <= CNStageIntLLROutputS4xD(3)(1);
  VNStageIntLLRInputS4xD(181)(0) <= CNStageIntLLROutputS4xD(3)(2);
  VNStageIntLLRInputS4xD(245)(0) <= CNStageIntLLROutputS4xD(3)(3);
  VNStageIntLLRInputS4xD(309)(0) <= CNStageIntLLROutputS4xD(3)(4);
  VNStageIntLLRInputS4xD(373)(0) <= CNStageIntLLROutputS4xD(3)(5);
  VNStageIntLLRInputS4xD(51)(0) <= CNStageIntLLROutputS4xD(4)(0);
  VNStageIntLLRInputS4xD(115)(0) <= CNStageIntLLROutputS4xD(4)(1);
  VNStageIntLLRInputS4xD(179)(0) <= CNStageIntLLROutputS4xD(4)(2);
  VNStageIntLLRInputS4xD(243)(0) <= CNStageIntLLROutputS4xD(4)(3);
  VNStageIntLLRInputS4xD(307)(0) <= CNStageIntLLROutputS4xD(4)(4);
  VNStageIntLLRInputS4xD(371)(0) <= CNStageIntLLROutputS4xD(4)(5);
  VNStageIntLLRInputS4xD(50)(0) <= CNStageIntLLROutputS4xD(5)(0);
  VNStageIntLLRInputS4xD(114)(0) <= CNStageIntLLROutputS4xD(5)(1);
  VNStageIntLLRInputS4xD(178)(0) <= CNStageIntLLROutputS4xD(5)(2);
  VNStageIntLLRInputS4xD(242)(0) <= CNStageIntLLROutputS4xD(5)(3);
  VNStageIntLLRInputS4xD(306)(0) <= CNStageIntLLROutputS4xD(5)(4);
  VNStageIntLLRInputS4xD(370)(0) <= CNStageIntLLROutputS4xD(5)(5);
  VNStageIntLLRInputS4xD(49)(0) <= CNStageIntLLROutputS4xD(6)(0);
  VNStageIntLLRInputS4xD(113)(0) <= CNStageIntLLROutputS4xD(6)(1);
  VNStageIntLLRInputS4xD(177)(0) <= CNStageIntLLROutputS4xD(6)(2);
  VNStageIntLLRInputS4xD(241)(0) <= CNStageIntLLROutputS4xD(6)(3);
  VNStageIntLLRInputS4xD(305)(0) <= CNStageIntLLROutputS4xD(6)(4);
  VNStageIntLLRInputS4xD(369)(0) <= CNStageIntLLROutputS4xD(6)(5);
  VNStageIntLLRInputS4xD(48)(0) <= CNStageIntLLROutputS4xD(7)(0);
  VNStageIntLLRInputS4xD(112)(0) <= CNStageIntLLROutputS4xD(7)(1);
  VNStageIntLLRInputS4xD(176)(0) <= CNStageIntLLROutputS4xD(7)(2);
  VNStageIntLLRInputS4xD(240)(0) <= CNStageIntLLROutputS4xD(7)(3);
  VNStageIntLLRInputS4xD(304)(0) <= CNStageIntLLROutputS4xD(7)(4);
  VNStageIntLLRInputS4xD(368)(0) <= CNStageIntLLROutputS4xD(7)(5);
  VNStageIntLLRInputS4xD(47)(0) <= CNStageIntLLROutputS4xD(8)(0);
  VNStageIntLLRInputS4xD(111)(0) <= CNStageIntLLROutputS4xD(8)(1);
  VNStageIntLLRInputS4xD(175)(0) <= CNStageIntLLROutputS4xD(8)(2);
  VNStageIntLLRInputS4xD(239)(0) <= CNStageIntLLROutputS4xD(8)(3);
  VNStageIntLLRInputS4xD(303)(0) <= CNStageIntLLROutputS4xD(8)(4);
  VNStageIntLLRInputS4xD(367)(0) <= CNStageIntLLROutputS4xD(8)(5);
  VNStageIntLLRInputS4xD(46)(0) <= CNStageIntLLROutputS4xD(9)(0);
  VNStageIntLLRInputS4xD(110)(0) <= CNStageIntLLROutputS4xD(9)(1);
  VNStageIntLLRInputS4xD(174)(0) <= CNStageIntLLROutputS4xD(9)(2);
  VNStageIntLLRInputS4xD(238)(0) <= CNStageIntLLROutputS4xD(9)(3);
  VNStageIntLLRInputS4xD(302)(0) <= CNStageIntLLROutputS4xD(9)(4);
  VNStageIntLLRInputS4xD(366)(0) <= CNStageIntLLROutputS4xD(9)(5);
  VNStageIntLLRInputS4xD(45)(0) <= CNStageIntLLROutputS4xD(10)(0);
  VNStageIntLLRInputS4xD(109)(0) <= CNStageIntLLROutputS4xD(10)(1);
  VNStageIntLLRInputS4xD(173)(0) <= CNStageIntLLROutputS4xD(10)(2);
  VNStageIntLLRInputS4xD(237)(0) <= CNStageIntLLROutputS4xD(10)(3);
  VNStageIntLLRInputS4xD(301)(0) <= CNStageIntLLROutputS4xD(10)(4);
  VNStageIntLLRInputS4xD(365)(0) <= CNStageIntLLROutputS4xD(10)(5);
  VNStageIntLLRInputS4xD(44)(0) <= CNStageIntLLROutputS4xD(11)(0);
  VNStageIntLLRInputS4xD(108)(0) <= CNStageIntLLROutputS4xD(11)(1);
  VNStageIntLLRInputS4xD(172)(0) <= CNStageIntLLROutputS4xD(11)(2);
  VNStageIntLLRInputS4xD(236)(0) <= CNStageIntLLROutputS4xD(11)(3);
  VNStageIntLLRInputS4xD(300)(0) <= CNStageIntLLROutputS4xD(11)(4);
  VNStageIntLLRInputS4xD(364)(0) <= CNStageIntLLROutputS4xD(11)(5);
  VNStageIntLLRInputS4xD(42)(0) <= CNStageIntLLROutputS4xD(12)(0);
  VNStageIntLLRInputS4xD(106)(0) <= CNStageIntLLROutputS4xD(12)(1);
  VNStageIntLLRInputS4xD(170)(0) <= CNStageIntLLROutputS4xD(12)(2);
  VNStageIntLLRInputS4xD(234)(0) <= CNStageIntLLROutputS4xD(12)(3);
  VNStageIntLLRInputS4xD(298)(0) <= CNStageIntLLROutputS4xD(12)(4);
  VNStageIntLLRInputS4xD(362)(0) <= CNStageIntLLROutputS4xD(12)(5);
  VNStageIntLLRInputS4xD(41)(0) <= CNStageIntLLROutputS4xD(13)(0);
  VNStageIntLLRInputS4xD(105)(0) <= CNStageIntLLROutputS4xD(13)(1);
  VNStageIntLLRInputS4xD(169)(0) <= CNStageIntLLROutputS4xD(13)(2);
  VNStageIntLLRInputS4xD(233)(0) <= CNStageIntLLROutputS4xD(13)(3);
  VNStageIntLLRInputS4xD(297)(0) <= CNStageIntLLROutputS4xD(13)(4);
  VNStageIntLLRInputS4xD(361)(0) <= CNStageIntLLROutputS4xD(13)(5);
  VNStageIntLLRInputS4xD(40)(0) <= CNStageIntLLROutputS4xD(14)(0);
  VNStageIntLLRInputS4xD(104)(0) <= CNStageIntLLROutputS4xD(14)(1);
  VNStageIntLLRInputS4xD(168)(0) <= CNStageIntLLROutputS4xD(14)(2);
  VNStageIntLLRInputS4xD(232)(0) <= CNStageIntLLROutputS4xD(14)(3);
  VNStageIntLLRInputS4xD(296)(0) <= CNStageIntLLROutputS4xD(14)(4);
  VNStageIntLLRInputS4xD(360)(0) <= CNStageIntLLROutputS4xD(14)(5);
  VNStageIntLLRInputS4xD(39)(0) <= CNStageIntLLROutputS4xD(15)(0);
  VNStageIntLLRInputS4xD(103)(0) <= CNStageIntLLROutputS4xD(15)(1);
  VNStageIntLLRInputS4xD(167)(0) <= CNStageIntLLROutputS4xD(15)(2);
  VNStageIntLLRInputS4xD(231)(0) <= CNStageIntLLROutputS4xD(15)(3);
  VNStageIntLLRInputS4xD(295)(0) <= CNStageIntLLROutputS4xD(15)(4);
  VNStageIntLLRInputS4xD(359)(0) <= CNStageIntLLROutputS4xD(15)(5);
  VNStageIntLLRInputS4xD(38)(0) <= CNStageIntLLROutputS4xD(16)(0);
  VNStageIntLLRInputS4xD(102)(0) <= CNStageIntLLROutputS4xD(16)(1);
  VNStageIntLLRInputS4xD(166)(0) <= CNStageIntLLROutputS4xD(16)(2);
  VNStageIntLLRInputS4xD(230)(0) <= CNStageIntLLROutputS4xD(16)(3);
  VNStageIntLLRInputS4xD(294)(0) <= CNStageIntLLROutputS4xD(16)(4);
  VNStageIntLLRInputS4xD(358)(0) <= CNStageIntLLROutputS4xD(16)(5);
  VNStageIntLLRInputS4xD(37)(0) <= CNStageIntLLROutputS4xD(17)(0);
  VNStageIntLLRInputS4xD(101)(0) <= CNStageIntLLROutputS4xD(17)(1);
  VNStageIntLLRInputS4xD(165)(0) <= CNStageIntLLROutputS4xD(17)(2);
  VNStageIntLLRInputS4xD(229)(0) <= CNStageIntLLROutputS4xD(17)(3);
  VNStageIntLLRInputS4xD(293)(0) <= CNStageIntLLROutputS4xD(17)(4);
  VNStageIntLLRInputS4xD(357)(0) <= CNStageIntLLROutputS4xD(17)(5);
  VNStageIntLLRInputS4xD(36)(0) <= CNStageIntLLROutputS4xD(18)(0);
  VNStageIntLLRInputS4xD(100)(0) <= CNStageIntLLROutputS4xD(18)(1);
  VNStageIntLLRInputS4xD(164)(0) <= CNStageIntLLROutputS4xD(18)(2);
  VNStageIntLLRInputS4xD(228)(0) <= CNStageIntLLROutputS4xD(18)(3);
  VNStageIntLLRInputS4xD(292)(0) <= CNStageIntLLROutputS4xD(18)(4);
  VNStageIntLLRInputS4xD(356)(0) <= CNStageIntLLROutputS4xD(18)(5);
  VNStageIntLLRInputS4xD(35)(0) <= CNStageIntLLROutputS4xD(19)(0);
  VNStageIntLLRInputS4xD(99)(0) <= CNStageIntLLROutputS4xD(19)(1);
  VNStageIntLLRInputS4xD(163)(0) <= CNStageIntLLROutputS4xD(19)(2);
  VNStageIntLLRInputS4xD(227)(0) <= CNStageIntLLROutputS4xD(19)(3);
  VNStageIntLLRInputS4xD(291)(0) <= CNStageIntLLROutputS4xD(19)(4);
  VNStageIntLLRInputS4xD(355)(0) <= CNStageIntLLROutputS4xD(19)(5);
  VNStageIntLLRInputS4xD(34)(0) <= CNStageIntLLROutputS4xD(20)(0);
  VNStageIntLLRInputS4xD(98)(0) <= CNStageIntLLROutputS4xD(20)(1);
  VNStageIntLLRInputS4xD(162)(0) <= CNStageIntLLROutputS4xD(20)(2);
  VNStageIntLLRInputS4xD(226)(0) <= CNStageIntLLROutputS4xD(20)(3);
  VNStageIntLLRInputS4xD(290)(0) <= CNStageIntLLROutputS4xD(20)(4);
  VNStageIntLLRInputS4xD(354)(0) <= CNStageIntLLROutputS4xD(20)(5);
  VNStageIntLLRInputS4xD(33)(0) <= CNStageIntLLROutputS4xD(21)(0);
  VNStageIntLLRInputS4xD(97)(0) <= CNStageIntLLROutputS4xD(21)(1);
  VNStageIntLLRInputS4xD(161)(0) <= CNStageIntLLROutputS4xD(21)(2);
  VNStageIntLLRInputS4xD(225)(0) <= CNStageIntLLROutputS4xD(21)(3);
  VNStageIntLLRInputS4xD(289)(0) <= CNStageIntLLROutputS4xD(21)(4);
  VNStageIntLLRInputS4xD(353)(0) <= CNStageIntLLROutputS4xD(21)(5);
  VNStageIntLLRInputS4xD(32)(0) <= CNStageIntLLROutputS4xD(22)(0);
  VNStageIntLLRInputS4xD(96)(0) <= CNStageIntLLROutputS4xD(22)(1);
  VNStageIntLLRInputS4xD(160)(0) <= CNStageIntLLROutputS4xD(22)(2);
  VNStageIntLLRInputS4xD(224)(0) <= CNStageIntLLROutputS4xD(22)(3);
  VNStageIntLLRInputS4xD(288)(0) <= CNStageIntLLROutputS4xD(22)(4);
  VNStageIntLLRInputS4xD(352)(0) <= CNStageIntLLROutputS4xD(22)(5);
  VNStageIntLLRInputS4xD(31)(0) <= CNStageIntLLROutputS4xD(23)(0);
  VNStageIntLLRInputS4xD(95)(0) <= CNStageIntLLROutputS4xD(23)(1);
  VNStageIntLLRInputS4xD(159)(0) <= CNStageIntLLROutputS4xD(23)(2);
  VNStageIntLLRInputS4xD(223)(0) <= CNStageIntLLROutputS4xD(23)(3);
  VNStageIntLLRInputS4xD(287)(0) <= CNStageIntLLROutputS4xD(23)(4);
  VNStageIntLLRInputS4xD(351)(0) <= CNStageIntLLROutputS4xD(23)(5);
  VNStageIntLLRInputS4xD(30)(0) <= CNStageIntLLROutputS4xD(24)(0);
  VNStageIntLLRInputS4xD(94)(0) <= CNStageIntLLROutputS4xD(24)(1);
  VNStageIntLLRInputS4xD(158)(0) <= CNStageIntLLROutputS4xD(24)(2);
  VNStageIntLLRInputS4xD(222)(0) <= CNStageIntLLROutputS4xD(24)(3);
  VNStageIntLLRInputS4xD(286)(0) <= CNStageIntLLROutputS4xD(24)(4);
  VNStageIntLLRInputS4xD(350)(0) <= CNStageIntLLROutputS4xD(24)(5);
  VNStageIntLLRInputS4xD(29)(0) <= CNStageIntLLROutputS4xD(25)(0);
  VNStageIntLLRInputS4xD(93)(0) <= CNStageIntLLROutputS4xD(25)(1);
  VNStageIntLLRInputS4xD(157)(0) <= CNStageIntLLROutputS4xD(25)(2);
  VNStageIntLLRInputS4xD(221)(0) <= CNStageIntLLROutputS4xD(25)(3);
  VNStageIntLLRInputS4xD(285)(0) <= CNStageIntLLROutputS4xD(25)(4);
  VNStageIntLLRInputS4xD(349)(0) <= CNStageIntLLROutputS4xD(25)(5);
  VNStageIntLLRInputS4xD(28)(0) <= CNStageIntLLROutputS4xD(26)(0);
  VNStageIntLLRInputS4xD(92)(0) <= CNStageIntLLROutputS4xD(26)(1);
  VNStageIntLLRInputS4xD(156)(0) <= CNStageIntLLROutputS4xD(26)(2);
  VNStageIntLLRInputS4xD(220)(0) <= CNStageIntLLROutputS4xD(26)(3);
  VNStageIntLLRInputS4xD(284)(0) <= CNStageIntLLROutputS4xD(26)(4);
  VNStageIntLLRInputS4xD(348)(0) <= CNStageIntLLROutputS4xD(26)(5);
  VNStageIntLLRInputS4xD(27)(0) <= CNStageIntLLROutputS4xD(27)(0);
  VNStageIntLLRInputS4xD(91)(0) <= CNStageIntLLROutputS4xD(27)(1);
  VNStageIntLLRInputS4xD(155)(0) <= CNStageIntLLROutputS4xD(27)(2);
  VNStageIntLLRInputS4xD(219)(0) <= CNStageIntLLROutputS4xD(27)(3);
  VNStageIntLLRInputS4xD(283)(0) <= CNStageIntLLROutputS4xD(27)(4);
  VNStageIntLLRInputS4xD(347)(0) <= CNStageIntLLROutputS4xD(27)(5);
  VNStageIntLLRInputS4xD(26)(0) <= CNStageIntLLROutputS4xD(28)(0);
  VNStageIntLLRInputS4xD(90)(0) <= CNStageIntLLROutputS4xD(28)(1);
  VNStageIntLLRInputS4xD(154)(0) <= CNStageIntLLROutputS4xD(28)(2);
  VNStageIntLLRInputS4xD(218)(0) <= CNStageIntLLROutputS4xD(28)(3);
  VNStageIntLLRInputS4xD(282)(0) <= CNStageIntLLROutputS4xD(28)(4);
  VNStageIntLLRInputS4xD(346)(0) <= CNStageIntLLROutputS4xD(28)(5);
  VNStageIntLLRInputS4xD(25)(0) <= CNStageIntLLROutputS4xD(29)(0);
  VNStageIntLLRInputS4xD(89)(0) <= CNStageIntLLROutputS4xD(29)(1);
  VNStageIntLLRInputS4xD(153)(0) <= CNStageIntLLROutputS4xD(29)(2);
  VNStageIntLLRInputS4xD(217)(0) <= CNStageIntLLROutputS4xD(29)(3);
  VNStageIntLLRInputS4xD(281)(0) <= CNStageIntLLROutputS4xD(29)(4);
  VNStageIntLLRInputS4xD(345)(0) <= CNStageIntLLROutputS4xD(29)(5);
  VNStageIntLLRInputS4xD(24)(0) <= CNStageIntLLROutputS4xD(30)(0);
  VNStageIntLLRInputS4xD(88)(0) <= CNStageIntLLROutputS4xD(30)(1);
  VNStageIntLLRInputS4xD(152)(0) <= CNStageIntLLROutputS4xD(30)(2);
  VNStageIntLLRInputS4xD(216)(0) <= CNStageIntLLROutputS4xD(30)(3);
  VNStageIntLLRInputS4xD(280)(0) <= CNStageIntLLROutputS4xD(30)(4);
  VNStageIntLLRInputS4xD(344)(0) <= CNStageIntLLROutputS4xD(30)(5);
  VNStageIntLLRInputS4xD(23)(0) <= CNStageIntLLROutputS4xD(31)(0);
  VNStageIntLLRInputS4xD(87)(0) <= CNStageIntLLROutputS4xD(31)(1);
  VNStageIntLLRInputS4xD(151)(0) <= CNStageIntLLROutputS4xD(31)(2);
  VNStageIntLLRInputS4xD(215)(0) <= CNStageIntLLROutputS4xD(31)(3);
  VNStageIntLLRInputS4xD(279)(0) <= CNStageIntLLROutputS4xD(31)(4);
  VNStageIntLLRInputS4xD(343)(0) <= CNStageIntLLROutputS4xD(31)(5);
  VNStageIntLLRInputS4xD(22)(0) <= CNStageIntLLROutputS4xD(32)(0);
  VNStageIntLLRInputS4xD(86)(0) <= CNStageIntLLROutputS4xD(32)(1);
  VNStageIntLLRInputS4xD(150)(0) <= CNStageIntLLROutputS4xD(32)(2);
  VNStageIntLLRInputS4xD(214)(0) <= CNStageIntLLROutputS4xD(32)(3);
  VNStageIntLLRInputS4xD(278)(0) <= CNStageIntLLROutputS4xD(32)(4);
  VNStageIntLLRInputS4xD(342)(0) <= CNStageIntLLROutputS4xD(32)(5);
  VNStageIntLLRInputS4xD(21)(0) <= CNStageIntLLROutputS4xD(33)(0);
  VNStageIntLLRInputS4xD(85)(0) <= CNStageIntLLROutputS4xD(33)(1);
  VNStageIntLLRInputS4xD(149)(0) <= CNStageIntLLROutputS4xD(33)(2);
  VNStageIntLLRInputS4xD(213)(0) <= CNStageIntLLROutputS4xD(33)(3);
  VNStageIntLLRInputS4xD(277)(0) <= CNStageIntLLROutputS4xD(33)(4);
  VNStageIntLLRInputS4xD(341)(0) <= CNStageIntLLROutputS4xD(33)(5);
  VNStageIntLLRInputS4xD(20)(0) <= CNStageIntLLROutputS4xD(34)(0);
  VNStageIntLLRInputS4xD(84)(0) <= CNStageIntLLROutputS4xD(34)(1);
  VNStageIntLLRInputS4xD(148)(0) <= CNStageIntLLROutputS4xD(34)(2);
  VNStageIntLLRInputS4xD(212)(0) <= CNStageIntLLROutputS4xD(34)(3);
  VNStageIntLLRInputS4xD(276)(0) <= CNStageIntLLROutputS4xD(34)(4);
  VNStageIntLLRInputS4xD(340)(0) <= CNStageIntLLROutputS4xD(34)(5);
  VNStageIntLLRInputS4xD(19)(0) <= CNStageIntLLROutputS4xD(35)(0);
  VNStageIntLLRInputS4xD(83)(0) <= CNStageIntLLROutputS4xD(35)(1);
  VNStageIntLLRInputS4xD(147)(0) <= CNStageIntLLROutputS4xD(35)(2);
  VNStageIntLLRInputS4xD(211)(0) <= CNStageIntLLROutputS4xD(35)(3);
  VNStageIntLLRInputS4xD(275)(0) <= CNStageIntLLROutputS4xD(35)(4);
  VNStageIntLLRInputS4xD(339)(0) <= CNStageIntLLROutputS4xD(35)(5);
  VNStageIntLLRInputS4xD(18)(0) <= CNStageIntLLROutputS4xD(36)(0);
  VNStageIntLLRInputS4xD(82)(0) <= CNStageIntLLROutputS4xD(36)(1);
  VNStageIntLLRInputS4xD(146)(0) <= CNStageIntLLROutputS4xD(36)(2);
  VNStageIntLLRInputS4xD(210)(0) <= CNStageIntLLROutputS4xD(36)(3);
  VNStageIntLLRInputS4xD(274)(0) <= CNStageIntLLROutputS4xD(36)(4);
  VNStageIntLLRInputS4xD(338)(0) <= CNStageIntLLROutputS4xD(36)(5);
  VNStageIntLLRInputS4xD(17)(0) <= CNStageIntLLROutputS4xD(37)(0);
  VNStageIntLLRInputS4xD(81)(0) <= CNStageIntLLROutputS4xD(37)(1);
  VNStageIntLLRInputS4xD(145)(0) <= CNStageIntLLROutputS4xD(37)(2);
  VNStageIntLLRInputS4xD(209)(0) <= CNStageIntLLROutputS4xD(37)(3);
  VNStageIntLLRInputS4xD(273)(0) <= CNStageIntLLROutputS4xD(37)(4);
  VNStageIntLLRInputS4xD(337)(0) <= CNStageIntLLROutputS4xD(37)(5);
  VNStageIntLLRInputS4xD(16)(0) <= CNStageIntLLROutputS4xD(38)(0);
  VNStageIntLLRInputS4xD(80)(0) <= CNStageIntLLROutputS4xD(38)(1);
  VNStageIntLLRInputS4xD(144)(0) <= CNStageIntLLROutputS4xD(38)(2);
  VNStageIntLLRInputS4xD(208)(0) <= CNStageIntLLROutputS4xD(38)(3);
  VNStageIntLLRInputS4xD(272)(0) <= CNStageIntLLROutputS4xD(38)(4);
  VNStageIntLLRInputS4xD(336)(0) <= CNStageIntLLROutputS4xD(38)(5);
  VNStageIntLLRInputS4xD(15)(0) <= CNStageIntLLROutputS4xD(39)(0);
  VNStageIntLLRInputS4xD(79)(0) <= CNStageIntLLROutputS4xD(39)(1);
  VNStageIntLLRInputS4xD(143)(0) <= CNStageIntLLROutputS4xD(39)(2);
  VNStageIntLLRInputS4xD(207)(0) <= CNStageIntLLROutputS4xD(39)(3);
  VNStageIntLLRInputS4xD(271)(0) <= CNStageIntLLROutputS4xD(39)(4);
  VNStageIntLLRInputS4xD(335)(0) <= CNStageIntLLROutputS4xD(39)(5);
  VNStageIntLLRInputS4xD(14)(0) <= CNStageIntLLROutputS4xD(40)(0);
  VNStageIntLLRInputS4xD(78)(0) <= CNStageIntLLROutputS4xD(40)(1);
  VNStageIntLLRInputS4xD(142)(0) <= CNStageIntLLROutputS4xD(40)(2);
  VNStageIntLLRInputS4xD(206)(0) <= CNStageIntLLROutputS4xD(40)(3);
  VNStageIntLLRInputS4xD(270)(0) <= CNStageIntLLROutputS4xD(40)(4);
  VNStageIntLLRInputS4xD(334)(0) <= CNStageIntLLROutputS4xD(40)(5);
  VNStageIntLLRInputS4xD(12)(0) <= CNStageIntLLROutputS4xD(41)(0);
  VNStageIntLLRInputS4xD(76)(0) <= CNStageIntLLROutputS4xD(41)(1);
  VNStageIntLLRInputS4xD(140)(0) <= CNStageIntLLROutputS4xD(41)(2);
  VNStageIntLLRInputS4xD(204)(0) <= CNStageIntLLROutputS4xD(41)(3);
  VNStageIntLLRInputS4xD(268)(0) <= CNStageIntLLROutputS4xD(41)(4);
  VNStageIntLLRInputS4xD(332)(0) <= CNStageIntLLROutputS4xD(41)(5);
  VNStageIntLLRInputS4xD(11)(0) <= CNStageIntLLROutputS4xD(42)(0);
  VNStageIntLLRInputS4xD(75)(0) <= CNStageIntLLROutputS4xD(42)(1);
  VNStageIntLLRInputS4xD(139)(0) <= CNStageIntLLROutputS4xD(42)(2);
  VNStageIntLLRInputS4xD(203)(0) <= CNStageIntLLROutputS4xD(42)(3);
  VNStageIntLLRInputS4xD(267)(0) <= CNStageIntLLROutputS4xD(42)(4);
  VNStageIntLLRInputS4xD(331)(0) <= CNStageIntLLROutputS4xD(42)(5);
  VNStageIntLLRInputS4xD(10)(0) <= CNStageIntLLROutputS4xD(43)(0);
  VNStageIntLLRInputS4xD(74)(0) <= CNStageIntLLROutputS4xD(43)(1);
  VNStageIntLLRInputS4xD(138)(0) <= CNStageIntLLROutputS4xD(43)(2);
  VNStageIntLLRInputS4xD(202)(0) <= CNStageIntLLROutputS4xD(43)(3);
  VNStageIntLLRInputS4xD(266)(0) <= CNStageIntLLROutputS4xD(43)(4);
  VNStageIntLLRInputS4xD(330)(0) <= CNStageIntLLROutputS4xD(43)(5);
  VNStageIntLLRInputS4xD(9)(0) <= CNStageIntLLROutputS4xD(44)(0);
  VNStageIntLLRInputS4xD(73)(0) <= CNStageIntLLROutputS4xD(44)(1);
  VNStageIntLLRInputS4xD(137)(0) <= CNStageIntLLROutputS4xD(44)(2);
  VNStageIntLLRInputS4xD(201)(0) <= CNStageIntLLROutputS4xD(44)(3);
  VNStageIntLLRInputS4xD(265)(0) <= CNStageIntLLROutputS4xD(44)(4);
  VNStageIntLLRInputS4xD(329)(0) <= CNStageIntLLROutputS4xD(44)(5);
  VNStageIntLLRInputS4xD(8)(0) <= CNStageIntLLROutputS4xD(45)(0);
  VNStageIntLLRInputS4xD(72)(0) <= CNStageIntLLROutputS4xD(45)(1);
  VNStageIntLLRInputS4xD(136)(0) <= CNStageIntLLROutputS4xD(45)(2);
  VNStageIntLLRInputS4xD(200)(0) <= CNStageIntLLROutputS4xD(45)(3);
  VNStageIntLLRInputS4xD(264)(0) <= CNStageIntLLROutputS4xD(45)(4);
  VNStageIntLLRInputS4xD(328)(0) <= CNStageIntLLROutputS4xD(45)(5);
  VNStageIntLLRInputS4xD(7)(0) <= CNStageIntLLROutputS4xD(46)(0);
  VNStageIntLLRInputS4xD(71)(0) <= CNStageIntLLROutputS4xD(46)(1);
  VNStageIntLLRInputS4xD(135)(0) <= CNStageIntLLROutputS4xD(46)(2);
  VNStageIntLLRInputS4xD(199)(0) <= CNStageIntLLROutputS4xD(46)(3);
  VNStageIntLLRInputS4xD(263)(0) <= CNStageIntLLROutputS4xD(46)(4);
  VNStageIntLLRInputS4xD(327)(0) <= CNStageIntLLROutputS4xD(46)(5);
  VNStageIntLLRInputS4xD(6)(0) <= CNStageIntLLROutputS4xD(47)(0);
  VNStageIntLLRInputS4xD(70)(0) <= CNStageIntLLROutputS4xD(47)(1);
  VNStageIntLLRInputS4xD(134)(0) <= CNStageIntLLROutputS4xD(47)(2);
  VNStageIntLLRInputS4xD(198)(0) <= CNStageIntLLROutputS4xD(47)(3);
  VNStageIntLLRInputS4xD(262)(0) <= CNStageIntLLROutputS4xD(47)(4);
  VNStageIntLLRInputS4xD(326)(0) <= CNStageIntLLROutputS4xD(47)(5);
  VNStageIntLLRInputS4xD(5)(0) <= CNStageIntLLROutputS4xD(48)(0);
  VNStageIntLLRInputS4xD(69)(0) <= CNStageIntLLROutputS4xD(48)(1);
  VNStageIntLLRInputS4xD(133)(0) <= CNStageIntLLROutputS4xD(48)(2);
  VNStageIntLLRInputS4xD(197)(0) <= CNStageIntLLROutputS4xD(48)(3);
  VNStageIntLLRInputS4xD(261)(0) <= CNStageIntLLROutputS4xD(48)(4);
  VNStageIntLLRInputS4xD(325)(0) <= CNStageIntLLROutputS4xD(48)(5);
  VNStageIntLLRInputS4xD(4)(0) <= CNStageIntLLROutputS4xD(49)(0);
  VNStageIntLLRInputS4xD(68)(0) <= CNStageIntLLROutputS4xD(49)(1);
  VNStageIntLLRInputS4xD(132)(0) <= CNStageIntLLROutputS4xD(49)(2);
  VNStageIntLLRInputS4xD(196)(0) <= CNStageIntLLROutputS4xD(49)(3);
  VNStageIntLLRInputS4xD(260)(0) <= CNStageIntLLROutputS4xD(49)(4);
  VNStageIntLLRInputS4xD(324)(0) <= CNStageIntLLROutputS4xD(49)(5);
  VNStageIntLLRInputS4xD(2)(0) <= CNStageIntLLROutputS4xD(50)(0);
  VNStageIntLLRInputS4xD(66)(0) <= CNStageIntLLROutputS4xD(50)(1);
  VNStageIntLLRInputS4xD(130)(0) <= CNStageIntLLROutputS4xD(50)(2);
  VNStageIntLLRInputS4xD(194)(0) <= CNStageIntLLROutputS4xD(50)(3);
  VNStageIntLLRInputS4xD(258)(0) <= CNStageIntLLROutputS4xD(50)(4);
  VNStageIntLLRInputS4xD(322)(0) <= CNStageIntLLROutputS4xD(50)(5);
  VNStageIntLLRInputS4xD(1)(0) <= CNStageIntLLROutputS4xD(51)(0);
  VNStageIntLLRInputS4xD(65)(0) <= CNStageIntLLROutputS4xD(51)(1);
  VNStageIntLLRInputS4xD(129)(0) <= CNStageIntLLROutputS4xD(51)(2);
  VNStageIntLLRInputS4xD(193)(0) <= CNStageIntLLROutputS4xD(51)(3);
  VNStageIntLLRInputS4xD(257)(0) <= CNStageIntLLROutputS4xD(51)(4);
  VNStageIntLLRInputS4xD(321)(0) <= CNStageIntLLROutputS4xD(51)(5);
  VNStageIntLLRInputS4xD(63)(0) <= CNStageIntLLROutputS4xD(52)(0);
  VNStageIntLLRInputS4xD(127)(0) <= CNStageIntLLROutputS4xD(52)(1);
  VNStageIntLLRInputS4xD(191)(0) <= CNStageIntLLROutputS4xD(52)(2);
  VNStageIntLLRInputS4xD(255)(0) <= CNStageIntLLROutputS4xD(52)(3);
  VNStageIntLLRInputS4xD(319)(0) <= CNStageIntLLROutputS4xD(52)(4);
  VNStageIntLLRInputS4xD(383)(0) <= CNStageIntLLROutputS4xD(52)(5);
  VNStageIntLLRInputS4xD(0)(0) <= CNStageIntLLROutputS4xD(53)(0);
  VNStageIntLLRInputS4xD(64)(0) <= CNStageIntLLROutputS4xD(53)(1);
  VNStageIntLLRInputS4xD(128)(0) <= CNStageIntLLROutputS4xD(53)(2);
  VNStageIntLLRInputS4xD(192)(0) <= CNStageIntLLROutputS4xD(53)(3);
  VNStageIntLLRInputS4xD(256)(0) <= CNStageIntLLROutputS4xD(53)(4);
  VNStageIntLLRInputS4xD(320)(0) <= CNStageIntLLROutputS4xD(53)(5);
  VNStageIntLLRInputS4xD(42)(1) <= CNStageIntLLROutputS4xD(54)(0);
  VNStageIntLLRInputS4xD(112)(1) <= CNStageIntLLROutputS4xD(54)(1);
  VNStageIntLLRInputS4xD(182)(1) <= CNStageIntLLROutputS4xD(54)(2);
  VNStageIntLLRInputS4xD(203)(1) <= CNStageIntLLROutputS4xD(54)(3);
  VNStageIntLLRInputS4xD(259)(0) <= CNStageIntLLROutputS4xD(54)(4);
  VNStageIntLLRInputS4xD(361)(1) <= CNStageIntLLROutputS4xD(54)(5);
  VNStageIntLLRInputS4xD(41)(1) <= CNStageIntLLROutputS4xD(55)(0);
  VNStageIntLLRInputS4xD(117)(1) <= CNStageIntLLROutputS4xD(55)(1);
  VNStageIntLLRInputS4xD(138)(1) <= CNStageIntLLROutputS4xD(55)(2);
  VNStageIntLLRInputS4xD(194)(1) <= CNStageIntLLROutputS4xD(55)(3);
  VNStageIntLLRInputS4xD(296)(1) <= CNStageIntLLROutputS4xD(55)(4);
  VNStageIntLLRInputS4xD(362)(1) <= CNStageIntLLROutputS4xD(55)(5);
  VNStageIntLLRInputS4xD(40)(1) <= CNStageIntLLROutputS4xD(56)(0);
  VNStageIntLLRInputS4xD(73)(1) <= CNStageIntLLROutputS4xD(56)(1);
  VNStageIntLLRInputS4xD(129)(1) <= CNStageIntLLROutputS4xD(56)(2);
  VNStageIntLLRInputS4xD(231)(1) <= CNStageIntLLROutputS4xD(56)(3);
  VNStageIntLLRInputS4xD(297)(1) <= CNStageIntLLROutputS4xD(56)(4);
  VNStageIntLLRInputS4xD(323)(0) <= CNStageIntLLROutputS4xD(56)(5);
  VNStageIntLLRInputS4xD(39)(1) <= CNStageIntLLROutputS4xD(57)(0);
  VNStageIntLLRInputS4xD(127)(1) <= CNStageIntLLROutputS4xD(57)(1);
  VNStageIntLLRInputS4xD(166)(1) <= CNStageIntLLROutputS4xD(57)(2);
  VNStageIntLLRInputS4xD(232)(1) <= CNStageIntLLROutputS4xD(57)(3);
  VNStageIntLLRInputS4xD(258)(1) <= CNStageIntLLROutputS4xD(57)(4);
  VNStageIntLLRInputS4xD(344)(1) <= CNStageIntLLROutputS4xD(57)(5);
  VNStageIntLLRInputS4xD(38)(1) <= CNStageIntLLROutputS4xD(58)(0);
  VNStageIntLLRInputS4xD(101)(1) <= CNStageIntLLROutputS4xD(58)(1);
  VNStageIntLLRInputS4xD(167)(1) <= CNStageIntLLROutputS4xD(58)(2);
  VNStageIntLLRInputS4xD(193)(1) <= CNStageIntLLROutputS4xD(58)(3);
  VNStageIntLLRInputS4xD(279)(1) <= CNStageIntLLROutputS4xD(58)(4);
  VNStageIntLLRInputS4xD(340)(1) <= CNStageIntLLROutputS4xD(58)(5);
  VNStageIntLLRInputS4xD(37)(1) <= CNStageIntLLROutputS4xD(59)(0);
  VNStageIntLLRInputS4xD(102)(1) <= CNStageIntLLROutputS4xD(59)(1);
  VNStageIntLLRInputS4xD(191)(1) <= CNStageIntLLROutputS4xD(59)(2);
  VNStageIntLLRInputS4xD(214)(1) <= CNStageIntLLROutputS4xD(59)(3);
  VNStageIntLLRInputS4xD(275)(1) <= CNStageIntLLROutputS4xD(59)(4);
  VNStageIntLLRInputS4xD(355)(1) <= CNStageIntLLROutputS4xD(59)(5);
  VNStageIntLLRInputS4xD(36)(1) <= CNStageIntLLROutputS4xD(60)(0);
  VNStageIntLLRInputS4xD(126)(0) <= CNStageIntLLROutputS4xD(60)(1);
  VNStageIntLLRInputS4xD(149)(1) <= CNStageIntLLROutputS4xD(60)(2);
  VNStageIntLLRInputS4xD(210)(1) <= CNStageIntLLROutputS4xD(60)(3);
  VNStageIntLLRInputS4xD(290)(1) <= CNStageIntLLROutputS4xD(60)(4);
  VNStageIntLLRInputS4xD(381)(0) <= CNStageIntLLROutputS4xD(60)(5);
  VNStageIntLLRInputS4xD(35)(1) <= CNStageIntLLROutputS4xD(61)(0);
  VNStageIntLLRInputS4xD(84)(1) <= CNStageIntLLROutputS4xD(61)(1);
  VNStageIntLLRInputS4xD(145)(1) <= CNStageIntLLROutputS4xD(61)(2);
  VNStageIntLLRInputS4xD(225)(1) <= CNStageIntLLROutputS4xD(61)(3);
  VNStageIntLLRInputS4xD(316)(0) <= CNStageIntLLROutputS4xD(61)(4);
  VNStageIntLLRInputS4xD(357)(1) <= CNStageIntLLROutputS4xD(61)(5);
  VNStageIntLLRInputS4xD(34)(1) <= CNStageIntLLROutputS4xD(62)(0);
  VNStageIntLLRInputS4xD(80)(1) <= CNStageIntLLROutputS4xD(62)(1);
  VNStageIntLLRInputS4xD(160)(1) <= CNStageIntLLROutputS4xD(62)(2);
  VNStageIntLLRInputS4xD(251)(0) <= CNStageIntLLROutputS4xD(62)(3);
  VNStageIntLLRInputS4xD(292)(1) <= CNStageIntLLROutputS4xD(62)(4);
  VNStageIntLLRInputS4xD(326)(1) <= CNStageIntLLROutputS4xD(62)(5);
  VNStageIntLLRInputS4xD(33)(1) <= CNStageIntLLROutputS4xD(63)(0);
  VNStageIntLLRInputS4xD(95)(1) <= CNStageIntLLROutputS4xD(63)(1);
  VNStageIntLLRInputS4xD(186)(0) <= CNStageIntLLROutputS4xD(63)(2);
  VNStageIntLLRInputS4xD(227)(1) <= CNStageIntLLROutputS4xD(63)(3);
  VNStageIntLLRInputS4xD(261)(1) <= CNStageIntLLROutputS4xD(63)(4);
  VNStageIntLLRInputS4xD(342)(1) <= CNStageIntLLROutputS4xD(63)(5);
  VNStageIntLLRInputS4xD(32)(1) <= CNStageIntLLROutputS4xD(64)(0);
  VNStageIntLLRInputS4xD(121)(0) <= CNStageIntLLROutputS4xD(64)(1);
  VNStageIntLLRInputS4xD(162)(1) <= CNStageIntLLROutputS4xD(64)(2);
  VNStageIntLLRInputS4xD(196)(1) <= CNStageIntLLROutputS4xD(64)(3);
  VNStageIntLLRInputS4xD(277)(1) <= CNStageIntLLROutputS4xD(64)(4);
  VNStageIntLLRInputS4xD(375)(1) <= CNStageIntLLROutputS4xD(64)(5);
  VNStageIntLLRInputS4xD(31)(1) <= CNStageIntLLROutputS4xD(65)(0);
  VNStageIntLLRInputS4xD(97)(1) <= CNStageIntLLROutputS4xD(65)(1);
  VNStageIntLLRInputS4xD(131)(0) <= CNStageIntLLROutputS4xD(65)(2);
  VNStageIntLLRInputS4xD(212)(1) <= CNStageIntLLROutputS4xD(65)(3);
  VNStageIntLLRInputS4xD(310)(1) <= CNStageIntLLROutputS4xD(65)(4);
  VNStageIntLLRInputS4xD(321)(1) <= CNStageIntLLROutputS4xD(65)(5);
  VNStageIntLLRInputS4xD(30)(1) <= CNStageIntLLROutputS4xD(66)(0);
  VNStageIntLLRInputS4xD(66)(1) <= CNStageIntLLROutputS4xD(66)(1);
  VNStageIntLLRInputS4xD(147)(1) <= CNStageIntLLROutputS4xD(66)(2);
  VNStageIntLLRInputS4xD(245)(1) <= CNStageIntLLROutputS4xD(66)(3);
  VNStageIntLLRInputS4xD(319)(1) <= CNStageIntLLROutputS4xD(66)(4);
  VNStageIntLLRInputS4xD(334)(1) <= CNStageIntLLROutputS4xD(66)(5);
  VNStageIntLLRInputS4xD(29)(1) <= CNStageIntLLROutputS4xD(67)(0);
  VNStageIntLLRInputS4xD(82)(1) <= CNStageIntLLROutputS4xD(67)(1);
  VNStageIntLLRInputS4xD(180)(0) <= CNStageIntLLROutputS4xD(67)(2);
  VNStageIntLLRInputS4xD(254)(0) <= CNStageIntLLROutputS4xD(67)(3);
  VNStageIntLLRInputS4xD(269)(0) <= CNStageIntLLROutputS4xD(67)(4);
  VNStageIntLLRInputS4xD(376)(1) <= CNStageIntLLROutputS4xD(67)(5);
  VNStageIntLLRInputS4xD(28)(1) <= CNStageIntLLROutputS4xD(68)(0);
  VNStageIntLLRInputS4xD(115)(1) <= CNStageIntLLROutputS4xD(68)(1);
  VNStageIntLLRInputS4xD(189)(0) <= CNStageIntLLROutputS4xD(68)(2);
  VNStageIntLLRInputS4xD(204)(1) <= CNStageIntLLROutputS4xD(68)(3);
  VNStageIntLLRInputS4xD(311)(1) <= CNStageIntLLROutputS4xD(68)(4);
  VNStageIntLLRInputS4xD(341)(1) <= CNStageIntLLROutputS4xD(68)(5);
  VNStageIntLLRInputS4xD(27)(1) <= CNStageIntLLROutputS4xD(69)(0);
  VNStageIntLLRInputS4xD(124)(0) <= CNStageIntLLROutputS4xD(69)(1);
  VNStageIntLLRInputS4xD(139)(1) <= CNStageIntLLROutputS4xD(69)(2);
  VNStageIntLLRInputS4xD(246)(1) <= CNStageIntLLROutputS4xD(69)(3);
  VNStageIntLLRInputS4xD(276)(1) <= CNStageIntLLROutputS4xD(69)(4);
  VNStageIntLLRInputS4xD(343)(1) <= CNStageIntLLROutputS4xD(69)(5);
  VNStageIntLLRInputS4xD(26)(1) <= CNStageIntLLROutputS4xD(70)(0);
  VNStageIntLLRInputS4xD(74)(1) <= CNStageIntLLROutputS4xD(70)(1);
  VNStageIntLLRInputS4xD(181)(1) <= CNStageIntLLROutputS4xD(70)(2);
  VNStageIntLLRInputS4xD(211)(1) <= CNStageIntLLROutputS4xD(70)(3);
  VNStageIntLLRInputS4xD(278)(1) <= CNStageIntLLROutputS4xD(70)(4);
  VNStageIntLLRInputS4xD(325)(1) <= CNStageIntLLROutputS4xD(70)(5);
  VNStageIntLLRInputS4xD(25)(1) <= CNStageIntLLROutputS4xD(71)(0);
  VNStageIntLLRInputS4xD(116)(0) <= CNStageIntLLROutputS4xD(71)(1);
  VNStageIntLLRInputS4xD(146)(1) <= CNStageIntLLROutputS4xD(71)(2);
  VNStageIntLLRInputS4xD(213)(1) <= CNStageIntLLROutputS4xD(71)(3);
  VNStageIntLLRInputS4xD(260)(1) <= CNStageIntLLROutputS4xD(71)(4);
  VNStageIntLLRInputS4xD(332)(1) <= CNStageIntLLROutputS4xD(71)(5);
  VNStageIntLLRInputS4xD(24)(1) <= CNStageIntLLROutputS4xD(72)(0);
  VNStageIntLLRInputS4xD(81)(1) <= CNStageIntLLROutputS4xD(72)(1);
  VNStageIntLLRInputS4xD(148)(1) <= CNStageIntLLROutputS4xD(72)(2);
  VNStageIntLLRInputS4xD(195)(0) <= CNStageIntLLROutputS4xD(72)(3);
  VNStageIntLLRInputS4xD(267)(1) <= CNStageIntLLROutputS4xD(72)(4);
  VNStageIntLLRInputS4xD(359)(1) <= CNStageIntLLROutputS4xD(72)(5);
  VNStageIntLLRInputS4xD(23)(1) <= CNStageIntLLROutputS4xD(73)(0);
  VNStageIntLLRInputS4xD(83)(1) <= CNStageIntLLROutputS4xD(73)(1);
  VNStageIntLLRInputS4xD(130)(1) <= CNStageIntLLROutputS4xD(73)(2);
  VNStageIntLLRInputS4xD(202)(1) <= CNStageIntLLROutputS4xD(73)(3);
  VNStageIntLLRInputS4xD(294)(1) <= CNStageIntLLROutputS4xD(73)(4);
  VNStageIntLLRInputS4xD(347)(1) <= CNStageIntLLROutputS4xD(73)(5);
  VNStageIntLLRInputS4xD(22)(1) <= CNStageIntLLROutputS4xD(74)(0);
  VNStageIntLLRInputS4xD(65)(1) <= CNStageIntLLROutputS4xD(74)(1);
  VNStageIntLLRInputS4xD(137)(1) <= CNStageIntLLROutputS4xD(74)(2);
  VNStageIntLLRInputS4xD(229)(1) <= CNStageIntLLROutputS4xD(74)(3);
  VNStageIntLLRInputS4xD(282)(1) <= CNStageIntLLROutputS4xD(74)(4);
  VNStageIntLLRInputS4xD(353)(1) <= CNStageIntLLROutputS4xD(74)(5);
  VNStageIntLLRInputS4xD(21)(1) <= CNStageIntLLROutputS4xD(75)(0);
  VNStageIntLLRInputS4xD(72)(1) <= CNStageIntLLROutputS4xD(75)(1);
  VNStageIntLLRInputS4xD(164)(1) <= CNStageIntLLROutputS4xD(75)(2);
  VNStageIntLLRInputS4xD(217)(1) <= CNStageIntLLROutputS4xD(75)(3);
  VNStageIntLLRInputS4xD(288)(1) <= CNStageIntLLROutputS4xD(75)(4);
  VNStageIntLLRInputS4xD(348)(1) <= CNStageIntLLROutputS4xD(75)(5);
  VNStageIntLLRInputS4xD(20)(1) <= CNStageIntLLROutputS4xD(76)(0);
  VNStageIntLLRInputS4xD(99)(1) <= CNStageIntLLROutputS4xD(76)(1);
  VNStageIntLLRInputS4xD(152)(1) <= CNStageIntLLROutputS4xD(76)(2);
  VNStageIntLLRInputS4xD(223)(1) <= CNStageIntLLROutputS4xD(76)(3);
  VNStageIntLLRInputS4xD(283)(1) <= CNStageIntLLROutputS4xD(76)(4);
  VNStageIntLLRInputS4xD(358)(1) <= CNStageIntLLROutputS4xD(76)(5);
  VNStageIntLLRInputS4xD(19)(1) <= CNStageIntLLROutputS4xD(77)(0);
  VNStageIntLLRInputS4xD(87)(1) <= CNStageIntLLROutputS4xD(77)(1);
  VNStageIntLLRInputS4xD(158)(1) <= CNStageIntLLROutputS4xD(77)(2);
  VNStageIntLLRInputS4xD(218)(1) <= CNStageIntLLROutputS4xD(77)(3);
  VNStageIntLLRInputS4xD(293)(1) <= CNStageIntLLROutputS4xD(77)(4);
  VNStageIntLLRInputS4xD(380)(0) <= CNStageIntLLROutputS4xD(77)(5);
  VNStageIntLLRInputS4xD(18)(1) <= CNStageIntLLROutputS4xD(78)(0);
  VNStageIntLLRInputS4xD(93)(1) <= CNStageIntLLROutputS4xD(78)(1);
  VNStageIntLLRInputS4xD(153)(1) <= CNStageIntLLROutputS4xD(78)(2);
  VNStageIntLLRInputS4xD(228)(1) <= CNStageIntLLROutputS4xD(78)(3);
  VNStageIntLLRInputS4xD(315)(0) <= CNStageIntLLROutputS4xD(78)(4);
  VNStageIntLLRInputS4xD(335)(1) <= CNStageIntLLROutputS4xD(78)(5);
  VNStageIntLLRInputS4xD(17)(1) <= CNStageIntLLROutputS4xD(79)(0);
  VNStageIntLLRInputS4xD(88)(1) <= CNStageIntLLROutputS4xD(79)(1);
  VNStageIntLLRInputS4xD(163)(1) <= CNStageIntLLROutputS4xD(79)(2);
  VNStageIntLLRInputS4xD(250)(0) <= CNStageIntLLROutputS4xD(79)(3);
  VNStageIntLLRInputS4xD(270)(1) <= CNStageIntLLROutputS4xD(79)(4);
  VNStageIntLLRInputS4xD(383)(1) <= CNStageIntLLROutputS4xD(79)(5);
  VNStageIntLLRInputS4xD(15)(1) <= CNStageIntLLROutputS4xD(80)(0);
  VNStageIntLLRInputS4xD(120)(1) <= CNStageIntLLROutputS4xD(80)(1);
  VNStageIntLLRInputS4xD(140)(1) <= CNStageIntLLROutputS4xD(80)(2);
  VNStageIntLLRInputS4xD(253)(0) <= CNStageIntLLROutputS4xD(80)(3);
  VNStageIntLLRInputS4xD(305)(1) <= CNStageIntLLROutputS4xD(80)(4);
  VNStageIntLLRInputS4xD(338)(1) <= CNStageIntLLROutputS4xD(80)(5);
  VNStageIntLLRInputS4xD(14)(1) <= CNStageIntLLROutputS4xD(81)(0);
  VNStageIntLLRInputS4xD(75)(1) <= CNStageIntLLROutputS4xD(81)(1);
  VNStageIntLLRInputS4xD(188)(0) <= CNStageIntLLROutputS4xD(81)(2);
  VNStageIntLLRInputS4xD(240)(1) <= CNStageIntLLROutputS4xD(81)(3);
  VNStageIntLLRInputS4xD(273)(1) <= CNStageIntLLROutputS4xD(81)(4);
  VNStageIntLLRInputS4xD(350)(1) <= CNStageIntLLROutputS4xD(81)(5);
  VNStageIntLLRInputS4xD(13)(0) <= CNStageIntLLROutputS4xD(82)(0);
  VNStageIntLLRInputS4xD(123)(0) <= CNStageIntLLROutputS4xD(82)(1);
  VNStageIntLLRInputS4xD(175)(1) <= CNStageIntLLROutputS4xD(82)(2);
  VNStageIntLLRInputS4xD(208)(1) <= CNStageIntLLROutputS4xD(82)(3);
  VNStageIntLLRInputS4xD(285)(1) <= CNStageIntLLROutputS4xD(82)(4);
  VNStageIntLLRInputS4xD(364)(1) <= CNStageIntLLROutputS4xD(82)(5);
  VNStageIntLLRInputS4xD(12)(1) <= CNStageIntLLROutputS4xD(83)(0);
  VNStageIntLLRInputS4xD(110)(1) <= CNStageIntLLROutputS4xD(83)(1);
  VNStageIntLLRInputS4xD(143)(1) <= CNStageIntLLROutputS4xD(83)(2);
  VNStageIntLLRInputS4xD(220)(1) <= CNStageIntLLROutputS4xD(83)(3);
  VNStageIntLLRInputS4xD(299)(0) <= CNStageIntLLROutputS4xD(83)(4);
  VNStageIntLLRInputS4xD(345)(1) <= CNStageIntLLROutputS4xD(83)(5);
  VNStageIntLLRInputS4xD(11)(1) <= CNStageIntLLROutputS4xD(84)(0);
  VNStageIntLLRInputS4xD(78)(1) <= CNStageIntLLROutputS4xD(84)(1);
  VNStageIntLLRInputS4xD(155)(1) <= CNStageIntLLROutputS4xD(84)(2);
  VNStageIntLLRInputS4xD(234)(1) <= CNStageIntLLROutputS4xD(84)(3);
  VNStageIntLLRInputS4xD(280)(1) <= CNStageIntLLROutputS4xD(84)(4);
  VNStageIntLLRInputS4xD(322)(1) <= CNStageIntLLROutputS4xD(84)(5);
  VNStageIntLLRInputS4xD(10)(1) <= CNStageIntLLROutputS4xD(85)(0);
  VNStageIntLLRInputS4xD(90)(1) <= CNStageIntLLROutputS4xD(85)(1);
  VNStageIntLLRInputS4xD(169)(1) <= CNStageIntLLROutputS4xD(85)(2);
  VNStageIntLLRInputS4xD(215)(1) <= CNStageIntLLROutputS4xD(85)(3);
  VNStageIntLLRInputS4xD(257)(1) <= CNStageIntLLROutputS4xD(85)(4);
  VNStageIntLLRInputS4xD(374)(1) <= CNStageIntLLROutputS4xD(85)(5);
  VNStageIntLLRInputS4xD(9)(1) <= CNStageIntLLROutputS4xD(86)(0);
  VNStageIntLLRInputS4xD(104)(1) <= CNStageIntLLROutputS4xD(86)(1);
  VNStageIntLLRInputS4xD(150)(1) <= CNStageIntLLROutputS4xD(86)(2);
  VNStageIntLLRInputS4xD(255)(1) <= CNStageIntLLROutputS4xD(86)(3);
  VNStageIntLLRInputS4xD(309)(1) <= CNStageIntLLROutputS4xD(86)(4);
  VNStageIntLLRInputS4xD(378)(0) <= CNStageIntLLROutputS4xD(86)(5);
  VNStageIntLLRInputS4xD(7)(1) <= CNStageIntLLROutputS4xD(87)(0);
  VNStageIntLLRInputS4xD(125)(0) <= CNStageIntLLROutputS4xD(87)(1);
  VNStageIntLLRInputS4xD(179)(1) <= CNStageIntLLROutputS4xD(87)(2);
  VNStageIntLLRInputS4xD(248)(1) <= CNStageIntLLROutputS4xD(87)(3);
  VNStageIntLLRInputS4xD(306)(1) <= CNStageIntLLROutputS4xD(87)(4);
  VNStageIntLLRInputS4xD(382)(0) <= CNStageIntLLROutputS4xD(87)(5);
  VNStageIntLLRInputS4xD(6)(1) <= CNStageIntLLROutputS4xD(88)(0);
  VNStageIntLLRInputS4xD(114)(1) <= CNStageIntLLROutputS4xD(88)(1);
  VNStageIntLLRInputS4xD(183)(1) <= CNStageIntLLROutputS4xD(88)(2);
  VNStageIntLLRInputS4xD(241)(1) <= CNStageIntLLROutputS4xD(88)(3);
  VNStageIntLLRInputS4xD(317)(0) <= CNStageIntLLROutputS4xD(88)(4);
  VNStageIntLLRInputS4xD(354)(1) <= CNStageIntLLROutputS4xD(88)(5);
  VNStageIntLLRInputS4xD(5)(1) <= CNStageIntLLROutputS4xD(89)(0);
  VNStageIntLLRInputS4xD(118)(1) <= CNStageIntLLROutputS4xD(89)(1);
  VNStageIntLLRInputS4xD(176)(1) <= CNStageIntLLROutputS4xD(89)(2);
  VNStageIntLLRInputS4xD(252)(0) <= CNStageIntLLROutputS4xD(89)(3);
  VNStageIntLLRInputS4xD(289)(1) <= CNStageIntLLROutputS4xD(89)(4);
  VNStageIntLLRInputS4xD(346)(1) <= CNStageIntLLROutputS4xD(89)(5);
  VNStageIntLLRInputS4xD(4)(1) <= CNStageIntLLROutputS4xD(90)(0);
  VNStageIntLLRInputS4xD(111)(1) <= CNStageIntLLROutputS4xD(90)(1);
  VNStageIntLLRInputS4xD(187)(0) <= CNStageIntLLROutputS4xD(90)(2);
  VNStageIntLLRInputS4xD(224)(1) <= CNStageIntLLROutputS4xD(90)(3);
  VNStageIntLLRInputS4xD(281)(1) <= CNStageIntLLROutputS4xD(90)(4);
  VNStageIntLLRInputS4xD(363)(0) <= CNStageIntLLROutputS4xD(90)(5);
  VNStageIntLLRInputS4xD(3)(0) <= CNStageIntLLROutputS4xD(91)(0);
  VNStageIntLLRInputS4xD(122)(0) <= CNStageIntLLROutputS4xD(91)(1);
  VNStageIntLLRInputS4xD(159)(1) <= CNStageIntLLROutputS4xD(91)(2);
  VNStageIntLLRInputS4xD(216)(1) <= CNStageIntLLROutputS4xD(91)(3);
  VNStageIntLLRInputS4xD(298)(1) <= CNStageIntLLROutputS4xD(91)(4);
  VNStageIntLLRInputS4xD(360)(1) <= CNStageIntLLROutputS4xD(91)(5);
  VNStageIntLLRInputS4xD(2)(1) <= CNStageIntLLROutputS4xD(92)(0);
  VNStageIntLLRInputS4xD(94)(1) <= CNStageIntLLROutputS4xD(92)(1);
  VNStageIntLLRInputS4xD(151)(1) <= CNStageIntLLROutputS4xD(92)(2);
  VNStageIntLLRInputS4xD(233)(1) <= CNStageIntLLROutputS4xD(92)(3);
  VNStageIntLLRInputS4xD(295)(1) <= CNStageIntLLROutputS4xD(92)(4);
  VNStageIntLLRInputS4xD(331)(1) <= CNStageIntLLROutputS4xD(92)(5);
  VNStageIntLLRInputS4xD(63)(1) <= CNStageIntLLROutputS4xD(93)(0);
  VNStageIntLLRInputS4xD(103)(1) <= CNStageIntLLROutputS4xD(93)(1);
  VNStageIntLLRInputS4xD(165)(1) <= CNStageIntLLROutputS4xD(93)(2);
  VNStageIntLLRInputS4xD(201)(1) <= CNStageIntLLROutputS4xD(93)(3);
  VNStageIntLLRInputS4xD(286)(1) <= CNStageIntLLROutputS4xD(93)(4);
  VNStageIntLLRInputS4xD(337)(1) <= CNStageIntLLROutputS4xD(93)(5);
  VNStageIntLLRInputS4xD(62)(0) <= CNStageIntLLROutputS4xD(94)(0);
  VNStageIntLLRInputS4xD(100)(1) <= CNStageIntLLROutputS4xD(94)(1);
  VNStageIntLLRInputS4xD(136)(1) <= CNStageIntLLROutputS4xD(94)(2);
  VNStageIntLLRInputS4xD(221)(1) <= CNStageIntLLROutputS4xD(94)(3);
  VNStageIntLLRInputS4xD(272)(1) <= CNStageIntLLROutputS4xD(94)(4);
  VNStageIntLLRInputS4xD(327)(1) <= CNStageIntLLROutputS4xD(94)(5);
  VNStageIntLLRInputS4xD(61)(0) <= CNStageIntLLROutputS4xD(95)(0);
  VNStageIntLLRInputS4xD(71)(1) <= CNStageIntLLROutputS4xD(95)(1);
  VNStageIntLLRInputS4xD(156)(1) <= CNStageIntLLROutputS4xD(95)(2);
  VNStageIntLLRInputS4xD(207)(1) <= CNStageIntLLROutputS4xD(95)(3);
  VNStageIntLLRInputS4xD(262)(1) <= CNStageIntLLROutputS4xD(95)(4);
  VNStageIntLLRInputS4xD(356)(1) <= CNStageIntLLROutputS4xD(95)(5);
  VNStageIntLLRInputS4xD(60)(0) <= CNStageIntLLROutputS4xD(96)(0);
  VNStageIntLLRInputS4xD(91)(1) <= CNStageIntLLROutputS4xD(96)(1);
  VNStageIntLLRInputS4xD(142)(1) <= CNStageIntLLROutputS4xD(96)(2);
  VNStageIntLLRInputS4xD(197)(1) <= CNStageIntLLROutputS4xD(96)(3);
  VNStageIntLLRInputS4xD(291)(1) <= CNStageIntLLROutputS4xD(96)(4);
  VNStageIntLLRInputS4xD(339)(1) <= CNStageIntLLROutputS4xD(96)(5);
  VNStageIntLLRInputS4xD(58)(0) <= CNStageIntLLROutputS4xD(97)(0);
  VNStageIntLLRInputS4xD(67)(0) <= CNStageIntLLROutputS4xD(97)(1);
  VNStageIntLLRInputS4xD(161)(1) <= CNStageIntLLROutputS4xD(97)(2);
  VNStageIntLLRInputS4xD(209)(1) <= CNStageIntLLROutputS4xD(97)(3);
  VNStageIntLLRInputS4xD(304)(1) <= CNStageIntLLROutputS4xD(97)(4);
  VNStageIntLLRInputS4xD(329)(1) <= CNStageIntLLROutputS4xD(97)(5);
  VNStageIntLLRInputS4xD(57)(0) <= CNStageIntLLROutputS4xD(98)(0);
  VNStageIntLLRInputS4xD(96)(1) <= CNStageIntLLROutputS4xD(98)(1);
  VNStageIntLLRInputS4xD(144)(1) <= CNStageIntLLROutputS4xD(98)(2);
  VNStageIntLLRInputS4xD(239)(1) <= CNStageIntLLROutputS4xD(98)(3);
  VNStageIntLLRInputS4xD(264)(1) <= CNStageIntLLROutputS4xD(98)(4);
  VNStageIntLLRInputS4xD(365)(1) <= CNStageIntLLROutputS4xD(98)(5);
  VNStageIntLLRInputS4xD(56)(1) <= CNStageIntLLROutputS4xD(99)(0);
  VNStageIntLLRInputS4xD(79)(1) <= CNStageIntLLROutputS4xD(99)(1);
  VNStageIntLLRInputS4xD(174)(1) <= CNStageIntLLROutputS4xD(99)(2);
  VNStageIntLLRInputS4xD(199)(1) <= CNStageIntLLROutputS4xD(99)(3);
  VNStageIntLLRInputS4xD(300)(1) <= CNStageIntLLROutputS4xD(99)(4);
  VNStageIntLLRInputS4xD(349)(1) <= CNStageIntLLROutputS4xD(99)(5);
  VNStageIntLLRInputS4xD(55)(1) <= CNStageIntLLROutputS4xD(100)(0);
  VNStageIntLLRInputS4xD(109)(1) <= CNStageIntLLROutputS4xD(100)(1);
  VNStageIntLLRInputS4xD(134)(1) <= CNStageIntLLROutputS4xD(100)(2);
  VNStageIntLLRInputS4xD(235)(0) <= CNStageIntLLROutputS4xD(100)(3);
  VNStageIntLLRInputS4xD(284)(1) <= CNStageIntLLROutputS4xD(100)(4);
  VNStageIntLLRInputS4xD(352)(1) <= CNStageIntLLROutputS4xD(100)(5);
  VNStageIntLLRInputS4xD(54)(1) <= CNStageIntLLROutputS4xD(101)(0);
  VNStageIntLLRInputS4xD(69)(1) <= CNStageIntLLROutputS4xD(101)(1);
  VNStageIntLLRInputS4xD(170)(1) <= CNStageIntLLROutputS4xD(101)(2);
  VNStageIntLLRInputS4xD(219)(1) <= CNStageIntLLROutputS4xD(101)(3);
  VNStageIntLLRInputS4xD(287)(1) <= CNStageIntLLROutputS4xD(101)(4);
  VNStageIntLLRInputS4xD(330)(1) <= CNStageIntLLROutputS4xD(101)(5);
  VNStageIntLLRInputS4xD(52)(0) <= CNStageIntLLROutputS4xD(102)(0);
  VNStageIntLLRInputS4xD(89)(1) <= CNStageIntLLROutputS4xD(102)(1);
  VNStageIntLLRInputS4xD(157)(1) <= CNStageIntLLROutputS4xD(102)(2);
  VNStageIntLLRInputS4xD(200)(1) <= CNStageIntLLROutputS4xD(102)(3);
  VNStageIntLLRInputS4xD(303)(1) <= CNStageIntLLROutputS4xD(102)(4);
  VNStageIntLLRInputS4xD(366)(1) <= CNStageIntLLROutputS4xD(102)(5);
  VNStageIntLLRInputS4xD(51)(1) <= CNStageIntLLROutputS4xD(103)(0);
  VNStageIntLLRInputS4xD(92)(1) <= CNStageIntLLROutputS4xD(103)(1);
  VNStageIntLLRInputS4xD(135)(1) <= CNStageIntLLROutputS4xD(103)(2);
  VNStageIntLLRInputS4xD(238)(1) <= CNStageIntLLROutputS4xD(103)(3);
  VNStageIntLLRInputS4xD(301)(1) <= CNStageIntLLROutputS4xD(103)(4);
  VNStageIntLLRInputS4xD(328)(1) <= CNStageIntLLROutputS4xD(103)(5);
  VNStageIntLLRInputS4xD(50)(1) <= CNStageIntLLROutputS4xD(104)(0);
  VNStageIntLLRInputS4xD(70)(1) <= CNStageIntLLROutputS4xD(104)(1);
  VNStageIntLLRInputS4xD(173)(1) <= CNStageIntLLROutputS4xD(104)(2);
  VNStageIntLLRInputS4xD(236)(1) <= CNStageIntLLROutputS4xD(104)(3);
  VNStageIntLLRInputS4xD(263)(1) <= CNStageIntLLROutputS4xD(104)(4);
  VNStageIntLLRInputS4xD(336)(1) <= CNStageIntLLROutputS4xD(104)(5);
  VNStageIntLLRInputS4xD(49)(1) <= CNStageIntLLROutputS4xD(105)(0);
  VNStageIntLLRInputS4xD(108)(1) <= CNStageIntLLROutputS4xD(105)(1);
  VNStageIntLLRInputS4xD(171)(0) <= CNStageIntLLROutputS4xD(105)(2);
  VNStageIntLLRInputS4xD(198)(1) <= CNStageIntLLROutputS4xD(105)(3);
  VNStageIntLLRInputS4xD(271)(1) <= CNStageIntLLROutputS4xD(105)(4);
  VNStageIntLLRInputS4xD(379)(0) <= CNStageIntLLROutputS4xD(105)(5);
  VNStageIntLLRInputS4xD(46)(1) <= CNStageIntLLROutputS4xD(106)(0);
  VNStageIntLLRInputS4xD(76)(1) <= CNStageIntLLROutputS4xD(106)(1);
  VNStageIntLLRInputS4xD(184)(1) <= CNStageIntLLROutputS4xD(106)(2);
  VNStageIntLLRInputS4xD(243)(1) <= CNStageIntLLROutputS4xD(106)(3);
  VNStageIntLLRInputS4xD(256)(1) <= CNStageIntLLROutputS4xD(106)(4);
  VNStageIntLLRInputS4xD(372)(0) <= CNStageIntLLROutputS4xD(106)(5);
  VNStageIntLLRInputS4xD(45)(1) <= CNStageIntLLROutputS4xD(107)(0);
  VNStageIntLLRInputS4xD(119)(1) <= CNStageIntLLROutputS4xD(107)(1);
  VNStageIntLLRInputS4xD(178)(1) <= CNStageIntLLROutputS4xD(107)(2);
  VNStageIntLLRInputS4xD(192)(1) <= CNStageIntLLROutputS4xD(107)(3);
  VNStageIntLLRInputS4xD(307)(1) <= CNStageIntLLROutputS4xD(107)(4);
  VNStageIntLLRInputS4xD(377)(0) <= CNStageIntLLROutputS4xD(107)(5);
  VNStageIntLLRInputS4xD(44)(1) <= CNStageIntLLROutputS4xD(108)(0);
  VNStageIntLLRInputS4xD(113)(1) <= CNStageIntLLROutputS4xD(108)(1);
  VNStageIntLLRInputS4xD(128)(1) <= CNStageIntLLROutputS4xD(108)(2);
  VNStageIntLLRInputS4xD(242)(1) <= CNStageIntLLROutputS4xD(108)(3);
  VNStageIntLLRInputS4xD(312)(1) <= CNStageIntLLROutputS4xD(108)(4);
  VNStageIntLLRInputS4xD(333)(0) <= CNStageIntLLROutputS4xD(108)(5);
  VNStageIntLLRInputS4xD(43)(0) <= CNStageIntLLROutputS4xD(109)(0);
  VNStageIntLLRInputS4xD(64)(1) <= CNStageIntLLROutputS4xD(109)(1);
  VNStageIntLLRInputS4xD(177)(1) <= CNStageIntLLROutputS4xD(109)(2);
  VNStageIntLLRInputS4xD(247)(1) <= CNStageIntLLROutputS4xD(109)(3);
  VNStageIntLLRInputS4xD(268)(1) <= CNStageIntLLROutputS4xD(109)(4);
  VNStageIntLLRInputS4xD(324)(1) <= CNStageIntLLROutputS4xD(109)(5);
  VNStageIntLLRInputS4xD(0)(1) <= CNStageIntLLROutputS4xD(110)(0);
  VNStageIntLLRInputS4xD(107)(0) <= CNStageIntLLROutputS4xD(110)(1);
  VNStageIntLLRInputS4xD(172)(1) <= CNStageIntLLROutputS4xD(110)(2);
  VNStageIntLLRInputS4xD(237)(1) <= CNStageIntLLROutputS4xD(110)(3);
  VNStageIntLLRInputS4xD(302)(1) <= CNStageIntLLROutputS4xD(110)(4);
  VNStageIntLLRInputS4xD(367)(1) <= CNStageIntLLROutputS4xD(110)(5);
  VNStageIntLLRInputS4xD(32)(2) <= CNStageIntLLROutputS4xD(111)(0);
  VNStageIntLLRInputS4xD(117)(2) <= CNStageIntLLROutputS4xD(111)(1);
  VNStageIntLLRInputS4xD(136)(2) <= CNStageIntLLROutputS4xD(111)(2);
  VNStageIntLLRInputS4xD(198)(2) <= CNStageIntLLROutputS4xD(111)(3);
  VNStageIntLLRInputS4xD(297)(2) <= CNStageIntLLROutputS4xD(111)(4);
  VNStageIntLLRInputS4xD(382)(1) <= CNStageIntLLROutputS4xD(111)(5);
  VNStageIntLLRInputS4xD(30)(2) <= CNStageIntLLROutputS4xD(112)(0);
  VNStageIntLLRInputS4xD(68)(1) <= CNStageIntLLROutputS4xD(112)(1);
  VNStageIntLLRInputS4xD(167)(2) <= CNStageIntLLROutputS4xD(112)(2);
  VNStageIntLLRInputS4xD(252)(1) <= CNStageIntLLROutputS4xD(112)(3);
  VNStageIntLLRInputS4xD(303)(2) <= CNStageIntLLROutputS4xD(112)(4);
  VNStageIntLLRInputS4xD(358)(2) <= CNStageIntLLROutputS4xD(112)(5);
  VNStageIntLLRInputS4xD(29)(2) <= CNStageIntLLROutputS4xD(113)(0);
  VNStageIntLLRInputS4xD(102)(2) <= CNStageIntLLROutputS4xD(113)(1);
  VNStageIntLLRInputS4xD(187)(1) <= CNStageIntLLROutputS4xD(113)(2);
  VNStageIntLLRInputS4xD(238)(2) <= CNStageIntLLROutputS4xD(113)(3);
  VNStageIntLLRInputS4xD(293)(2) <= CNStageIntLLROutputS4xD(113)(4);
  VNStageIntLLRInputS4xD(324)(2) <= CNStageIntLLROutputS4xD(113)(5);
  VNStageIntLLRInputS4xD(28)(2) <= CNStageIntLLROutputS4xD(114)(0);
  VNStageIntLLRInputS4xD(122)(1) <= CNStageIntLLROutputS4xD(114)(1);
  VNStageIntLLRInputS4xD(173)(2) <= CNStageIntLLROutputS4xD(114)(2);
  VNStageIntLLRInputS4xD(228)(2) <= CNStageIntLLROutputS4xD(114)(3);
  VNStageIntLLRInputS4xD(259)(1) <= CNStageIntLLROutputS4xD(114)(4);
  VNStageIntLLRInputS4xD(370)(1) <= CNStageIntLLROutputS4xD(114)(5);
  VNStageIntLLRInputS4xD(27)(2) <= CNStageIntLLROutputS4xD(115)(0);
  VNStageIntLLRInputS4xD(108)(2) <= CNStageIntLLROutputS4xD(115)(1);
  VNStageIntLLRInputS4xD(163)(2) <= CNStageIntLLROutputS4xD(115)(2);
  VNStageIntLLRInputS4xD(194)(2) <= CNStageIntLLROutputS4xD(115)(3);
  VNStageIntLLRInputS4xD(305)(2) <= CNStageIntLLROutputS4xD(115)(4);
  VNStageIntLLRInputS4xD(337)(2) <= CNStageIntLLROutputS4xD(115)(5);
  VNStageIntLLRInputS4xD(26)(2) <= CNStageIntLLROutputS4xD(116)(0);
  VNStageIntLLRInputS4xD(98)(1) <= CNStageIntLLROutputS4xD(116)(1);
  VNStageIntLLRInputS4xD(129)(2) <= CNStageIntLLROutputS4xD(116)(2);
  VNStageIntLLRInputS4xD(240)(2) <= CNStageIntLLROutputS4xD(116)(3);
  VNStageIntLLRInputS4xD(272)(2) <= CNStageIntLLROutputS4xD(116)(4);
  VNStageIntLLRInputS4xD(360)(2) <= CNStageIntLLROutputS4xD(116)(5);
  VNStageIntLLRInputS4xD(25)(2) <= CNStageIntLLROutputS4xD(117)(0);
  VNStageIntLLRInputS4xD(127)(2) <= CNStageIntLLROutputS4xD(117)(1);
  VNStageIntLLRInputS4xD(175)(2) <= CNStageIntLLROutputS4xD(117)(2);
  VNStageIntLLRInputS4xD(207)(2) <= CNStageIntLLROutputS4xD(117)(3);
  VNStageIntLLRInputS4xD(295)(2) <= CNStageIntLLROutputS4xD(117)(4);
  VNStageIntLLRInputS4xD(333)(1) <= CNStageIntLLROutputS4xD(117)(5);
  VNStageIntLLRInputS4xD(24)(2) <= CNStageIntLLROutputS4xD(118)(0);
  VNStageIntLLRInputS4xD(110)(2) <= CNStageIntLLROutputS4xD(118)(1);
  VNStageIntLLRInputS4xD(142)(2) <= CNStageIntLLROutputS4xD(118)(2);
  VNStageIntLLRInputS4xD(230)(1) <= CNStageIntLLROutputS4xD(118)(3);
  VNStageIntLLRInputS4xD(268)(2) <= CNStageIntLLROutputS4xD(118)(4);
  VNStageIntLLRInputS4xD(380)(1) <= CNStageIntLLROutputS4xD(118)(5);
  VNStageIntLLRInputS4xD(23)(2) <= CNStageIntLLROutputS4xD(119)(0);
  VNStageIntLLRInputS4xD(77)(0) <= CNStageIntLLROutputS4xD(119)(1);
  VNStageIntLLRInputS4xD(165)(2) <= CNStageIntLLROutputS4xD(119)(2);
  VNStageIntLLRInputS4xD(203)(2) <= CNStageIntLLROutputS4xD(119)(3);
  VNStageIntLLRInputS4xD(315)(1) <= CNStageIntLLROutputS4xD(119)(4);
  VNStageIntLLRInputS4xD(383)(2) <= CNStageIntLLROutputS4xD(119)(5);
  VNStageIntLLRInputS4xD(22)(2) <= CNStageIntLLROutputS4xD(120)(0);
  VNStageIntLLRInputS4xD(100)(2) <= CNStageIntLLROutputS4xD(120)(1);
  VNStageIntLLRInputS4xD(138)(2) <= CNStageIntLLROutputS4xD(120)(2);
  VNStageIntLLRInputS4xD(250)(1) <= CNStageIntLLROutputS4xD(120)(3);
  VNStageIntLLRInputS4xD(318)(0) <= CNStageIntLLROutputS4xD(120)(4);
  VNStageIntLLRInputS4xD(361)(2) <= CNStageIntLLROutputS4xD(120)(5);
  VNStageIntLLRInputS4xD(21)(2) <= CNStageIntLLROutputS4xD(121)(0);
  VNStageIntLLRInputS4xD(73)(2) <= CNStageIntLLROutputS4xD(121)(1);
  VNStageIntLLRInputS4xD(185)(0) <= CNStageIntLLROutputS4xD(121)(2);
  VNStageIntLLRInputS4xD(253)(1) <= CNStageIntLLROutputS4xD(121)(3);
  VNStageIntLLRInputS4xD(296)(2) <= CNStageIntLLROutputS4xD(121)(4);
  VNStageIntLLRInputS4xD(336)(2) <= CNStageIntLLROutputS4xD(121)(5);
  VNStageIntLLRInputS4xD(19)(2) <= CNStageIntLLROutputS4xD(122)(0);
  VNStageIntLLRInputS4xD(123)(1) <= CNStageIntLLROutputS4xD(122)(1);
  VNStageIntLLRInputS4xD(166)(2) <= CNStageIntLLROutputS4xD(122)(2);
  VNStageIntLLRInputS4xD(206)(1) <= CNStageIntLLROutputS4xD(122)(3);
  VNStageIntLLRInputS4xD(269)(1) <= CNStageIntLLROutputS4xD(122)(4);
  VNStageIntLLRInputS4xD(359)(2) <= CNStageIntLLROutputS4xD(122)(5);
  VNStageIntLLRInputS4xD(18)(2) <= CNStageIntLLROutputS4xD(123)(0);
  VNStageIntLLRInputS4xD(101)(2) <= CNStageIntLLROutputS4xD(123)(1);
  VNStageIntLLRInputS4xD(141)(0) <= CNStageIntLLROutputS4xD(123)(2);
  VNStageIntLLRInputS4xD(204)(2) <= CNStageIntLLROutputS4xD(123)(3);
  VNStageIntLLRInputS4xD(294)(2) <= CNStageIntLLROutputS4xD(123)(4);
  VNStageIntLLRInputS4xD(367)(2) <= CNStageIntLLROutputS4xD(123)(5);
  VNStageIntLLRInputS4xD(17)(2) <= CNStageIntLLROutputS4xD(124)(0);
  VNStageIntLLRInputS4xD(76)(2) <= CNStageIntLLROutputS4xD(124)(1);
  VNStageIntLLRInputS4xD(139)(2) <= CNStageIntLLROutputS4xD(124)(2);
  VNStageIntLLRInputS4xD(229)(2) <= CNStageIntLLROutputS4xD(124)(3);
  VNStageIntLLRInputS4xD(302)(2) <= CNStageIntLLROutputS4xD(124)(4);
  VNStageIntLLRInputS4xD(347)(2) <= CNStageIntLLROutputS4xD(124)(5);
  VNStageIntLLRInputS4xD(16)(1) <= CNStageIntLLROutputS4xD(125)(0);
  VNStageIntLLRInputS4xD(74)(2) <= CNStageIntLLROutputS4xD(125)(1);
  VNStageIntLLRInputS4xD(164)(2) <= CNStageIntLLROutputS4xD(125)(2);
  VNStageIntLLRInputS4xD(237)(2) <= CNStageIntLLROutputS4xD(125)(3);
  VNStageIntLLRInputS4xD(282)(2) <= CNStageIntLLROutputS4xD(125)(4);
  VNStageIntLLRInputS4xD(341)(2) <= CNStageIntLLROutputS4xD(125)(5);
  VNStageIntLLRInputS4xD(15)(2) <= CNStageIntLLROutputS4xD(126)(0);
  VNStageIntLLRInputS4xD(99)(2) <= CNStageIntLLROutputS4xD(126)(1);
  VNStageIntLLRInputS4xD(172)(2) <= CNStageIntLLROutputS4xD(126)(2);
  VNStageIntLLRInputS4xD(217)(2) <= CNStageIntLLROutputS4xD(126)(3);
  VNStageIntLLRInputS4xD(276)(2) <= CNStageIntLLROutputS4xD(126)(4);
  VNStageIntLLRInputS4xD(320)(1) <= CNStageIntLLROutputS4xD(126)(5);
  VNStageIntLLRInputS4xD(14)(2) <= CNStageIntLLROutputS4xD(127)(0);
  VNStageIntLLRInputS4xD(107)(1) <= CNStageIntLLROutputS4xD(127)(1);
  VNStageIntLLRInputS4xD(152)(2) <= CNStageIntLLROutputS4xD(127)(2);
  VNStageIntLLRInputS4xD(211)(2) <= CNStageIntLLROutputS4xD(127)(3);
  VNStageIntLLRInputS4xD(256)(2) <= CNStageIntLLROutputS4xD(127)(4);
  VNStageIntLLRInputS4xD(340)(2) <= CNStageIntLLROutputS4xD(127)(5);
  VNStageIntLLRInputS4xD(13)(1) <= CNStageIntLLROutputS4xD(128)(0);
  VNStageIntLLRInputS4xD(87)(2) <= CNStageIntLLROutputS4xD(128)(1);
  VNStageIntLLRInputS4xD(146)(2) <= CNStageIntLLROutputS4xD(128)(2);
  VNStageIntLLRInputS4xD(192)(2) <= CNStageIntLLROutputS4xD(128)(3);
  VNStageIntLLRInputS4xD(275)(2) <= CNStageIntLLROutputS4xD(128)(4);
  VNStageIntLLRInputS4xD(345)(2) <= CNStageIntLLROutputS4xD(128)(5);
  VNStageIntLLRInputS4xD(12)(2) <= CNStageIntLLROutputS4xD(129)(0);
  VNStageIntLLRInputS4xD(81)(2) <= CNStageIntLLROutputS4xD(129)(1);
  VNStageIntLLRInputS4xD(128)(2) <= CNStageIntLLROutputS4xD(129)(2);
  VNStageIntLLRInputS4xD(210)(2) <= CNStageIntLLROutputS4xD(129)(3);
  VNStageIntLLRInputS4xD(280)(2) <= CNStageIntLLROutputS4xD(129)(4);
  VNStageIntLLRInputS4xD(364)(2) <= CNStageIntLLROutputS4xD(129)(5);
  VNStageIntLLRInputS4xD(11)(2) <= CNStageIntLLROutputS4xD(130)(0);
  VNStageIntLLRInputS4xD(64)(2) <= CNStageIntLLROutputS4xD(130)(1);
  VNStageIntLLRInputS4xD(145)(2) <= CNStageIntLLROutputS4xD(130)(2);
  VNStageIntLLRInputS4xD(215)(2) <= CNStageIntLLROutputS4xD(130)(3);
  VNStageIntLLRInputS4xD(299)(1) <= CNStageIntLLROutputS4xD(130)(4);
  VNStageIntLLRInputS4xD(355)(2) <= CNStageIntLLROutputS4xD(130)(5);
  VNStageIntLLRInputS4xD(10)(2) <= CNStageIntLLROutputS4xD(131)(0);
  VNStageIntLLRInputS4xD(80)(2) <= CNStageIntLLROutputS4xD(131)(1);
  VNStageIntLLRInputS4xD(150)(2) <= CNStageIntLLROutputS4xD(131)(2);
  VNStageIntLLRInputS4xD(234)(2) <= CNStageIntLLROutputS4xD(131)(3);
  VNStageIntLLRInputS4xD(290)(2) <= CNStageIntLLROutputS4xD(131)(4);
  VNStageIntLLRInputS4xD(329)(2) <= CNStageIntLLROutputS4xD(131)(5);
  VNStageIntLLRInputS4xD(9)(2) <= CNStageIntLLROutputS4xD(132)(0);
  VNStageIntLLRInputS4xD(85)(1) <= CNStageIntLLROutputS4xD(132)(1);
  VNStageIntLLRInputS4xD(169)(2) <= CNStageIntLLROutputS4xD(132)(2);
  VNStageIntLLRInputS4xD(225)(2) <= CNStageIntLLROutputS4xD(132)(3);
  VNStageIntLLRInputS4xD(264)(2) <= CNStageIntLLROutputS4xD(132)(4);
  VNStageIntLLRInputS4xD(330)(2) <= CNStageIntLLROutputS4xD(132)(5);
  VNStageIntLLRInputS4xD(8)(1) <= CNStageIntLLROutputS4xD(133)(0);
  VNStageIntLLRInputS4xD(104)(2) <= CNStageIntLLROutputS4xD(133)(1);
  VNStageIntLLRInputS4xD(160)(2) <= CNStageIntLLROutputS4xD(133)(2);
  VNStageIntLLRInputS4xD(199)(2) <= CNStageIntLLROutputS4xD(133)(3);
  VNStageIntLLRInputS4xD(265)(1) <= CNStageIntLLROutputS4xD(133)(4);
  VNStageIntLLRInputS4xD(354)(2) <= CNStageIntLLROutputS4xD(133)(5);
  VNStageIntLLRInputS4xD(7)(2) <= CNStageIntLLROutputS4xD(134)(0);
  VNStageIntLLRInputS4xD(95)(2) <= CNStageIntLLROutputS4xD(134)(1);
  VNStageIntLLRInputS4xD(134)(2) <= CNStageIntLLROutputS4xD(134)(2);
  VNStageIntLLRInputS4xD(200)(2) <= CNStageIntLLROutputS4xD(134)(3);
  VNStageIntLLRInputS4xD(289)(2) <= CNStageIntLLROutputS4xD(134)(4);
  VNStageIntLLRInputS4xD(375)(2) <= CNStageIntLLROutputS4xD(134)(5);
  VNStageIntLLRInputS4xD(6)(2) <= CNStageIntLLROutputS4xD(135)(0);
  VNStageIntLLRInputS4xD(69)(2) <= CNStageIntLLROutputS4xD(135)(1);
  VNStageIntLLRInputS4xD(135)(2) <= CNStageIntLLROutputS4xD(135)(2);
  VNStageIntLLRInputS4xD(224)(2) <= CNStageIntLLROutputS4xD(135)(3);
  VNStageIntLLRInputS4xD(310)(2) <= CNStageIntLLROutputS4xD(135)(4);
  VNStageIntLLRInputS4xD(371)(1) <= CNStageIntLLROutputS4xD(135)(5);
  VNStageIntLLRInputS4xD(5)(2) <= CNStageIntLLROutputS4xD(136)(0);
  VNStageIntLLRInputS4xD(70)(2) <= CNStageIntLLROutputS4xD(136)(1);
  VNStageIntLLRInputS4xD(159)(2) <= CNStageIntLLROutputS4xD(136)(2);
  VNStageIntLLRInputS4xD(245)(2) <= CNStageIntLLROutputS4xD(136)(3);
  VNStageIntLLRInputS4xD(306)(2) <= CNStageIntLLROutputS4xD(136)(4);
  VNStageIntLLRInputS4xD(323)(1) <= CNStageIntLLROutputS4xD(136)(5);
  VNStageIntLLRInputS4xD(3)(1) <= CNStageIntLLROutputS4xD(137)(0);
  VNStageIntLLRInputS4xD(115)(2) <= CNStageIntLLROutputS4xD(137)(1);
  VNStageIntLLRInputS4xD(176)(2) <= CNStageIntLLROutputS4xD(137)(2);
  VNStageIntLLRInputS4xD(193)(2) <= CNStageIntLLROutputS4xD(137)(3);
  VNStageIntLLRInputS4xD(284)(2) <= CNStageIntLLROutputS4xD(137)(4);
  VNStageIntLLRInputS4xD(325)(2) <= CNStageIntLLROutputS4xD(137)(5);
  VNStageIntLLRInputS4xD(2)(2) <= CNStageIntLLROutputS4xD(138)(0);
  VNStageIntLLRInputS4xD(111)(2) <= CNStageIntLLROutputS4xD(138)(1);
  VNStageIntLLRInputS4xD(191)(2) <= CNStageIntLLROutputS4xD(138)(2);
  VNStageIntLLRInputS4xD(219)(2) <= CNStageIntLLROutputS4xD(138)(3);
  VNStageIntLLRInputS4xD(260)(2) <= CNStageIntLLROutputS4xD(138)(4);
  VNStageIntLLRInputS4xD(357)(2) <= CNStageIntLLROutputS4xD(138)(5);
  VNStageIntLLRInputS4xD(1)(1) <= CNStageIntLLROutputS4xD(139)(0);
  VNStageIntLLRInputS4xD(126)(1) <= CNStageIntLLROutputS4xD(139)(1);
  VNStageIntLLRInputS4xD(154)(1) <= CNStageIntLLROutputS4xD(139)(2);
  VNStageIntLLRInputS4xD(195)(1) <= CNStageIntLLROutputS4xD(139)(3);
  VNStageIntLLRInputS4xD(292)(2) <= CNStageIntLLROutputS4xD(139)(4);
  VNStageIntLLRInputS4xD(373)(1) <= CNStageIntLLROutputS4xD(139)(5);
  VNStageIntLLRInputS4xD(63)(2) <= CNStageIntLLROutputS4xD(140)(0);
  VNStageIntLLRInputS4xD(89)(2) <= CNStageIntLLROutputS4xD(140)(1);
  VNStageIntLLRInputS4xD(130)(2) <= CNStageIntLLROutputS4xD(140)(2);
  VNStageIntLLRInputS4xD(227)(2) <= CNStageIntLLROutputS4xD(140)(3);
  VNStageIntLLRInputS4xD(308)(0) <= CNStageIntLLROutputS4xD(140)(4);
  VNStageIntLLRInputS4xD(343)(2) <= CNStageIntLLROutputS4xD(140)(5);
  VNStageIntLLRInputS4xD(62)(1) <= CNStageIntLLROutputS4xD(141)(0);
  VNStageIntLLRInputS4xD(65)(2) <= CNStageIntLLROutputS4xD(141)(1);
  VNStageIntLLRInputS4xD(162)(2) <= CNStageIntLLROutputS4xD(141)(2);
  VNStageIntLLRInputS4xD(243)(2) <= CNStageIntLLROutputS4xD(141)(3);
  VNStageIntLLRInputS4xD(278)(2) <= CNStageIntLLROutputS4xD(141)(4);
  VNStageIntLLRInputS4xD(352)(2) <= CNStageIntLLROutputS4xD(141)(5);
  VNStageIntLLRInputS4xD(61)(1) <= CNStageIntLLROutputS4xD(142)(0);
  VNStageIntLLRInputS4xD(97)(2) <= CNStageIntLLROutputS4xD(142)(1);
  VNStageIntLLRInputS4xD(178)(2) <= CNStageIntLLROutputS4xD(142)(2);
  VNStageIntLLRInputS4xD(213)(2) <= CNStageIntLLROutputS4xD(142)(3);
  VNStageIntLLRInputS4xD(287)(2) <= CNStageIntLLROutputS4xD(142)(4);
  VNStageIntLLRInputS4xD(365)(2) <= CNStageIntLLROutputS4xD(142)(5);
  VNStageIntLLRInputS4xD(60)(1) <= CNStageIntLLROutputS4xD(143)(0);
  VNStageIntLLRInputS4xD(113)(2) <= CNStageIntLLROutputS4xD(143)(1);
  VNStageIntLLRInputS4xD(148)(2) <= CNStageIntLLROutputS4xD(143)(2);
  VNStageIntLLRInputS4xD(222)(1) <= CNStageIntLLROutputS4xD(143)(3);
  VNStageIntLLRInputS4xD(300)(2) <= CNStageIntLLROutputS4xD(143)(4);
  VNStageIntLLRInputS4xD(344)(2) <= CNStageIntLLROutputS4xD(143)(5);
  VNStageIntLLRInputS4xD(59)(0) <= CNStageIntLLROutputS4xD(144)(0);
  VNStageIntLLRInputS4xD(83)(2) <= CNStageIntLLROutputS4xD(144)(1);
  VNStageIntLLRInputS4xD(157)(2) <= CNStageIntLLROutputS4xD(144)(2);
  VNStageIntLLRInputS4xD(235)(1) <= CNStageIntLLROutputS4xD(144)(3);
  VNStageIntLLRInputS4xD(279)(2) <= CNStageIntLLROutputS4xD(144)(4);
  VNStageIntLLRInputS4xD(372)(1) <= CNStageIntLLROutputS4xD(144)(5);
  VNStageIntLLRInputS4xD(58)(1) <= CNStageIntLLROutputS4xD(145)(0);
  VNStageIntLLRInputS4xD(92)(2) <= CNStageIntLLROutputS4xD(145)(1);
  VNStageIntLLRInputS4xD(170)(2) <= CNStageIntLLROutputS4xD(145)(2);
  VNStageIntLLRInputS4xD(214)(2) <= CNStageIntLLROutputS4xD(145)(3);
  VNStageIntLLRInputS4xD(307)(2) <= CNStageIntLLROutputS4xD(145)(4);
  VNStageIntLLRInputS4xD(374)(2) <= CNStageIntLLROutputS4xD(145)(5);
  VNStageIntLLRInputS4xD(57)(1) <= CNStageIntLLROutputS4xD(146)(0);
  VNStageIntLLRInputS4xD(105)(1) <= CNStageIntLLROutputS4xD(146)(1);
  VNStageIntLLRInputS4xD(149)(2) <= CNStageIntLLROutputS4xD(146)(2);
  VNStageIntLLRInputS4xD(242)(2) <= CNStageIntLLROutputS4xD(146)(3);
  VNStageIntLLRInputS4xD(309)(2) <= CNStageIntLLROutputS4xD(146)(4);
  VNStageIntLLRInputS4xD(356)(2) <= CNStageIntLLROutputS4xD(146)(5);
  VNStageIntLLRInputS4xD(56)(2) <= CNStageIntLLROutputS4xD(147)(0);
  VNStageIntLLRInputS4xD(84)(2) <= CNStageIntLLROutputS4xD(147)(1);
  VNStageIntLLRInputS4xD(177)(2) <= CNStageIntLLROutputS4xD(147)(2);
  VNStageIntLLRInputS4xD(244)(0) <= CNStageIntLLROutputS4xD(147)(3);
  VNStageIntLLRInputS4xD(291)(2) <= CNStageIntLLROutputS4xD(147)(4);
  VNStageIntLLRInputS4xD(363)(1) <= CNStageIntLLROutputS4xD(147)(5);
  VNStageIntLLRInputS4xD(55)(2) <= CNStageIntLLROutputS4xD(148)(0);
  VNStageIntLLRInputS4xD(112)(2) <= CNStageIntLLROutputS4xD(148)(1);
  VNStageIntLLRInputS4xD(179)(2) <= CNStageIntLLROutputS4xD(148)(2);
  VNStageIntLLRInputS4xD(226)(1) <= CNStageIntLLROutputS4xD(148)(3);
  VNStageIntLLRInputS4xD(298)(2) <= CNStageIntLLROutputS4xD(148)(4);
  VNStageIntLLRInputS4xD(327)(2) <= CNStageIntLLROutputS4xD(148)(5);
  VNStageIntLLRInputS4xD(54)(2) <= CNStageIntLLROutputS4xD(149)(0);
  VNStageIntLLRInputS4xD(114)(2) <= CNStageIntLLROutputS4xD(149)(1);
  VNStageIntLLRInputS4xD(161)(2) <= CNStageIntLLROutputS4xD(149)(2);
  VNStageIntLLRInputS4xD(233)(2) <= CNStageIntLLROutputS4xD(149)(3);
  VNStageIntLLRInputS4xD(262)(2) <= CNStageIntLLROutputS4xD(149)(4);
  VNStageIntLLRInputS4xD(378)(1) <= CNStageIntLLROutputS4xD(149)(5);
  VNStageIntLLRInputS4xD(53)(1) <= CNStageIntLLROutputS4xD(150)(0);
  VNStageIntLLRInputS4xD(96)(2) <= CNStageIntLLROutputS4xD(150)(1);
  VNStageIntLLRInputS4xD(168)(1) <= CNStageIntLLROutputS4xD(150)(2);
  VNStageIntLLRInputS4xD(197)(2) <= CNStageIntLLROutputS4xD(150)(3);
  VNStageIntLLRInputS4xD(313)(0) <= CNStageIntLLROutputS4xD(150)(4);
  VNStageIntLLRInputS4xD(321)(2) <= CNStageIntLLROutputS4xD(150)(5);
  VNStageIntLLRInputS4xD(52)(1) <= CNStageIntLLROutputS4xD(151)(0);
  VNStageIntLLRInputS4xD(103)(2) <= CNStageIntLLROutputS4xD(151)(1);
  VNStageIntLLRInputS4xD(132)(1) <= CNStageIntLLROutputS4xD(151)(2);
  VNStageIntLLRInputS4xD(248)(2) <= CNStageIntLLROutputS4xD(151)(3);
  VNStageIntLLRInputS4xD(319)(2) <= CNStageIntLLROutputS4xD(151)(4);
  VNStageIntLLRInputS4xD(379)(1) <= CNStageIntLLROutputS4xD(151)(5);
  VNStageIntLLRInputS4xD(50)(2) <= CNStageIntLLROutputS4xD(152)(0);
  VNStageIntLLRInputS4xD(118)(2) <= CNStageIntLLROutputS4xD(152)(1);
  VNStageIntLLRInputS4xD(189)(1) <= CNStageIntLLROutputS4xD(152)(2);
  VNStageIntLLRInputS4xD(249)(0) <= CNStageIntLLROutputS4xD(152)(3);
  VNStageIntLLRInputS4xD(261)(2) <= CNStageIntLLROutputS4xD(152)(4);
  VNStageIntLLRInputS4xD(348)(2) <= CNStageIntLLROutputS4xD(152)(5);
  VNStageIntLLRInputS4xD(49)(2) <= CNStageIntLLROutputS4xD(153)(0);
  VNStageIntLLRInputS4xD(124)(1) <= CNStageIntLLROutputS4xD(153)(1);
  VNStageIntLLRInputS4xD(184)(2) <= CNStageIntLLROutputS4xD(153)(2);
  VNStageIntLLRInputS4xD(196)(2) <= CNStageIntLLROutputS4xD(153)(3);
  VNStageIntLLRInputS4xD(283)(2) <= CNStageIntLLROutputS4xD(153)(4);
  VNStageIntLLRInputS4xD(366)(2) <= CNStageIntLLROutputS4xD(153)(5);
  VNStageIntLLRInputS4xD(48)(1) <= CNStageIntLLROutputS4xD(154)(0);
  VNStageIntLLRInputS4xD(119)(2) <= CNStageIntLLROutputS4xD(154)(1);
  VNStageIntLLRInputS4xD(131)(1) <= CNStageIntLLROutputS4xD(154)(2);
  VNStageIntLLRInputS4xD(218)(2) <= CNStageIntLLROutputS4xD(154)(3);
  VNStageIntLLRInputS4xD(301)(2) <= CNStageIntLLROutputS4xD(154)(4);
  VNStageIntLLRInputS4xD(351)(1) <= CNStageIntLLROutputS4xD(154)(5);
  VNStageIntLLRInputS4xD(47)(1) <= CNStageIntLLROutputS4xD(155)(0);
  VNStageIntLLRInputS4xD(66)(2) <= CNStageIntLLROutputS4xD(155)(1);
  VNStageIntLLRInputS4xD(153)(2) <= CNStageIntLLROutputS4xD(155)(2);
  VNStageIntLLRInputS4xD(236)(2) <= CNStageIntLLROutputS4xD(155)(3);
  VNStageIntLLRInputS4xD(286)(2) <= CNStageIntLLROutputS4xD(155)(4);
  VNStageIntLLRInputS4xD(338)(2) <= CNStageIntLLROutputS4xD(155)(5);
  VNStageIntLLRInputS4xD(46)(2) <= CNStageIntLLROutputS4xD(156)(0);
  VNStageIntLLRInputS4xD(88)(2) <= CNStageIntLLROutputS4xD(156)(1);
  VNStageIntLLRInputS4xD(171)(1) <= CNStageIntLLROutputS4xD(156)(2);
  VNStageIntLLRInputS4xD(221)(2) <= CNStageIntLLROutputS4xD(156)(3);
  VNStageIntLLRInputS4xD(273)(2) <= CNStageIntLLROutputS4xD(156)(4);
  VNStageIntLLRInputS4xD(369)(1) <= CNStageIntLLROutputS4xD(156)(5);
  VNStageIntLLRInputS4xD(45)(2) <= CNStageIntLLROutputS4xD(157)(0);
  VNStageIntLLRInputS4xD(106)(1) <= CNStageIntLLROutputS4xD(157)(1);
  VNStageIntLLRInputS4xD(156)(2) <= CNStageIntLLROutputS4xD(157)(2);
  VNStageIntLLRInputS4xD(208)(2) <= CNStageIntLLROutputS4xD(157)(3);
  VNStageIntLLRInputS4xD(304)(2) <= CNStageIntLLROutputS4xD(157)(4);
  VNStageIntLLRInputS4xD(381)(1) <= CNStageIntLLROutputS4xD(157)(5);
  VNStageIntLLRInputS4xD(44)(2) <= CNStageIntLLROutputS4xD(158)(0);
  VNStageIntLLRInputS4xD(91)(2) <= CNStageIntLLROutputS4xD(158)(1);
  VNStageIntLLRInputS4xD(143)(2) <= CNStageIntLLROutputS4xD(158)(2);
  VNStageIntLLRInputS4xD(239)(2) <= CNStageIntLLROutputS4xD(158)(3);
  VNStageIntLLRInputS4xD(316)(1) <= CNStageIntLLROutputS4xD(158)(4);
  VNStageIntLLRInputS4xD(332)(2) <= CNStageIntLLROutputS4xD(158)(5);
  VNStageIntLLRInputS4xD(43)(1) <= CNStageIntLLROutputS4xD(159)(0);
  VNStageIntLLRInputS4xD(78)(2) <= CNStageIntLLROutputS4xD(159)(1);
  VNStageIntLLRInputS4xD(174)(2) <= CNStageIntLLROutputS4xD(159)(2);
  VNStageIntLLRInputS4xD(251)(1) <= CNStageIntLLROutputS4xD(159)(3);
  VNStageIntLLRInputS4xD(267)(2) <= CNStageIntLLROutputS4xD(159)(4);
  VNStageIntLLRInputS4xD(376)(2) <= CNStageIntLLROutputS4xD(159)(5);
  VNStageIntLLRInputS4xD(42)(2) <= CNStageIntLLROutputS4xD(160)(0);
  VNStageIntLLRInputS4xD(109)(2) <= CNStageIntLLROutputS4xD(160)(1);
  VNStageIntLLRInputS4xD(186)(1) <= CNStageIntLLROutputS4xD(160)(2);
  VNStageIntLLRInputS4xD(202)(2) <= CNStageIntLLROutputS4xD(160)(3);
  VNStageIntLLRInputS4xD(311)(2) <= CNStageIntLLROutputS4xD(160)(4);
  VNStageIntLLRInputS4xD(353)(2) <= CNStageIntLLROutputS4xD(160)(5);
  VNStageIntLLRInputS4xD(41)(2) <= CNStageIntLLROutputS4xD(161)(0);
  VNStageIntLLRInputS4xD(121)(1) <= CNStageIntLLROutputS4xD(161)(1);
  VNStageIntLLRInputS4xD(137)(2) <= CNStageIntLLROutputS4xD(161)(2);
  VNStageIntLLRInputS4xD(246)(2) <= CNStageIntLLROutputS4xD(161)(3);
  VNStageIntLLRInputS4xD(288)(2) <= CNStageIntLLROutputS4xD(161)(4);
  VNStageIntLLRInputS4xD(342)(2) <= CNStageIntLLROutputS4xD(161)(5);
  VNStageIntLLRInputS4xD(40)(2) <= CNStageIntLLROutputS4xD(162)(0);
  VNStageIntLLRInputS4xD(72)(2) <= CNStageIntLLROutputS4xD(162)(1);
  VNStageIntLLRInputS4xD(181)(2) <= CNStageIntLLROutputS4xD(162)(2);
  VNStageIntLLRInputS4xD(223)(2) <= CNStageIntLLROutputS4xD(162)(3);
  VNStageIntLLRInputS4xD(277)(2) <= CNStageIntLLROutputS4xD(162)(4);
  VNStageIntLLRInputS4xD(346)(2) <= CNStageIntLLROutputS4xD(162)(5);
  VNStageIntLLRInputS4xD(39)(2) <= CNStageIntLLROutputS4xD(163)(0);
  VNStageIntLLRInputS4xD(116)(1) <= CNStageIntLLROutputS4xD(163)(1);
  VNStageIntLLRInputS4xD(158)(2) <= CNStageIntLLROutputS4xD(163)(2);
  VNStageIntLLRInputS4xD(212)(2) <= CNStageIntLLROutputS4xD(163)(3);
  VNStageIntLLRInputS4xD(281)(2) <= CNStageIntLLROutputS4xD(163)(4);
  VNStageIntLLRInputS4xD(339)(2) <= CNStageIntLLROutputS4xD(163)(5);
  VNStageIntLLRInputS4xD(38)(2) <= CNStageIntLLROutputS4xD(164)(0);
  VNStageIntLLRInputS4xD(93)(2) <= CNStageIntLLROutputS4xD(164)(1);
  VNStageIntLLRInputS4xD(147)(2) <= CNStageIntLLROutputS4xD(164)(2);
  VNStageIntLLRInputS4xD(216)(2) <= CNStageIntLLROutputS4xD(164)(3);
  VNStageIntLLRInputS4xD(274)(1) <= CNStageIntLLROutputS4xD(164)(4);
  VNStageIntLLRInputS4xD(350)(2) <= CNStageIntLLROutputS4xD(164)(5);
  VNStageIntLLRInputS4xD(37)(2) <= CNStageIntLLROutputS4xD(165)(0);
  VNStageIntLLRInputS4xD(82)(2) <= CNStageIntLLROutputS4xD(165)(1);
  VNStageIntLLRInputS4xD(151)(2) <= CNStageIntLLROutputS4xD(165)(2);
  VNStageIntLLRInputS4xD(209)(2) <= CNStageIntLLROutputS4xD(165)(3);
  VNStageIntLLRInputS4xD(285)(2) <= CNStageIntLLROutputS4xD(165)(4);
  VNStageIntLLRInputS4xD(322)(2) <= CNStageIntLLROutputS4xD(165)(5);
  VNStageIntLLRInputS4xD(36)(2) <= CNStageIntLLROutputS4xD(166)(0);
  VNStageIntLLRInputS4xD(86)(1) <= CNStageIntLLROutputS4xD(166)(1);
  VNStageIntLLRInputS4xD(144)(2) <= CNStageIntLLROutputS4xD(166)(2);
  VNStageIntLLRInputS4xD(220)(2) <= CNStageIntLLROutputS4xD(166)(3);
  VNStageIntLLRInputS4xD(257)(2) <= CNStageIntLLROutputS4xD(166)(4);
  VNStageIntLLRInputS4xD(377)(1) <= CNStageIntLLROutputS4xD(166)(5);
  VNStageIntLLRInputS4xD(35)(2) <= CNStageIntLLROutputS4xD(167)(0);
  VNStageIntLLRInputS4xD(79)(2) <= CNStageIntLLROutputS4xD(167)(1);
  VNStageIntLLRInputS4xD(155)(2) <= CNStageIntLLROutputS4xD(167)(2);
  VNStageIntLLRInputS4xD(255)(2) <= CNStageIntLLROutputS4xD(167)(3);
  VNStageIntLLRInputS4xD(312)(2) <= CNStageIntLLROutputS4xD(167)(4);
  VNStageIntLLRInputS4xD(331)(2) <= CNStageIntLLROutputS4xD(167)(5);
  VNStageIntLLRInputS4xD(34)(2) <= CNStageIntLLROutputS4xD(168)(0);
  VNStageIntLLRInputS4xD(90)(2) <= CNStageIntLLROutputS4xD(168)(1);
  VNStageIntLLRInputS4xD(190)(0) <= CNStageIntLLROutputS4xD(168)(2);
  VNStageIntLLRInputS4xD(247)(2) <= CNStageIntLLROutputS4xD(168)(3);
  VNStageIntLLRInputS4xD(266)(1) <= CNStageIntLLROutputS4xD(168)(4);
  VNStageIntLLRInputS4xD(328)(2) <= CNStageIntLLROutputS4xD(168)(5);
  VNStageIntLLRInputS4xD(33)(2) <= CNStageIntLLROutputS4xD(169)(0);
  VNStageIntLLRInputS4xD(125)(1) <= CNStageIntLLROutputS4xD(169)(1);
  VNStageIntLLRInputS4xD(182)(2) <= CNStageIntLLROutputS4xD(169)(2);
  VNStageIntLLRInputS4xD(201)(2) <= CNStageIntLLROutputS4xD(169)(3);
  VNStageIntLLRInputS4xD(263)(2) <= CNStageIntLLROutputS4xD(169)(4);
  VNStageIntLLRInputS4xD(362)(2) <= CNStageIntLLROutputS4xD(169)(5);
  VNStageIntLLRInputS4xD(0)(2) <= CNStageIntLLROutputS4xD(170)(0);
  VNStageIntLLRInputS4xD(75)(2) <= CNStageIntLLROutputS4xD(170)(1);
  VNStageIntLLRInputS4xD(140)(2) <= CNStageIntLLROutputS4xD(170)(2);
  VNStageIntLLRInputS4xD(205)(0) <= CNStageIntLLROutputS4xD(170)(3);
  VNStageIntLLRInputS4xD(270)(2) <= CNStageIntLLROutputS4xD(170)(4);
  VNStageIntLLRInputS4xD(335)(2) <= CNStageIntLLROutputS4xD(170)(5);
  VNStageIntLLRInputS4xD(62)(2) <= CNStageIntLLROutputS4xD(171)(0);
  VNStageIntLLRInputS4xD(109)(3) <= CNStageIntLLROutputS4xD(171)(1);
  VNStageIntLLRInputS4xD(161)(3) <= CNStageIntLLROutputS4xD(171)(2);
  VNStageIntLLRInputS4xD(194)(3) <= CNStageIntLLROutputS4xD(171)(3);
  VNStageIntLLRInputS4xD(271)(2) <= CNStageIntLLROutputS4xD(171)(4);
  VNStageIntLLRInputS4xD(350)(3) <= CNStageIntLLROutputS4xD(171)(5);
  VNStageIntLLRInputS4xD(61)(2) <= CNStageIntLLROutputS4xD(172)(0);
  VNStageIntLLRInputS4xD(96)(3) <= CNStageIntLLROutputS4xD(172)(1);
  VNStageIntLLRInputS4xD(129)(3) <= CNStageIntLLROutputS4xD(172)(2);
  VNStageIntLLRInputS4xD(206)(2) <= CNStageIntLLROutputS4xD(172)(3);
  VNStageIntLLRInputS4xD(285)(3) <= CNStageIntLLROutputS4xD(172)(4);
  VNStageIntLLRInputS4xD(331)(3) <= CNStageIntLLROutputS4xD(172)(5);
  VNStageIntLLRInputS4xD(60)(2) <= CNStageIntLLROutputS4xD(173)(0);
  VNStageIntLLRInputS4xD(127)(3) <= CNStageIntLLROutputS4xD(173)(1);
  VNStageIntLLRInputS4xD(141)(1) <= CNStageIntLLROutputS4xD(173)(2);
  VNStageIntLLRInputS4xD(220)(3) <= CNStageIntLLROutputS4xD(173)(3);
  VNStageIntLLRInputS4xD(266)(2) <= CNStageIntLLROutputS4xD(173)(4);
  VNStageIntLLRInputS4xD(371)(2) <= CNStageIntLLROutputS4xD(173)(5);
  VNStageIntLLRInputS4xD(59)(1) <= CNStageIntLLROutputS4xD(174)(0);
  VNStageIntLLRInputS4xD(76)(3) <= CNStageIntLLROutputS4xD(174)(1);
  VNStageIntLLRInputS4xD(155)(3) <= CNStageIntLLROutputS4xD(174)(2);
  VNStageIntLLRInputS4xD(201)(3) <= CNStageIntLLROutputS4xD(174)(3);
  VNStageIntLLRInputS4xD(306)(3) <= CNStageIntLLROutputS4xD(174)(4);
  VNStageIntLLRInputS4xD(360)(3) <= CNStageIntLLROutputS4xD(174)(5);
  VNStageIntLLRInputS4xD(58)(2) <= CNStageIntLLROutputS4xD(175)(0);
  VNStageIntLLRInputS4xD(90)(3) <= CNStageIntLLROutputS4xD(175)(1);
  VNStageIntLLRInputS4xD(136)(3) <= CNStageIntLLROutputS4xD(175)(2);
  VNStageIntLLRInputS4xD(241)(2) <= CNStageIntLLROutputS4xD(175)(3);
  VNStageIntLLRInputS4xD(295)(3) <= CNStageIntLLROutputS4xD(175)(4);
  VNStageIntLLRInputS4xD(364)(3) <= CNStageIntLLROutputS4xD(175)(5);
  VNStageIntLLRInputS4xD(57)(2) <= CNStageIntLLROutputS4xD(176)(0);
  VNStageIntLLRInputS4xD(71)(2) <= CNStageIntLLROutputS4xD(176)(1);
  VNStageIntLLRInputS4xD(176)(3) <= CNStageIntLLROutputS4xD(176)(2);
  VNStageIntLLRInputS4xD(230)(2) <= CNStageIntLLROutputS4xD(176)(3);
  VNStageIntLLRInputS4xD(299)(2) <= CNStageIntLLROutputS4xD(176)(4);
  VNStageIntLLRInputS4xD(357)(3) <= CNStageIntLLROutputS4xD(176)(5);
  VNStageIntLLRInputS4xD(56)(3) <= CNStageIntLLROutputS4xD(177)(0);
  VNStageIntLLRInputS4xD(111)(3) <= CNStageIntLLROutputS4xD(177)(1);
  VNStageIntLLRInputS4xD(165)(3) <= CNStageIntLLROutputS4xD(177)(2);
  VNStageIntLLRInputS4xD(234)(3) <= CNStageIntLLROutputS4xD(177)(3);
  VNStageIntLLRInputS4xD(292)(3) <= CNStageIntLLROutputS4xD(177)(4);
  VNStageIntLLRInputS4xD(368)(1) <= CNStageIntLLROutputS4xD(177)(5);
  VNStageIntLLRInputS4xD(55)(3) <= CNStageIntLLROutputS4xD(178)(0);
  VNStageIntLLRInputS4xD(100)(3) <= CNStageIntLLROutputS4xD(178)(1);
  VNStageIntLLRInputS4xD(169)(3) <= CNStageIntLLROutputS4xD(178)(2);
  VNStageIntLLRInputS4xD(227)(3) <= CNStageIntLLROutputS4xD(178)(3);
  VNStageIntLLRInputS4xD(303)(3) <= CNStageIntLLROutputS4xD(178)(4);
  VNStageIntLLRInputS4xD(340)(3) <= CNStageIntLLROutputS4xD(178)(5);
  VNStageIntLLRInputS4xD(54)(3) <= CNStageIntLLROutputS4xD(179)(0);
  VNStageIntLLRInputS4xD(104)(3) <= CNStageIntLLROutputS4xD(179)(1);
  VNStageIntLLRInputS4xD(162)(3) <= CNStageIntLLROutputS4xD(179)(2);
  VNStageIntLLRInputS4xD(238)(3) <= CNStageIntLLROutputS4xD(179)(3);
  VNStageIntLLRInputS4xD(275)(3) <= CNStageIntLLROutputS4xD(179)(4);
  VNStageIntLLRInputS4xD(332)(3) <= CNStageIntLLROutputS4xD(179)(5);
  VNStageIntLLRInputS4xD(53)(2) <= CNStageIntLLROutputS4xD(180)(0);
  VNStageIntLLRInputS4xD(97)(3) <= CNStageIntLLROutputS4xD(180)(1);
  VNStageIntLLRInputS4xD(173)(3) <= CNStageIntLLROutputS4xD(180)(2);
  VNStageIntLLRInputS4xD(210)(3) <= CNStageIntLLROutputS4xD(180)(3);
  VNStageIntLLRInputS4xD(267)(3) <= CNStageIntLLROutputS4xD(180)(4);
  VNStageIntLLRInputS4xD(349)(2) <= CNStageIntLLROutputS4xD(180)(5);
  VNStageIntLLRInputS4xD(52)(2) <= CNStageIntLLROutputS4xD(181)(0);
  VNStageIntLLRInputS4xD(108)(3) <= CNStageIntLLROutputS4xD(181)(1);
  VNStageIntLLRInputS4xD(145)(3) <= CNStageIntLLROutputS4xD(181)(2);
  VNStageIntLLRInputS4xD(202)(3) <= CNStageIntLLROutputS4xD(181)(3);
  VNStageIntLLRInputS4xD(284)(3) <= CNStageIntLLROutputS4xD(181)(4);
  VNStageIntLLRInputS4xD(346)(3) <= CNStageIntLLROutputS4xD(181)(5);
  VNStageIntLLRInputS4xD(51)(2) <= CNStageIntLLROutputS4xD(182)(0);
  VNStageIntLLRInputS4xD(80)(3) <= CNStageIntLLROutputS4xD(182)(1);
  VNStageIntLLRInputS4xD(137)(3) <= CNStageIntLLROutputS4xD(182)(2);
  VNStageIntLLRInputS4xD(219)(3) <= CNStageIntLLROutputS4xD(182)(3);
  VNStageIntLLRInputS4xD(281)(3) <= CNStageIntLLROutputS4xD(182)(4);
  VNStageIntLLRInputS4xD(380)(2) <= CNStageIntLLROutputS4xD(182)(5);
  VNStageIntLLRInputS4xD(50)(3) <= CNStageIntLLROutputS4xD(183)(0);
  VNStageIntLLRInputS4xD(72)(3) <= CNStageIntLLROutputS4xD(183)(1);
  VNStageIntLLRInputS4xD(154)(2) <= CNStageIntLLROutputS4xD(183)(2);
  VNStageIntLLRInputS4xD(216)(3) <= CNStageIntLLROutputS4xD(183)(3);
  VNStageIntLLRInputS4xD(315)(2) <= CNStageIntLLROutputS4xD(183)(4);
  VNStageIntLLRInputS4xD(337)(3) <= CNStageIntLLROutputS4xD(183)(5);
  VNStageIntLLRInputS4xD(49)(3) <= CNStageIntLLROutputS4xD(184)(0);
  VNStageIntLLRInputS4xD(89)(3) <= CNStageIntLLROutputS4xD(184)(1);
  VNStageIntLLRInputS4xD(151)(3) <= CNStageIntLLROutputS4xD(184)(2);
  VNStageIntLLRInputS4xD(250)(2) <= CNStageIntLLROutputS4xD(184)(3);
  VNStageIntLLRInputS4xD(272)(3) <= CNStageIntLLROutputS4xD(184)(4);
  VNStageIntLLRInputS4xD(323)(2) <= CNStageIntLLROutputS4xD(184)(5);
  VNStageIntLLRInputS4xD(46)(3) <= CNStageIntLLROutputS4xD(185)(0);
  VNStageIntLLRInputS4xD(77)(1) <= CNStageIntLLROutputS4xD(185)(1);
  VNStageIntLLRInputS4xD(191)(3) <= CNStageIntLLROutputS4xD(185)(2);
  VNStageIntLLRInputS4xD(246)(3) <= CNStageIntLLROutputS4xD(185)(3);
  VNStageIntLLRInputS4xD(277)(3) <= CNStageIntLLROutputS4xD(185)(4);
  VNStageIntLLRInputS4xD(325)(3) <= CNStageIntLLROutputS4xD(185)(5);
  VNStageIntLLRInputS4xD(45)(3) <= CNStageIntLLROutputS4xD(186)(0);
  VNStageIntLLRInputS4xD(126)(2) <= CNStageIntLLROutputS4xD(186)(1);
  VNStageIntLLRInputS4xD(181)(3) <= CNStageIntLLROutputS4xD(186)(2);
  VNStageIntLLRInputS4xD(212)(3) <= CNStageIntLLROutputS4xD(186)(3);
  VNStageIntLLRInputS4xD(260)(3) <= CNStageIntLLROutputS4xD(186)(4);
  VNStageIntLLRInputS4xD(355)(3) <= CNStageIntLLROutputS4xD(186)(5);
  VNStageIntLLRInputS4xD(44)(3) <= CNStageIntLLROutputS4xD(187)(0);
  VNStageIntLLRInputS4xD(116)(2) <= CNStageIntLLROutputS4xD(187)(1);
  VNStageIntLLRInputS4xD(147)(3) <= CNStageIntLLROutputS4xD(187)(2);
  VNStageIntLLRInputS4xD(195)(2) <= CNStageIntLLROutputS4xD(187)(3);
  VNStageIntLLRInputS4xD(290)(3) <= CNStageIntLLROutputS4xD(187)(4);
  VNStageIntLLRInputS4xD(378)(2) <= CNStageIntLLROutputS4xD(187)(5);
  VNStageIntLLRInputS4xD(43)(2) <= CNStageIntLLROutputS4xD(188)(0);
  VNStageIntLLRInputS4xD(82)(3) <= CNStageIntLLROutputS4xD(188)(1);
  VNStageIntLLRInputS4xD(130)(3) <= CNStageIntLLROutputS4xD(188)(2);
  VNStageIntLLRInputS4xD(225)(3) <= CNStageIntLLROutputS4xD(188)(3);
  VNStageIntLLRInputS4xD(313)(1) <= CNStageIntLLROutputS4xD(188)(4);
  VNStageIntLLRInputS4xD(351)(2) <= CNStageIntLLROutputS4xD(188)(5);
  VNStageIntLLRInputS4xD(42)(3) <= CNStageIntLLROutputS4xD(189)(0);
  VNStageIntLLRInputS4xD(65)(3) <= CNStageIntLLROutputS4xD(189)(1);
  VNStageIntLLRInputS4xD(160)(3) <= CNStageIntLLROutputS4xD(189)(2);
  VNStageIntLLRInputS4xD(248)(3) <= CNStageIntLLROutputS4xD(189)(3);
  VNStageIntLLRInputS4xD(286)(3) <= CNStageIntLLROutputS4xD(189)(4);
  VNStageIntLLRInputS4xD(335)(3) <= CNStageIntLLROutputS4xD(189)(5);
  VNStageIntLLRInputS4xD(41)(3) <= CNStageIntLLROutputS4xD(190)(0);
  VNStageIntLLRInputS4xD(95)(3) <= CNStageIntLLROutputS4xD(190)(1);
  VNStageIntLLRInputS4xD(183)(2) <= CNStageIntLLROutputS4xD(190)(2);
  VNStageIntLLRInputS4xD(221)(3) <= CNStageIntLLROutputS4xD(190)(3);
  VNStageIntLLRInputS4xD(270)(3) <= CNStageIntLLROutputS4xD(190)(4);
  VNStageIntLLRInputS4xD(338)(3) <= CNStageIntLLROutputS4xD(190)(5);
  VNStageIntLLRInputS4xD(39)(3) <= CNStageIntLLROutputS4xD(191)(0);
  VNStageIntLLRInputS4xD(91)(3) <= CNStageIntLLROutputS4xD(191)(1);
  VNStageIntLLRInputS4xD(140)(3) <= CNStageIntLLROutputS4xD(191)(2);
  VNStageIntLLRInputS4xD(208)(3) <= CNStageIntLLROutputS4xD(191)(3);
  VNStageIntLLRInputS4xD(314)(0) <= CNStageIntLLROutputS4xD(191)(4);
  VNStageIntLLRInputS4xD(354)(3) <= CNStageIntLLROutputS4xD(191)(5);
  VNStageIntLLRInputS4xD(38)(3) <= CNStageIntLLROutputS4xD(192)(0);
  VNStageIntLLRInputS4xD(75)(3) <= CNStageIntLLROutputS4xD(192)(1);
  VNStageIntLLRInputS4xD(143)(3) <= CNStageIntLLROutputS4xD(192)(2);
  VNStageIntLLRInputS4xD(249)(1) <= CNStageIntLLROutputS4xD(192)(3);
  VNStageIntLLRInputS4xD(289)(3) <= CNStageIntLLROutputS4xD(192)(4);
  VNStageIntLLRInputS4xD(352)(3) <= CNStageIntLLROutputS4xD(192)(5);
  VNStageIntLLRInputS4xD(37)(3) <= CNStageIntLLROutputS4xD(193)(0);
  VNStageIntLLRInputS4xD(78)(3) <= CNStageIntLLROutputS4xD(193)(1);
  VNStageIntLLRInputS4xD(184)(3) <= CNStageIntLLROutputS4xD(193)(2);
  VNStageIntLLRInputS4xD(224)(3) <= CNStageIntLLROutputS4xD(193)(3);
  VNStageIntLLRInputS4xD(287)(3) <= CNStageIntLLROutputS4xD(193)(4);
  VNStageIntLLRInputS4xD(377)(2) <= CNStageIntLLROutputS4xD(193)(5);
  VNStageIntLLRInputS4xD(35)(3) <= CNStageIntLLROutputS4xD(194)(0);
  VNStageIntLLRInputS4xD(94)(2) <= CNStageIntLLROutputS4xD(194)(1);
  VNStageIntLLRInputS4xD(157)(3) <= CNStageIntLLROutputS4xD(194)(2);
  VNStageIntLLRInputS4xD(247)(3) <= CNStageIntLLROutputS4xD(194)(3);
  VNStageIntLLRInputS4xD(257)(3) <= CNStageIntLLROutputS4xD(194)(4);
  VNStageIntLLRInputS4xD(365)(3) <= CNStageIntLLROutputS4xD(194)(5);
  VNStageIntLLRInputS4xD(34)(3) <= CNStageIntLLROutputS4xD(195)(0);
  VNStageIntLLRInputS4xD(92)(3) <= CNStageIntLLROutputS4xD(195)(1);
  VNStageIntLLRInputS4xD(182)(3) <= CNStageIntLLROutputS4xD(195)(2);
  VNStageIntLLRInputS4xD(255)(3) <= CNStageIntLLROutputS4xD(195)(3);
  VNStageIntLLRInputS4xD(300)(3) <= CNStageIntLLROutputS4xD(195)(4);
  VNStageIntLLRInputS4xD(359)(3) <= CNStageIntLLROutputS4xD(195)(5);
  VNStageIntLLRInputS4xD(33)(3) <= CNStageIntLLROutputS4xD(196)(0);
  VNStageIntLLRInputS4xD(117)(3) <= CNStageIntLLROutputS4xD(196)(1);
  VNStageIntLLRInputS4xD(190)(1) <= CNStageIntLLROutputS4xD(196)(2);
  VNStageIntLLRInputS4xD(235)(2) <= CNStageIntLLROutputS4xD(196)(3);
  VNStageIntLLRInputS4xD(294)(3) <= CNStageIntLLROutputS4xD(196)(4);
  VNStageIntLLRInputS4xD(320)(2) <= CNStageIntLLROutputS4xD(196)(5);
  VNStageIntLLRInputS4xD(31)(2) <= CNStageIntLLROutputS4xD(197)(0);
  VNStageIntLLRInputS4xD(105)(2) <= CNStageIntLLROutputS4xD(197)(1);
  VNStageIntLLRInputS4xD(164)(3) <= CNStageIntLLROutputS4xD(197)(2);
  VNStageIntLLRInputS4xD(192)(3) <= CNStageIntLLROutputS4xD(197)(3);
  VNStageIntLLRInputS4xD(293)(3) <= CNStageIntLLROutputS4xD(197)(4);
  VNStageIntLLRInputS4xD(363)(2) <= CNStageIntLLROutputS4xD(197)(5);
  VNStageIntLLRInputS4xD(30)(3) <= CNStageIntLLROutputS4xD(198)(0);
  VNStageIntLLRInputS4xD(99)(3) <= CNStageIntLLROutputS4xD(198)(1);
  VNStageIntLLRInputS4xD(128)(3) <= CNStageIntLLROutputS4xD(198)(2);
  VNStageIntLLRInputS4xD(228)(3) <= CNStageIntLLROutputS4xD(198)(3);
  VNStageIntLLRInputS4xD(298)(3) <= CNStageIntLLROutputS4xD(198)(4);
  VNStageIntLLRInputS4xD(382)(2) <= CNStageIntLLROutputS4xD(198)(5);
  VNStageIntLLRInputS4xD(28)(3) <= CNStageIntLLROutputS4xD(199)(0);
  VNStageIntLLRInputS4xD(98)(2) <= CNStageIntLLROutputS4xD(199)(1);
  VNStageIntLLRInputS4xD(168)(2) <= CNStageIntLLROutputS4xD(199)(2);
  VNStageIntLLRInputS4xD(252)(2) <= CNStageIntLLROutputS4xD(199)(3);
  VNStageIntLLRInputS4xD(308)(1) <= CNStageIntLLROutputS4xD(199)(4);
  VNStageIntLLRInputS4xD(347)(3) <= CNStageIntLLROutputS4xD(199)(5);
  VNStageIntLLRInputS4xD(27)(3) <= CNStageIntLLROutputS4xD(200)(0);
  VNStageIntLLRInputS4xD(103)(3) <= CNStageIntLLROutputS4xD(200)(1);
  VNStageIntLLRInputS4xD(187)(2) <= CNStageIntLLROutputS4xD(200)(2);
  VNStageIntLLRInputS4xD(243)(3) <= CNStageIntLLROutputS4xD(200)(3);
  VNStageIntLLRInputS4xD(282)(3) <= CNStageIntLLROutputS4xD(200)(4);
  VNStageIntLLRInputS4xD(348)(3) <= CNStageIntLLROutputS4xD(200)(5);
  VNStageIntLLRInputS4xD(26)(3) <= CNStageIntLLROutputS4xD(201)(0);
  VNStageIntLLRInputS4xD(122)(2) <= CNStageIntLLROutputS4xD(201)(1);
  VNStageIntLLRInputS4xD(178)(3) <= CNStageIntLLROutputS4xD(201)(2);
  VNStageIntLLRInputS4xD(217)(3) <= CNStageIntLLROutputS4xD(201)(3);
  VNStageIntLLRInputS4xD(283)(3) <= CNStageIntLLROutputS4xD(201)(4);
  VNStageIntLLRInputS4xD(372)(2) <= CNStageIntLLROutputS4xD(201)(5);
  VNStageIntLLRInputS4xD(25)(3) <= CNStageIntLLROutputS4xD(202)(0);
  VNStageIntLLRInputS4xD(113)(3) <= CNStageIntLLROutputS4xD(202)(1);
  VNStageIntLLRInputS4xD(152)(3) <= CNStageIntLLROutputS4xD(202)(2);
  VNStageIntLLRInputS4xD(218)(3) <= CNStageIntLLROutputS4xD(202)(3);
  VNStageIntLLRInputS4xD(307)(3) <= CNStageIntLLROutputS4xD(202)(4);
  VNStageIntLLRInputS4xD(330)(3) <= CNStageIntLLROutputS4xD(202)(5);
  VNStageIntLLRInputS4xD(24)(3) <= CNStageIntLLROutputS4xD(203)(0);
  VNStageIntLLRInputS4xD(87)(3) <= CNStageIntLLROutputS4xD(203)(1);
  VNStageIntLLRInputS4xD(153)(3) <= CNStageIntLLROutputS4xD(203)(2);
  VNStageIntLLRInputS4xD(242)(3) <= CNStageIntLLROutputS4xD(203)(3);
  VNStageIntLLRInputS4xD(265)(2) <= CNStageIntLLROutputS4xD(203)(4);
  VNStageIntLLRInputS4xD(326)(2) <= CNStageIntLLROutputS4xD(203)(5);
  VNStageIntLLRInputS4xD(23)(3) <= CNStageIntLLROutputS4xD(204)(0);
  VNStageIntLLRInputS4xD(88)(3) <= CNStageIntLLROutputS4xD(204)(1);
  VNStageIntLLRInputS4xD(177)(3) <= CNStageIntLLROutputS4xD(204)(2);
  VNStageIntLLRInputS4xD(200)(3) <= CNStageIntLLROutputS4xD(204)(3);
  VNStageIntLLRInputS4xD(261)(3) <= CNStageIntLLROutputS4xD(204)(4);
  VNStageIntLLRInputS4xD(341)(3) <= CNStageIntLLROutputS4xD(204)(5);
  VNStageIntLLRInputS4xD(22)(3) <= CNStageIntLLROutputS4xD(205)(0);
  VNStageIntLLRInputS4xD(112)(3) <= CNStageIntLLROutputS4xD(205)(1);
  VNStageIntLLRInputS4xD(135)(3) <= CNStageIntLLROutputS4xD(205)(2);
  VNStageIntLLRInputS4xD(196)(3) <= CNStageIntLLROutputS4xD(205)(3);
  VNStageIntLLRInputS4xD(276)(3) <= CNStageIntLLROutputS4xD(205)(4);
  VNStageIntLLRInputS4xD(367)(3) <= CNStageIntLLROutputS4xD(205)(5);
  VNStageIntLLRInputS4xD(21)(3) <= CNStageIntLLROutputS4xD(206)(0);
  VNStageIntLLRInputS4xD(70)(3) <= CNStageIntLLROutputS4xD(206)(1);
  VNStageIntLLRInputS4xD(131)(2) <= CNStageIntLLROutputS4xD(206)(2);
  VNStageIntLLRInputS4xD(211)(3) <= CNStageIntLLROutputS4xD(206)(3);
  VNStageIntLLRInputS4xD(302)(3) <= CNStageIntLLROutputS4xD(206)(4);
  VNStageIntLLRInputS4xD(343)(3) <= CNStageIntLLROutputS4xD(206)(5);
  VNStageIntLLRInputS4xD(18)(3) <= CNStageIntLLROutputS4xD(207)(0);
  VNStageIntLLRInputS4xD(107)(2) <= CNStageIntLLROutputS4xD(207)(1);
  VNStageIntLLRInputS4xD(148)(3) <= CNStageIntLLROutputS4xD(207)(2);
  VNStageIntLLRInputS4xD(245)(3) <= CNStageIntLLROutputS4xD(207)(3);
  VNStageIntLLRInputS4xD(263)(3) <= CNStageIntLLROutputS4xD(207)(4);
  VNStageIntLLRInputS4xD(361)(3) <= CNStageIntLLROutputS4xD(207)(5);
  VNStageIntLLRInputS4xD(17)(3) <= CNStageIntLLROutputS4xD(208)(0);
  VNStageIntLLRInputS4xD(83)(3) <= CNStageIntLLROutputS4xD(208)(1);
  VNStageIntLLRInputS4xD(180)(1) <= CNStageIntLLROutputS4xD(208)(2);
  VNStageIntLLRInputS4xD(198)(3) <= CNStageIntLLROutputS4xD(208)(3);
  VNStageIntLLRInputS4xD(296)(3) <= CNStageIntLLROutputS4xD(208)(4);
  VNStageIntLLRInputS4xD(370)(2) <= CNStageIntLLROutputS4xD(208)(5);
  VNStageIntLLRInputS4xD(16)(2) <= CNStageIntLLROutputS4xD(209)(0);
  VNStageIntLLRInputS4xD(115)(3) <= CNStageIntLLROutputS4xD(209)(1);
  VNStageIntLLRInputS4xD(133)(1) <= CNStageIntLLROutputS4xD(209)(2);
  VNStageIntLLRInputS4xD(231)(2) <= CNStageIntLLROutputS4xD(209)(3);
  VNStageIntLLRInputS4xD(305)(3) <= CNStageIntLLROutputS4xD(209)(4);
  VNStageIntLLRInputS4xD(383)(3) <= CNStageIntLLROutputS4xD(209)(5);
  VNStageIntLLRInputS4xD(15)(3) <= CNStageIntLLROutputS4xD(210)(0);
  VNStageIntLLRInputS4xD(68)(2) <= CNStageIntLLROutputS4xD(210)(1);
  VNStageIntLLRInputS4xD(166)(3) <= CNStageIntLLROutputS4xD(210)(2);
  VNStageIntLLRInputS4xD(240)(3) <= CNStageIntLLROutputS4xD(210)(3);
  VNStageIntLLRInputS4xD(318)(1) <= CNStageIntLLROutputS4xD(210)(4);
  VNStageIntLLRInputS4xD(362)(3) <= CNStageIntLLROutputS4xD(210)(5);
  VNStageIntLLRInputS4xD(14)(3) <= CNStageIntLLROutputS4xD(211)(0);
  VNStageIntLLRInputS4xD(101)(3) <= CNStageIntLLROutputS4xD(211)(1);
  VNStageIntLLRInputS4xD(175)(3) <= CNStageIntLLROutputS4xD(211)(2);
  VNStageIntLLRInputS4xD(253)(2) <= CNStageIntLLROutputS4xD(211)(3);
  VNStageIntLLRInputS4xD(297)(3) <= CNStageIntLLROutputS4xD(211)(4);
  VNStageIntLLRInputS4xD(327)(3) <= CNStageIntLLROutputS4xD(211)(5);
  VNStageIntLLRInputS4xD(13)(2) <= CNStageIntLLROutputS4xD(212)(0);
  VNStageIntLLRInputS4xD(110)(3) <= CNStageIntLLROutputS4xD(212)(1);
  VNStageIntLLRInputS4xD(188)(1) <= CNStageIntLLROutputS4xD(212)(2);
  VNStageIntLLRInputS4xD(232)(2) <= CNStageIntLLROutputS4xD(212)(3);
  VNStageIntLLRInputS4xD(262)(3) <= CNStageIntLLROutputS4xD(212)(4);
  VNStageIntLLRInputS4xD(329)(3) <= CNStageIntLLROutputS4xD(212)(5);
  VNStageIntLLRInputS4xD(12)(3) <= CNStageIntLLROutputS4xD(213)(0);
  VNStageIntLLRInputS4xD(123)(2) <= CNStageIntLLROutputS4xD(213)(1);
  VNStageIntLLRInputS4xD(167)(3) <= CNStageIntLLROutputS4xD(213)(2);
  VNStageIntLLRInputS4xD(197)(3) <= CNStageIntLLROutputS4xD(213)(3);
  VNStageIntLLRInputS4xD(264)(3) <= CNStageIntLLROutputS4xD(213)(4);
  VNStageIntLLRInputS4xD(374)(3) <= CNStageIntLLROutputS4xD(213)(5);
  VNStageIntLLRInputS4xD(11)(3) <= CNStageIntLLROutputS4xD(214)(0);
  VNStageIntLLRInputS4xD(102)(3) <= CNStageIntLLROutputS4xD(214)(1);
  VNStageIntLLRInputS4xD(132)(2) <= CNStageIntLLROutputS4xD(214)(2);
  VNStageIntLLRInputS4xD(199)(3) <= CNStageIntLLROutputS4xD(214)(3);
  VNStageIntLLRInputS4xD(309)(3) <= CNStageIntLLROutputS4xD(214)(4);
  VNStageIntLLRInputS4xD(381)(2) <= CNStageIntLLROutputS4xD(214)(5);
  VNStageIntLLRInputS4xD(9)(3) <= CNStageIntLLROutputS4xD(215)(0);
  VNStageIntLLRInputS4xD(69)(3) <= CNStageIntLLROutputS4xD(215)(1);
  VNStageIntLLRInputS4xD(179)(3) <= CNStageIntLLROutputS4xD(215)(2);
  VNStageIntLLRInputS4xD(251)(2) <= CNStageIntLLROutputS4xD(215)(3);
  VNStageIntLLRInputS4xD(280)(3) <= CNStageIntLLROutputS4xD(215)(4);
  VNStageIntLLRInputS4xD(333)(2) <= CNStageIntLLROutputS4xD(215)(5);
  VNStageIntLLRInputS4xD(8)(2) <= CNStageIntLLROutputS4xD(216)(0);
  VNStageIntLLRInputS4xD(114)(3) <= CNStageIntLLROutputS4xD(216)(1);
  VNStageIntLLRInputS4xD(186)(2) <= CNStageIntLLROutputS4xD(216)(2);
  VNStageIntLLRInputS4xD(215)(3) <= CNStageIntLLROutputS4xD(216)(3);
  VNStageIntLLRInputS4xD(268)(3) <= CNStageIntLLROutputS4xD(216)(4);
  VNStageIntLLRInputS4xD(339)(3) <= CNStageIntLLROutputS4xD(216)(5);
  VNStageIntLLRInputS4xD(7)(3) <= CNStageIntLLROutputS4xD(217)(0);
  VNStageIntLLRInputS4xD(121)(2) <= CNStageIntLLROutputS4xD(217)(1);
  VNStageIntLLRInputS4xD(150)(3) <= CNStageIntLLROutputS4xD(217)(2);
  VNStageIntLLRInputS4xD(203)(3) <= CNStageIntLLROutputS4xD(217)(3);
  VNStageIntLLRInputS4xD(274)(2) <= CNStageIntLLROutputS4xD(217)(4);
  VNStageIntLLRInputS4xD(334)(2) <= CNStageIntLLROutputS4xD(217)(5);
  VNStageIntLLRInputS4xD(6)(3) <= CNStageIntLLROutputS4xD(218)(0);
  VNStageIntLLRInputS4xD(85)(2) <= CNStageIntLLROutputS4xD(218)(1);
  VNStageIntLLRInputS4xD(138)(3) <= CNStageIntLLROutputS4xD(218)(2);
  VNStageIntLLRInputS4xD(209)(3) <= CNStageIntLLROutputS4xD(218)(3);
  VNStageIntLLRInputS4xD(269)(2) <= CNStageIntLLROutputS4xD(218)(4);
  VNStageIntLLRInputS4xD(344)(3) <= CNStageIntLLROutputS4xD(218)(5);
  VNStageIntLLRInputS4xD(5)(3) <= CNStageIntLLROutputS4xD(219)(0);
  VNStageIntLLRInputS4xD(73)(3) <= CNStageIntLLROutputS4xD(219)(1);
  VNStageIntLLRInputS4xD(144)(3) <= CNStageIntLLROutputS4xD(219)(2);
  VNStageIntLLRInputS4xD(204)(3) <= CNStageIntLLROutputS4xD(219)(3);
  VNStageIntLLRInputS4xD(279)(3) <= CNStageIntLLROutputS4xD(219)(4);
  VNStageIntLLRInputS4xD(366)(3) <= CNStageIntLLROutputS4xD(219)(5);
  VNStageIntLLRInputS4xD(4)(2) <= CNStageIntLLROutputS4xD(220)(0);
  VNStageIntLLRInputS4xD(79)(3) <= CNStageIntLLROutputS4xD(220)(1);
  VNStageIntLLRInputS4xD(139)(3) <= CNStageIntLLROutputS4xD(220)(2);
  VNStageIntLLRInputS4xD(214)(3) <= CNStageIntLLROutputS4xD(220)(3);
  VNStageIntLLRInputS4xD(301)(3) <= CNStageIntLLROutputS4xD(220)(4);
  VNStageIntLLRInputS4xD(321)(3) <= CNStageIntLLROutputS4xD(220)(5);
  VNStageIntLLRInputS4xD(3)(2) <= CNStageIntLLROutputS4xD(221)(0);
  VNStageIntLLRInputS4xD(74)(3) <= CNStageIntLLROutputS4xD(221)(1);
  VNStageIntLLRInputS4xD(149)(3) <= CNStageIntLLROutputS4xD(221)(2);
  VNStageIntLLRInputS4xD(236)(3) <= CNStageIntLLROutputS4xD(221)(3);
  VNStageIntLLRInputS4xD(319)(3) <= CNStageIntLLROutputS4xD(221)(4);
  VNStageIntLLRInputS4xD(369)(2) <= CNStageIntLLROutputS4xD(221)(5);
  VNStageIntLLRInputS4xD(2)(3) <= CNStageIntLLROutputS4xD(222)(0);
  VNStageIntLLRInputS4xD(84)(3) <= CNStageIntLLROutputS4xD(222)(1);
  VNStageIntLLRInputS4xD(171)(2) <= CNStageIntLLROutputS4xD(222)(2);
  VNStageIntLLRInputS4xD(254)(1) <= CNStageIntLLROutputS4xD(222)(3);
  VNStageIntLLRInputS4xD(304)(3) <= CNStageIntLLROutputS4xD(222)(4);
  VNStageIntLLRInputS4xD(356)(3) <= CNStageIntLLROutputS4xD(222)(5);
  VNStageIntLLRInputS4xD(1)(2) <= CNStageIntLLROutputS4xD(223)(0);
  VNStageIntLLRInputS4xD(106)(2) <= CNStageIntLLROutputS4xD(223)(1);
  VNStageIntLLRInputS4xD(189)(2) <= CNStageIntLLROutputS4xD(223)(2);
  VNStageIntLLRInputS4xD(239)(3) <= CNStageIntLLROutputS4xD(223)(3);
  VNStageIntLLRInputS4xD(291)(3) <= CNStageIntLLROutputS4xD(223)(4);
  VNStageIntLLRInputS4xD(324)(3) <= CNStageIntLLROutputS4xD(223)(5);
  VNStageIntLLRInputS4xD(0)(3) <= CNStageIntLLROutputS4xD(224)(0);
  VNStageIntLLRInputS4xD(93)(3) <= CNStageIntLLROutputS4xD(224)(1);
  VNStageIntLLRInputS4xD(158)(3) <= CNStageIntLLROutputS4xD(224)(2);
  VNStageIntLLRInputS4xD(223)(3) <= CNStageIntLLROutputS4xD(224)(3);
  VNStageIntLLRInputS4xD(288)(3) <= CNStageIntLLROutputS4xD(224)(4);
  VNStageIntLLRInputS4xD(353)(3) <= CNStageIntLLROutputS4xD(224)(5);
  VNStageIntLLRInputS4xD(18)(4) <= CNStageIntLLROutputS4xD(225)(0);
  VNStageIntLLRInputS4xD(110)(4) <= CNStageIntLLROutputS4xD(225)(1);
  VNStageIntLLRInputS4xD(167)(4) <= CNStageIntLLROutputS4xD(225)(2);
  VNStageIntLLRInputS4xD(249)(2) <= CNStageIntLLROutputS4xD(225)(3);
  VNStageIntLLRInputS4xD(311)(3) <= CNStageIntLLROutputS4xD(225)(4);
  VNStageIntLLRInputS4xD(347)(4) <= CNStageIntLLROutputS4xD(225)(5);
  VNStageIntLLRInputS4xD(17)(4) <= CNStageIntLLROutputS4xD(226)(0);
  VNStageIntLLRInputS4xD(102)(4) <= CNStageIntLLROutputS4xD(226)(1);
  VNStageIntLLRInputS4xD(184)(4) <= CNStageIntLLROutputS4xD(226)(2);
  VNStageIntLLRInputS4xD(246)(4) <= CNStageIntLLROutputS4xD(226)(3);
  VNStageIntLLRInputS4xD(282)(4) <= CNStageIntLLROutputS4xD(226)(4);
  VNStageIntLLRInputS4xD(367)(4) <= CNStageIntLLROutputS4xD(226)(5);
  VNStageIntLLRInputS4xD(16)(3) <= CNStageIntLLROutputS4xD(227)(0);
  VNStageIntLLRInputS4xD(119)(3) <= CNStageIntLLROutputS4xD(227)(1);
  VNStageIntLLRInputS4xD(181)(4) <= CNStageIntLLROutputS4xD(227)(2);
  VNStageIntLLRInputS4xD(217)(4) <= CNStageIntLLROutputS4xD(227)(3);
  VNStageIntLLRInputS4xD(302)(4) <= CNStageIntLLROutputS4xD(227)(4);
  VNStageIntLLRInputS4xD(353)(4) <= CNStageIntLLROutputS4xD(227)(5);
  VNStageIntLLRInputS4xD(15)(4) <= CNStageIntLLROutputS4xD(228)(0);
  VNStageIntLLRInputS4xD(116)(3) <= CNStageIntLLROutputS4xD(228)(1);
  VNStageIntLLRInputS4xD(152)(4) <= CNStageIntLLROutputS4xD(228)(2);
  VNStageIntLLRInputS4xD(237)(3) <= CNStageIntLLROutputS4xD(228)(3);
  VNStageIntLLRInputS4xD(288)(4) <= CNStageIntLLROutputS4xD(228)(4);
  VNStageIntLLRInputS4xD(343)(4) <= CNStageIntLLROutputS4xD(228)(5);
  VNStageIntLLRInputS4xD(14)(4) <= CNStageIntLLROutputS4xD(229)(0);
  VNStageIntLLRInputS4xD(87)(4) <= CNStageIntLLROutputS4xD(229)(1);
  VNStageIntLLRInputS4xD(172)(3) <= CNStageIntLLROutputS4xD(229)(2);
  VNStageIntLLRInputS4xD(223)(4) <= CNStageIntLLROutputS4xD(229)(3);
  VNStageIntLLRInputS4xD(278)(3) <= CNStageIntLLROutputS4xD(229)(4);
  VNStageIntLLRInputS4xD(372)(3) <= CNStageIntLLROutputS4xD(229)(5);
  VNStageIntLLRInputS4xD(13)(3) <= CNStageIntLLROutputS4xD(230)(0);
  VNStageIntLLRInputS4xD(107)(3) <= CNStageIntLLROutputS4xD(230)(1);
  VNStageIntLLRInputS4xD(158)(4) <= CNStageIntLLROutputS4xD(230)(2);
  VNStageIntLLRInputS4xD(213)(3) <= CNStageIntLLROutputS4xD(230)(3);
  VNStageIntLLRInputS4xD(307)(4) <= CNStageIntLLROutputS4xD(230)(4);
  VNStageIntLLRInputS4xD(355)(4) <= CNStageIntLLROutputS4xD(230)(5);
  VNStageIntLLRInputS4xD(12)(4) <= CNStageIntLLROutputS4xD(231)(0);
  VNStageIntLLRInputS4xD(93)(4) <= CNStageIntLLROutputS4xD(231)(1);
  VNStageIntLLRInputS4xD(148)(4) <= CNStageIntLLROutputS4xD(231)(2);
  VNStageIntLLRInputS4xD(242)(4) <= CNStageIntLLROutputS4xD(231)(3);
  VNStageIntLLRInputS4xD(290)(4) <= CNStageIntLLROutputS4xD(231)(4);
  VNStageIntLLRInputS4xD(322)(3) <= CNStageIntLLROutputS4xD(231)(5);
  VNStageIntLLRInputS4xD(11)(4) <= CNStageIntLLROutputS4xD(232)(0);
  VNStageIntLLRInputS4xD(83)(4) <= CNStageIntLLROutputS4xD(232)(1);
  VNStageIntLLRInputS4xD(177)(4) <= CNStageIntLLROutputS4xD(232)(2);
  VNStageIntLLRInputS4xD(225)(4) <= CNStageIntLLROutputS4xD(232)(3);
  VNStageIntLLRInputS4xD(257)(4) <= CNStageIntLLROutputS4xD(232)(4);
  VNStageIntLLRInputS4xD(345)(3) <= CNStageIntLLROutputS4xD(232)(5);
  VNStageIntLLRInputS4xD(10)(3) <= CNStageIntLLROutputS4xD(233)(0);
  VNStageIntLLRInputS4xD(112)(4) <= CNStageIntLLROutputS4xD(233)(1);
  VNStageIntLLRInputS4xD(160)(4) <= CNStageIntLLROutputS4xD(233)(2);
  VNStageIntLLRInputS4xD(255)(4) <= CNStageIntLLROutputS4xD(233)(3);
  VNStageIntLLRInputS4xD(280)(4) <= CNStageIntLLROutputS4xD(233)(4);
  VNStageIntLLRInputS4xD(381)(3) <= CNStageIntLLROutputS4xD(233)(5);
  VNStageIntLLRInputS4xD(9)(4) <= CNStageIntLLROutputS4xD(234)(0);
  VNStageIntLLRInputS4xD(95)(4) <= CNStageIntLLROutputS4xD(234)(1);
  VNStageIntLLRInputS4xD(190)(2) <= CNStageIntLLROutputS4xD(234)(2);
  VNStageIntLLRInputS4xD(215)(4) <= CNStageIntLLROutputS4xD(234)(3);
  VNStageIntLLRInputS4xD(316)(2) <= CNStageIntLLROutputS4xD(234)(4);
  VNStageIntLLRInputS4xD(365)(4) <= CNStageIntLLROutputS4xD(234)(5);
  VNStageIntLLRInputS4xD(7)(4) <= CNStageIntLLROutputS4xD(235)(0);
  VNStageIntLLRInputS4xD(85)(3) <= CNStageIntLLROutputS4xD(235)(1);
  VNStageIntLLRInputS4xD(186)(3) <= CNStageIntLLROutputS4xD(235)(2);
  VNStageIntLLRInputS4xD(235)(3) <= CNStageIntLLROutputS4xD(235)(3);
  VNStageIntLLRInputS4xD(303)(4) <= CNStageIntLLROutputS4xD(235)(4);
  VNStageIntLLRInputS4xD(346)(4) <= CNStageIntLLROutputS4xD(235)(5);
  VNStageIntLLRInputS4xD(6)(4) <= CNStageIntLLROutputS4xD(236)(0);
  VNStageIntLLRInputS4xD(121)(3) <= CNStageIntLLROutputS4xD(236)(1);
  VNStageIntLLRInputS4xD(170)(3) <= CNStageIntLLROutputS4xD(236)(2);
  VNStageIntLLRInputS4xD(238)(4) <= CNStageIntLLROutputS4xD(236)(3);
  VNStageIntLLRInputS4xD(281)(4) <= CNStageIntLLROutputS4xD(236)(4);
  VNStageIntLLRInputS4xD(321)(4) <= CNStageIntLLROutputS4xD(236)(5);
  VNStageIntLLRInputS4xD(5)(4) <= CNStageIntLLROutputS4xD(237)(0);
  VNStageIntLLRInputS4xD(105)(3) <= CNStageIntLLROutputS4xD(237)(1);
  VNStageIntLLRInputS4xD(173)(4) <= CNStageIntLLROutputS4xD(237)(2);
  VNStageIntLLRInputS4xD(216)(4) <= CNStageIntLLROutputS4xD(237)(3);
  VNStageIntLLRInputS4xD(319)(4) <= CNStageIntLLROutputS4xD(237)(4);
  VNStageIntLLRInputS4xD(382)(3) <= CNStageIntLLROutputS4xD(237)(5);
  VNStageIntLLRInputS4xD(4)(3) <= CNStageIntLLROutputS4xD(238)(0);
  VNStageIntLLRInputS4xD(108)(4) <= CNStageIntLLROutputS4xD(238)(1);
  VNStageIntLLRInputS4xD(151)(4) <= CNStageIntLLROutputS4xD(238)(2);
  VNStageIntLLRInputS4xD(254)(2) <= CNStageIntLLROutputS4xD(238)(3);
  VNStageIntLLRInputS4xD(317)(1) <= CNStageIntLLROutputS4xD(238)(4);
  VNStageIntLLRInputS4xD(344)(4) <= CNStageIntLLROutputS4xD(238)(5);
  VNStageIntLLRInputS4xD(3)(3) <= CNStageIntLLROutputS4xD(239)(0);
  VNStageIntLLRInputS4xD(86)(2) <= CNStageIntLLROutputS4xD(239)(1);
  VNStageIntLLRInputS4xD(189)(3) <= CNStageIntLLROutputS4xD(239)(2);
  VNStageIntLLRInputS4xD(252)(3) <= CNStageIntLLROutputS4xD(239)(3);
  VNStageIntLLRInputS4xD(279)(4) <= CNStageIntLLROutputS4xD(239)(4);
  VNStageIntLLRInputS4xD(352)(4) <= CNStageIntLLROutputS4xD(239)(5);
  VNStageIntLLRInputS4xD(2)(4) <= CNStageIntLLROutputS4xD(240)(0);
  VNStageIntLLRInputS4xD(124)(2) <= CNStageIntLLROutputS4xD(240)(1);
  VNStageIntLLRInputS4xD(187)(3) <= CNStageIntLLROutputS4xD(240)(2);
  VNStageIntLLRInputS4xD(214)(4) <= CNStageIntLLROutputS4xD(240)(3);
  VNStageIntLLRInputS4xD(287)(4) <= CNStageIntLLROutputS4xD(240)(4);
  VNStageIntLLRInputS4xD(332)(4) <= CNStageIntLLROutputS4xD(240)(5);
  VNStageIntLLRInputS4xD(1)(3) <= CNStageIntLLROutputS4xD(241)(0);
  VNStageIntLLRInputS4xD(122)(3) <= CNStageIntLLROutputS4xD(241)(1);
  VNStageIntLLRInputS4xD(149)(4) <= CNStageIntLLROutputS4xD(241)(2);
  VNStageIntLLRInputS4xD(222)(2) <= CNStageIntLLROutputS4xD(241)(3);
  VNStageIntLLRInputS4xD(267)(4) <= CNStageIntLLROutputS4xD(241)(4);
  VNStageIntLLRInputS4xD(326)(3) <= CNStageIntLLROutputS4xD(241)(5);
  VNStageIntLLRInputS4xD(62)(3) <= CNStageIntLLROutputS4xD(242)(0);
  VNStageIntLLRInputS4xD(92)(4) <= CNStageIntLLROutputS4xD(242)(1);
  VNStageIntLLRInputS4xD(137)(4) <= CNStageIntLLROutputS4xD(242)(2);
  VNStageIntLLRInputS4xD(196)(4) <= CNStageIntLLROutputS4xD(242)(3);
  VNStageIntLLRInputS4xD(256)(3) <= CNStageIntLLROutputS4xD(242)(4);
  VNStageIntLLRInputS4xD(325)(4) <= CNStageIntLLROutputS4xD(242)(5);
  VNStageIntLLRInputS4xD(61)(3) <= CNStageIntLLROutputS4xD(243)(0);
  VNStageIntLLRInputS4xD(72)(4) <= CNStageIntLLROutputS4xD(243)(1);
  VNStageIntLLRInputS4xD(131)(3) <= CNStageIntLLROutputS4xD(243)(2);
  VNStageIntLLRInputS4xD(192)(4) <= CNStageIntLLROutputS4xD(243)(3);
  VNStageIntLLRInputS4xD(260)(4) <= CNStageIntLLROutputS4xD(243)(4);
  VNStageIntLLRInputS4xD(330)(4) <= CNStageIntLLROutputS4xD(243)(5);
  VNStageIntLLRInputS4xD(60)(3) <= CNStageIntLLROutputS4xD(244)(0);
  VNStageIntLLRInputS4xD(66)(3) <= CNStageIntLLROutputS4xD(244)(1);
  VNStageIntLLRInputS4xD(128)(4) <= CNStageIntLLROutputS4xD(244)(2);
  VNStageIntLLRInputS4xD(195)(3) <= CNStageIntLLROutputS4xD(244)(3);
  VNStageIntLLRInputS4xD(265)(3) <= CNStageIntLLROutputS4xD(244)(4);
  VNStageIntLLRInputS4xD(349)(3) <= CNStageIntLLROutputS4xD(244)(5);
  VNStageIntLLRInputS4xD(59)(2) <= CNStageIntLLROutputS4xD(245)(0);
  VNStageIntLLRInputS4xD(64)(3) <= CNStageIntLLROutputS4xD(245)(1);
  VNStageIntLLRInputS4xD(130)(4) <= CNStageIntLLROutputS4xD(245)(2);
  VNStageIntLLRInputS4xD(200)(4) <= CNStageIntLLROutputS4xD(245)(3);
  VNStageIntLLRInputS4xD(284)(4) <= CNStageIntLLROutputS4xD(245)(4);
  VNStageIntLLRInputS4xD(340)(4) <= CNStageIntLLROutputS4xD(245)(5);
  VNStageIntLLRInputS4xD(57)(3) <= CNStageIntLLROutputS4xD(246)(0);
  VNStageIntLLRInputS4xD(70)(4) <= CNStageIntLLROutputS4xD(246)(1);
  VNStageIntLLRInputS4xD(154)(3) <= CNStageIntLLROutputS4xD(246)(2);
  VNStageIntLLRInputS4xD(210)(4) <= CNStageIntLLROutputS4xD(246)(3);
  VNStageIntLLRInputS4xD(312)(3) <= CNStageIntLLROutputS4xD(246)(4);
  VNStageIntLLRInputS4xD(378)(3) <= CNStageIntLLROutputS4xD(246)(5);
  VNStageIntLLRInputS4xD(56)(4) <= CNStageIntLLROutputS4xD(247)(0);
  VNStageIntLLRInputS4xD(89)(4) <= CNStageIntLLROutputS4xD(247)(1);
  VNStageIntLLRInputS4xD(145)(4) <= CNStageIntLLROutputS4xD(247)(2);
  VNStageIntLLRInputS4xD(247)(4) <= CNStageIntLLROutputS4xD(247)(3);
  VNStageIntLLRInputS4xD(313)(2) <= CNStageIntLLROutputS4xD(247)(4);
  VNStageIntLLRInputS4xD(339)(4) <= CNStageIntLLROutputS4xD(247)(5);
  VNStageIntLLRInputS4xD(55)(4) <= CNStageIntLLROutputS4xD(248)(0);
  VNStageIntLLRInputS4xD(80)(4) <= CNStageIntLLROutputS4xD(248)(1);
  VNStageIntLLRInputS4xD(182)(4) <= CNStageIntLLROutputS4xD(248)(2);
  VNStageIntLLRInputS4xD(248)(4) <= CNStageIntLLROutputS4xD(248)(3);
  VNStageIntLLRInputS4xD(274)(3) <= CNStageIntLLROutputS4xD(248)(4);
  VNStageIntLLRInputS4xD(360)(4) <= CNStageIntLLROutputS4xD(248)(5);
  VNStageIntLLRInputS4xD(53)(3) <= CNStageIntLLROutputS4xD(249)(0);
  VNStageIntLLRInputS4xD(118)(3) <= CNStageIntLLROutputS4xD(249)(1);
  VNStageIntLLRInputS4xD(144)(4) <= CNStageIntLLROutputS4xD(249)(2);
  VNStageIntLLRInputS4xD(230)(3) <= CNStageIntLLROutputS4xD(249)(3);
  VNStageIntLLRInputS4xD(291)(4) <= CNStageIntLLROutputS4xD(249)(4);
  VNStageIntLLRInputS4xD(371)(3) <= CNStageIntLLROutputS4xD(249)(5);
  VNStageIntLLRInputS4xD(51)(3) <= CNStageIntLLROutputS4xD(250)(0);
  VNStageIntLLRInputS4xD(100)(4) <= CNStageIntLLROutputS4xD(250)(1);
  VNStageIntLLRInputS4xD(161)(4) <= CNStageIntLLROutputS4xD(250)(2);
  VNStageIntLLRInputS4xD(241)(3) <= CNStageIntLLROutputS4xD(250)(3);
  VNStageIntLLRInputS4xD(269)(3) <= CNStageIntLLROutputS4xD(250)(4);
  VNStageIntLLRInputS4xD(373)(2) <= CNStageIntLLROutputS4xD(250)(5);
  VNStageIntLLRInputS4xD(50)(4) <= CNStageIntLLROutputS4xD(251)(0);
  VNStageIntLLRInputS4xD(96)(4) <= CNStageIntLLROutputS4xD(251)(1);
  VNStageIntLLRInputS4xD(176)(4) <= CNStageIntLLROutputS4xD(251)(2);
  VNStageIntLLRInputS4xD(204)(4) <= CNStageIntLLROutputS4xD(251)(3);
  VNStageIntLLRInputS4xD(308)(2) <= CNStageIntLLROutputS4xD(251)(4);
  VNStageIntLLRInputS4xD(342)(3) <= CNStageIntLLROutputS4xD(251)(5);
  VNStageIntLLRInputS4xD(49)(4) <= CNStageIntLLROutputS4xD(252)(0);
  VNStageIntLLRInputS4xD(111)(4) <= CNStageIntLLROutputS4xD(252)(1);
  VNStageIntLLRInputS4xD(139)(4) <= CNStageIntLLROutputS4xD(252)(2);
  VNStageIntLLRInputS4xD(243)(4) <= CNStageIntLLROutputS4xD(252)(3);
  VNStageIntLLRInputS4xD(277)(4) <= CNStageIntLLROutputS4xD(252)(4);
  VNStageIntLLRInputS4xD(358)(3) <= CNStageIntLLROutputS4xD(252)(5);
  VNStageIntLLRInputS4xD(47)(2) <= CNStageIntLLROutputS4xD(253)(0);
  VNStageIntLLRInputS4xD(113)(4) <= CNStageIntLLROutputS4xD(253)(1);
  VNStageIntLLRInputS4xD(147)(4) <= CNStageIntLLROutputS4xD(253)(2);
  VNStageIntLLRInputS4xD(228)(4) <= CNStageIntLLROutputS4xD(253)(3);
  VNStageIntLLRInputS4xD(263)(4) <= CNStageIntLLROutputS4xD(253)(4);
  VNStageIntLLRInputS4xD(337)(4) <= CNStageIntLLROutputS4xD(253)(5);
  VNStageIntLLRInputS4xD(46)(4) <= CNStageIntLLROutputS4xD(254)(0);
  VNStageIntLLRInputS4xD(82)(4) <= CNStageIntLLROutputS4xD(254)(1);
  VNStageIntLLRInputS4xD(163)(3) <= CNStageIntLLROutputS4xD(254)(2);
  VNStageIntLLRInputS4xD(198)(4) <= CNStageIntLLROutputS4xD(254)(3);
  VNStageIntLLRInputS4xD(272)(4) <= CNStageIntLLROutputS4xD(254)(4);
  VNStageIntLLRInputS4xD(350)(4) <= CNStageIntLLROutputS4xD(254)(5);
  VNStageIntLLRInputS4xD(45)(4) <= CNStageIntLLROutputS4xD(255)(0);
  VNStageIntLLRInputS4xD(98)(3) <= CNStageIntLLROutputS4xD(255)(1);
  VNStageIntLLRInputS4xD(133)(2) <= CNStageIntLLROutputS4xD(255)(2);
  VNStageIntLLRInputS4xD(207)(3) <= CNStageIntLLROutputS4xD(255)(3);
  VNStageIntLLRInputS4xD(285)(4) <= CNStageIntLLROutputS4xD(255)(4);
  VNStageIntLLRInputS4xD(329)(4) <= CNStageIntLLROutputS4xD(255)(5);
  VNStageIntLLRInputS4xD(44)(4) <= CNStageIntLLROutputS4xD(256)(0);
  VNStageIntLLRInputS4xD(68)(3) <= CNStageIntLLROutputS4xD(256)(1);
  VNStageIntLLRInputS4xD(142)(3) <= CNStageIntLLROutputS4xD(256)(2);
  VNStageIntLLRInputS4xD(220)(4) <= CNStageIntLLROutputS4xD(256)(3);
  VNStageIntLLRInputS4xD(264)(4) <= CNStageIntLLROutputS4xD(256)(4);
  VNStageIntLLRInputS4xD(357)(4) <= CNStageIntLLROutputS4xD(256)(5);
  VNStageIntLLRInputS4xD(43)(3) <= CNStageIntLLROutputS4xD(257)(0);
  VNStageIntLLRInputS4xD(77)(2) <= CNStageIntLLROutputS4xD(257)(1);
  VNStageIntLLRInputS4xD(155)(4) <= CNStageIntLLROutputS4xD(257)(2);
  VNStageIntLLRInputS4xD(199)(4) <= CNStageIntLLROutputS4xD(257)(3);
  VNStageIntLLRInputS4xD(292)(4) <= CNStageIntLLROutputS4xD(257)(4);
  VNStageIntLLRInputS4xD(359)(4) <= CNStageIntLLROutputS4xD(257)(5);
  VNStageIntLLRInputS4xD(42)(4) <= CNStageIntLLROutputS4xD(258)(0);
  VNStageIntLLRInputS4xD(90)(4) <= CNStageIntLLROutputS4xD(258)(1);
  VNStageIntLLRInputS4xD(134)(3) <= CNStageIntLLROutputS4xD(258)(2);
  VNStageIntLLRInputS4xD(227)(4) <= CNStageIntLLROutputS4xD(258)(3);
  VNStageIntLLRInputS4xD(294)(4) <= CNStageIntLLROutputS4xD(258)(4);
  VNStageIntLLRInputS4xD(341)(4) <= CNStageIntLLROutputS4xD(258)(5);
  VNStageIntLLRInputS4xD(41)(4) <= CNStageIntLLROutputS4xD(259)(0);
  VNStageIntLLRInputS4xD(69)(4) <= CNStageIntLLROutputS4xD(259)(1);
  VNStageIntLLRInputS4xD(162)(4) <= CNStageIntLLROutputS4xD(259)(2);
  VNStageIntLLRInputS4xD(229)(3) <= CNStageIntLLROutputS4xD(259)(3);
  VNStageIntLLRInputS4xD(276)(4) <= CNStageIntLLROutputS4xD(259)(4);
  VNStageIntLLRInputS4xD(348)(4) <= CNStageIntLLROutputS4xD(259)(5);
  VNStageIntLLRInputS4xD(40)(3) <= CNStageIntLLROutputS4xD(260)(0);
  VNStageIntLLRInputS4xD(97)(4) <= CNStageIntLLROutputS4xD(260)(1);
  VNStageIntLLRInputS4xD(164)(4) <= CNStageIntLLROutputS4xD(260)(2);
  VNStageIntLLRInputS4xD(211)(4) <= CNStageIntLLROutputS4xD(260)(3);
  VNStageIntLLRInputS4xD(283)(4) <= CNStageIntLLROutputS4xD(260)(4);
  VNStageIntLLRInputS4xD(375)(3) <= CNStageIntLLROutputS4xD(260)(5);
  VNStageIntLLRInputS4xD(39)(4) <= CNStageIntLLROutputS4xD(261)(0);
  VNStageIntLLRInputS4xD(99)(4) <= CNStageIntLLROutputS4xD(261)(1);
  VNStageIntLLRInputS4xD(146)(3) <= CNStageIntLLROutputS4xD(261)(2);
  VNStageIntLLRInputS4xD(218)(4) <= CNStageIntLLROutputS4xD(261)(3);
  VNStageIntLLRInputS4xD(310)(3) <= CNStageIntLLROutputS4xD(261)(4);
  VNStageIntLLRInputS4xD(363)(3) <= CNStageIntLLROutputS4xD(261)(5);
  VNStageIntLLRInputS4xD(38)(4) <= CNStageIntLLROutputS4xD(262)(0);
  VNStageIntLLRInputS4xD(81)(3) <= CNStageIntLLROutputS4xD(262)(1);
  VNStageIntLLRInputS4xD(153)(4) <= CNStageIntLLROutputS4xD(262)(2);
  VNStageIntLLRInputS4xD(245)(4) <= CNStageIntLLROutputS4xD(262)(3);
  VNStageIntLLRInputS4xD(298)(4) <= CNStageIntLLROutputS4xD(262)(4);
  VNStageIntLLRInputS4xD(369)(3) <= CNStageIntLLROutputS4xD(262)(5);
  VNStageIntLLRInputS4xD(37)(4) <= CNStageIntLLROutputS4xD(263)(0);
  VNStageIntLLRInputS4xD(88)(4) <= CNStageIntLLROutputS4xD(263)(1);
  VNStageIntLLRInputS4xD(180)(2) <= CNStageIntLLROutputS4xD(263)(2);
  VNStageIntLLRInputS4xD(233)(3) <= CNStageIntLLROutputS4xD(263)(3);
  VNStageIntLLRInputS4xD(304)(4) <= CNStageIntLLROutputS4xD(263)(4);
  VNStageIntLLRInputS4xD(364)(4) <= CNStageIntLLROutputS4xD(263)(5);
  VNStageIntLLRInputS4xD(36)(3) <= CNStageIntLLROutputS4xD(264)(0);
  VNStageIntLLRInputS4xD(115)(4) <= CNStageIntLLROutputS4xD(264)(1);
  VNStageIntLLRInputS4xD(168)(3) <= CNStageIntLLROutputS4xD(264)(2);
  VNStageIntLLRInputS4xD(239)(4) <= CNStageIntLLROutputS4xD(264)(3);
  VNStageIntLLRInputS4xD(299)(3) <= CNStageIntLLROutputS4xD(264)(4);
  VNStageIntLLRInputS4xD(374)(4) <= CNStageIntLLROutputS4xD(264)(5);
  VNStageIntLLRInputS4xD(35)(4) <= CNStageIntLLROutputS4xD(265)(0);
  VNStageIntLLRInputS4xD(103)(4) <= CNStageIntLLROutputS4xD(265)(1);
  VNStageIntLLRInputS4xD(174)(3) <= CNStageIntLLROutputS4xD(265)(2);
  VNStageIntLLRInputS4xD(234)(4) <= CNStageIntLLROutputS4xD(265)(3);
  VNStageIntLLRInputS4xD(309)(4) <= CNStageIntLLROutputS4xD(265)(4);
  VNStageIntLLRInputS4xD(333)(3) <= CNStageIntLLROutputS4xD(265)(5);
  VNStageIntLLRInputS4xD(34)(4) <= CNStageIntLLROutputS4xD(266)(0);
  VNStageIntLLRInputS4xD(109)(4) <= CNStageIntLLROutputS4xD(266)(1);
  VNStageIntLLRInputS4xD(169)(4) <= CNStageIntLLROutputS4xD(266)(2);
  VNStageIntLLRInputS4xD(244)(1) <= CNStageIntLLROutputS4xD(266)(3);
  VNStageIntLLRInputS4xD(268)(4) <= CNStageIntLLROutputS4xD(266)(4);
  VNStageIntLLRInputS4xD(351)(3) <= CNStageIntLLROutputS4xD(266)(5);
  VNStageIntLLRInputS4xD(33)(4) <= CNStageIntLLROutputS4xD(267)(0);
  VNStageIntLLRInputS4xD(104)(4) <= CNStageIntLLROutputS4xD(267)(1);
  VNStageIntLLRInputS4xD(179)(4) <= CNStageIntLLROutputS4xD(267)(2);
  VNStageIntLLRInputS4xD(203)(4) <= CNStageIntLLROutputS4xD(267)(3);
  VNStageIntLLRInputS4xD(286)(4) <= CNStageIntLLROutputS4xD(267)(4);
  VNStageIntLLRInputS4xD(336)(3) <= CNStageIntLLROutputS4xD(267)(5);
  VNStageIntLLRInputS4xD(32)(3) <= CNStageIntLLROutputS4xD(268)(0);
  VNStageIntLLRInputS4xD(114)(4) <= CNStageIntLLROutputS4xD(268)(1);
  VNStageIntLLRInputS4xD(138)(4) <= CNStageIntLLROutputS4xD(268)(2);
  VNStageIntLLRInputS4xD(221)(4) <= CNStageIntLLROutputS4xD(268)(3);
  VNStageIntLLRInputS4xD(271)(3) <= CNStageIntLLROutputS4xD(268)(4);
  VNStageIntLLRInputS4xD(323)(3) <= CNStageIntLLROutputS4xD(268)(5);
  VNStageIntLLRInputS4xD(30)(4) <= CNStageIntLLROutputS4xD(269)(0);
  VNStageIntLLRInputS4xD(91)(4) <= CNStageIntLLROutputS4xD(269)(1);
  VNStageIntLLRInputS4xD(141)(2) <= CNStageIntLLROutputS4xD(269)(2);
  VNStageIntLLRInputS4xD(193)(3) <= CNStageIntLLROutputS4xD(269)(3);
  VNStageIntLLRInputS4xD(289)(4) <= CNStageIntLLROutputS4xD(269)(4);
  VNStageIntLLRInputS4xD(366)(4) <= CNStageIntLLROutputS4xD(269)(5);
  VNStageIntLLRInputS4xD(29)(3) <= CNStageIntLLROutputS4xD(270)(0);
  VNStageIntLLRInputS4xD(76)(4) <= CNStageIntLLROutputS4xD(270)(1);
  VNStageIntLLRInputS4xD(191)(4) <= CNStageIntLLROutputS4xD(270)(2);
  VNStageIntLLRInputS4xD(224)(4) <= CNStageIntLLROutputS4xD(270)(3);
  VNStageIntLLRInputS4xD(301)(4) <= CNStageIntLLROutputS4xD(270)(4);
  VNStageIntLLRInputS4xD(380)(3) <= CNStageIntLLROutputS4xD(270)(5);
  VNStageIntLLRInputS4xD(28)(4) <= CNStageIntLLROutputS4xD(271)(0);
  VNStageIntLLRInputS4xD(126)(3) <= CNStageIntLLROutputS4xD(271)(1);
  VNStageIntLLRInputS4xD(159)(3) <= CNStageIntLLROutputS4xD(271)(2);
  VNStageIntLLRInputS4xD(236)(4) <= CNStageIntLLROutputS4xD(271)(3);
  VNStageIntLLRInputS4xD(315)(3) <= CNStageIntLLROutputS4xD(271)(4);
  VNStageIntLLRInputS4xD(361)(4) <= CNStageIntLLROutputS4xD(271)(5);
  VNStageIntLLRInputS4xD(26)(4) <= CNStageIntLLROutputS4xD(272)(0);
  VNStageIntLLRInputS4xD(106)(3) <= CNStageIntLLROutputS4xD(272)(1);
  VNStageIntLLRInputS4xD(185)(1) <= CNStageIntLLROutputS4xD(272)(2);
  VNStageIntLLRInputS4xD(231)(3) <= CNStageIntLLROutputS4xD(272)(3);
  VNStageIntLLRInputS4xD(273)(3) <= CNStageIntLLROutputS4xD(272)(4);
  VNStageIntLLRInputS4xD(327)(4) <= CNStageIntLLROutputS4xD(272)(5);
  VNStageIntLLRInputS4xD(24)(4) <= CNStageIntLLROutputS4xD(273)(0);
  VNStageIntLLRInputS4xD(101)(4) <= CNStageIntLLROutputS4xD(273)(1);
  VNStageIntLLRInputS4xD(143)(4) <= CNStageIntLLROutputS4xD(273)(2);
  VNStageIntLLRInputS4xD(197)(4) <= CNStageIntLLROutputS4xD(273)(3);
  VNStageIntLLRInputS4xD(266)(3) <= CNStageIntLLROutputS4xD(273)(4);
  VNStageIntLLRInputS4xD(324)(4) <= CNStageIntLLROutputS4xD(273)(5);
  VNStageIntLLRInputS4xD(23)(4) <= CNStageIntLLROutputS4xD(274)(0);
  VNStageIntLLRInputS4xD(78)(4) <= CNStageIntLLROutputS4xD(274)(1);
  VNStageIntLLRInputS4xD(132)(3) <= CNStageIntLLROutputS4xD(274)(2);
  VNStageIntLLRInputS4xD(201)(4) <= CNStageIntLLROutputS4xD(274)(3);
  VNStageIntLLRInputS4xD(259)(2) <= CNStageIntLLROutputS4xD(274)(4);
  VNStageIntLLRInputS4xD(335)(4) <= CNStageIntLLROutputS4xD(274)(5);
  VNStageIntLLRInputS4xD(22)(4) <= CNStageIntLLROutputS4xD(275)(0);
  VNStageIntLLRInputS4xD(67)(1) <= CNStageIntLLROutputS4xD(275)(1);
  VNStageIntLLRInputS4xD(136)(4) <= CNStageIntLLROutputS4xD(275)(2);
  VNStageIntLLRInputS4xD(194)(4) <= CNStageIntLLROutputS4xD(275)(3);
  VNStageIntLLRInputS4xD(270)(4) <= CNStageIntLLROutputS4xD(275)(4);
  VNStageIntLLRInputS4xD(370)(3) <= CNStageIntLLROutputS4xD(275)(5);
  VNStageIntLLRInputS4xD(21)(4) <= CNStageIntLLROutputS4xD(276)(0);
  VNStageIntLLRInputS4xD(71)(3) <= CNStageIntLLROutputS4xD(276)(1);
  VNStageIntLLRInputS4xD(129)(4) <= CNStageIntLLROutputS4xD(276)(2);
  VNStageIntLLRInputS4xD(205)(1) <= CNStageIntLLROutputS4xD(276)(3);
  VNStageIntLLRInputS4xD(305)(4) <= CNStageIntLLROutputS4xD(276)(4);
  VNStageIntLLRInputS4xD(362)(4) <= CNStageIntLLROutputS4xD(276)(5);
  VNStageIntLLRInputS4xD(20)(2) <= CNStageIntLLROutputS4xD(277)(0);
  VNStageIntLLRInputS4xD(127)(4) <= CNStageIntLLROutputS4xD(277)(1);
  VNStageIntLLRInputS4xD(140)(4) <= CNStageIntLLROutputS4xD(277)(2);
  VNStageIntLLRInputS4xD(240)(4) <= CNStageIntLLROutputS4xD(277)(3);
  VNStageIntLLRInputS4xD(297)(4) <= CNStageIntLLROutputS4xD(277)(4);
  VNStageIntLLRInputS4xD(379)(2) <= CNStageIntLLROutputS4xD(277)(5);
  VNStageIntLLRInputS4xD(19)(3) <= CNStageIntLLROutputS4xD(278)(0);
  VNStageIntLLRInputS4xD(75)(4) <= CNStageIntLLROutputS4xD(278)(1);
  VNStageIntLLRInputS4xD(175)(4) <= CNStageIntLLROutputS4xD(278)(2);
  VNStageIntLLRInputS4xD(232)(3) <= CNStageIntLLROutputS4xD(278)(3);
  VNStageIntLLRInputS4xD(314)(1) <= CNStageIntLLROutputS4xD(278)(4);
  VNStageIntLLRInputS4xD(376)(3) <= CNStageIntLLROutputS4xD(278)(5);
  VNStageIntLLRInputS4xD(0)(4) <= CNStageIntLLROutputS4xD(279)(0);
  VNStageIntLLRInputS4xD(123)(3) <= CNStageIntLLROutputS4xD(279)(1);
  VNStageIntLLRInputS4xD(188)(2) <= CNStageIntLLROutputS4xD(279)(2);
  VNStageIntLLRInputS4xD(253)(3) <= CNStageIntLLROutputS4xD(279)(3);
  VNStageIntLLRInputS4xD(318)(2) <= CNStageIntLLROutputS4xD(279)(4);
  VNStageIntLLRInputS4xD(383)(4) <= CNStageIntLLROutputS4xD(279)(5);
  VNStageIntLLRInputS4xD(35)(5) <= CNStageIntLLROutputS4xD(280)(0);
  VNStageIntLLRInputS4xD(91)(5) <= CNStageIntLLROutputS4xD(280)(1);
  VNStageIntLLRInputS4xD(191)(5) <= CNStageIntLLROutputS4xD(280)(2);
  VNStageIntLLRInputS4xD(248)(5) <= CNStageIntLLROutputS4xD(280)(3);
  VNStageIntLLRInputS4xD(267)(5) <= CNStageIntLLROutputS4xD(280)(4);
  VNStageIntLLRInputS4xD(329)(5) <= CNStageIntLLROutputS4xD(280)(5);
  VNStageIntLLRInputS4xD(34)(5) <= CNStageIntLLROutputS4xD(281)(0);
  VNStageIntLLRInputS4xD(126)(4) <= CNStageIntLLROutputS4xD(281)(1);
  VNStageIntLLRInputS4xD(183)(3) <= CNStageIntLLROutputS4xD(281)(2);
  VNStageIntLLRInputS4xD(202)(4) <= CNStageIntLLROutputS4xD(281)(3);
  VNStageIntLLRInputS4xD(264)(5) <= CNStageIntLLROutputS4xD(281)(4);
  VNStageIntLLRInputS4xD(363)(4) <= CNStageIntLLROutputS4xD(281)(5);
  VNStageIntLLRInputS4xD(33)(5) <= CNStageIntLLROutputS4xD(282)(0);
  VNStageIntLLRInputS4xD(118)(4) <= CNStageIntLLROutputS4xD(282)(1);
  VNStageIntLLRInputS4xD(137)(5) <= CNStageIntLLROutputS4xD(282)(2);
  VNStageIntLLRInputS4xD(199)(5) <= CNStageIntLLROutputS4xD(282)(3);
  VNStageIntLLRInputS4xD(298)(5) <= CNStageIntLLROutputS4xD(282)(4);
  VNStageIntLLRInputS4xD(383)(5) <= CNStageIntLLROutputS4xD(282)(5);
  VNStageIntLLRInputS4xD(31)(3) <= CNStageIntLLROutputS4xD(283)(0);
  VNStageIntLLRInputS4xD(69)(5) <= CNStageIntLLROutputS4xD(283)(1);
  VNStageIntLLRInputS4xD(168)(4) <= CNStageIntLLROutputS4xD(283)(2);
  VNStageIntLLRInputS4xD(253)(4) <= CNStageIntLLROutputS4xD(283)(3);
  VNStageIntLLRInputS4xD(304)(5) <= CNStageIntLLROutputS4xD(283)(4);
  VNStageIntLLRInputS4xD(359)(5) <= CNStageIntLLROutputS4xD(283)(5);
  VNStageIntLLRInputS4xD(30)(5) <= CNStageIntLLROutputS4xD(284)(0);
  VNStageIntLLRInputS4xD(103)(5) <= CNStageIntLLROutputS4xD(284)(1);
  VNStageIntLLRInputS4xD(188)(3) <= CNStageIntLLROutputS4xD(284)(2);
  VNStageIntLLRInputS4xD(239)(5) <= CNStageIntLLROutputS4xD(284)(3);
  VNStageIntLLRInputS4xD(294)(5) <= CNStageIntLLROutputS4xD(284)(4);
  VNStageIntLLRInputS4xD(325)(5) <= CNStageIntLLROutputS4xD(284)(5);
  VNStageIntLLRInputS4xD(27)(4) <= CNStageIntLLROutputS4xD(285)(0);
  VNStageIntLLRInputS4xD(99)(5) <= CNStageIntLLROutputS4xD(285)(1);
  VNStageIntLLRInputS4xD(130)(5) <= CNStageIntLLROutputS4xD(285)(2);
  VNStageIntLLRInputS4xD(241)(4) <= CNStageIntLLROutputS4xD(285)(3);
  VNStageIntLLRInputS4xD(273)(4) <= CNStageIntLLROutputS4xD(285)(4);
  VNStageIntLLRInputS4xD(361)(5) <= CNStageIntLLROutputS4xD(285)(5);
  VNStageIntLLRInputS4xD(26)(5) <= CNStageIntLLROutputS4xD(286)(0);
  VNStageIntLLRInputS4xD(65)(4) <= CNStageIntLLROutputS4xD(286)(1);
  VNStageIntLLRInputS4xD(176)(5) <= CNStageIntLLROutputS4xD(286)(2);
  VNStageIntLLRInputS4xD(208)(4) <= CNStageIntLLROutputS4xD(286)(3);
  VNStageIntLLRInputS4xD(296)(4) <= CNStageIntLLROutputS4xD(286)(4);
  VNStageIntLLRInputS4xD(334)(3) <= CNStageIntLLROutputS4xD(286)(5);
  VNStageIntLLRInputS4xD(25)(4) <= CNStageIntLLROutputS4xD(287)(0);
  VNStageIntLLRInputS4xD(111)(5) <= CNStageIntLLROutputS4xD(287)(1);
  VNStageIntLLRInputS4xD(143)(5) <= CNStageIntLLROutputS4xD(287)(2);
  VNStageIntLLRInputS4xD(231)(4) <= CNStageIntLLROutputS4xD(287)(3);
  VNStageIntLLRInputS4xD(269)(4) <= CNStageIntLLROutputS4xD(287)(4);
  VNStageIntLLRInputS4xD(381)(4) <= CNStageIntLLROutputS4xD(287)(5);
  VNStageIntLLRInputS4xD(24)(5) <= CNStageIntLLROutputS4xD(288)(0);
  VNStageIntLLRInputS4xD(78)(5) <= CNStageIntLLROutputS4xD(288)(1);
  VNStageIntLLRInputS4xD(166)(4) <= CNStageIntLLROutputS4xD(288)(2);
  VNStageIntLLRInputS4xD(204)(5) <= CNStageIntLLROutputS4xD(288)(3);
  VNStageIntLLRInputS4xD(316)(3) <= CNStageIntLLROutputS4xD(288)(4);
  VNStageIntLLRInputS4xD(321)(5) <= CNStageIntLLROutputS4xD(288)(5);
  VNStageIntLLRInputS4xD(23)(5) <= CNStageIntLLROutputS4xD(289)(0);
  VNStageIntLLRInputS4xD(101)(5) <= CNStageIntLLROutputS4xD(289)(1);
  VNStageIntLLRInputS4xD(139)(5) <= CNStageIntLLROutputS4xD(289)(2);
  VNStageIntLLRInputS4xD(251)(3) <= CNStageIntLLROutputS4xD(289)(3);
  VNStageIntLLRInputS4xD(319)(5) <= CNStageIntLLROutputS4xD(289)(4);
  VNStageIntLLRInputS4xD(362)(5) <= CNStageIntLLROutputS4xD(289)(5);
  VNStageIntLLRInputS4xD(22)(5) <= CNStageIntLLROutputS4xD(290)(0);
  VNStageIntLLRInputS4xD(74)(4) <= CNStageIntLLROutputS4xD(290)(1);
  VNStageIntLLRInputS4xD(186)(4) <= CNStageIntLLROutputS4xD(290)(2);
  VNStageIntLLRInputS4xD(254)(3) <= CNStageIntLLROutputS4xD(290)(3);
  VNStageIntLLRInputS4xD(297)(5) <= CNStageIntLLROutputS4xD(290)(4);
  VNStageIntLLRInputS4xD(337)(5) <= CNStageIntLLROutputS4xD(290)(5);
  VNStageIntLLRInputS4xD(21)(5) <= CNStageIntLLROutputS4xD(291)(0);
  VNStageIntLLRInputS4xD(121)(4) <= CNStageIntLLROutputS4xD(291)(1);
  VNStageIntLLRInputS4xD(189)(4) <= CNStageIntLLROutputS4xD(291)(2);
  VNStageIntLLRInputS4xD(232)(4) <= CNStageIntLLROutputS4xD(291)(3);
  VNStageIntLLRInputS4xD(272)(5) <= CNStageIntLLROutputS4xD(291)(4);
  VNStageIntLLRInputS4xD(335)(5) <= CNStageIntLLROutputS4xD(291)(5);
  VNStageIntLLRInputS4xD(20)(3) <= CNStageIntLLROutputS4xD(292)(0);
  VNStageIntLLRInputS4xD(124)(3) <= CNStageIntLLROutputS4xD(292)(1);
  VNStageIntLLRInputS4xD(167)(5) <= CNStageIntLLROutputS4xD(292)(2);
  VNStageIntLLRInputS4xD(207)(4) <= CNStageIntLLROutputS4xD(292)(3);
  VNStageIntLLRInputS4xD(270)(5) <= CNStageIntLLROutputS4xD(292)(4);
  VNStageIntLLRInputS4xD(360)(5) <= CNStageIntLLROutputS4xD(292)(5);
  VNStageIntLLRInputS4xD(18)(5) <= CNStageIntLLROutputS4xD(293)(0);
  VNStageIntLLRInputS4xD(77)(3) <= CNStageIntLLROutputS4xD(293)(1);
  VNStageIntLLRInputS4xD(140)(5) <= CNStageIntLLROutputS4xD(293)(2);
  VNStageIntLLRInputS4xD(230)(4) <= CNStageIntLLROutputS4xD(293)(3);
  VNStageIntLLRInputS4xD(303)(5) <= CNStageIntLLROutputS4xD(293)(4);
  VNStageIntLLRInputS4xD(348)(5) <= CNStageIntLLROutputS4xD(293)(5);
  VNStageIntLLRInputS4xD(17)(5) <= CNStageIntLLROutputS4xD(294)(0);
  VNStageIntLLRInputS4xD(75)(5) <= CNStageIntLLROutputS4xD(294)(1);
  VNStageIntLLRInputS4xD(165)(4) <= CNStageIntLLROutputS4xD(294)(2);
  VNStageIntLLRInputS4xD(238)(5) <= CNStageIntLLROutputS4xD(294)(3);
  VNStageIntLLRInputS4xD(283)(5) <= CNStageIntLLROutputS4xD(294)(4);
  VNStageIntLLRInputS4xD(342)(4) <= CNStageIntLLROutputS4xD(294)(5);
  VNStageIntLLRInputS4xD(16)(4) <= CNStageIntLLROutputS4xD(295)(0);
  VNStageIntLLRInputS4xD(100)(5) <= CNStageIntLLROutputS4xD(295)(1);
  VNStageIntLLRInputS4xD(173)(5) <= CNStageIntLLROutputS4xD(295)(2);
  VNStageIntLLRInputS4xD(218)(5) <= CNStageIntLLROutputS4xD(295)(3);
  VNStageIntLLRInputS4xD(277)(5) <= CNStageIntLLROutputS4xD(295)(4);
  VNStageIntLLRInputS4xD(320)(3) <= CNStageIntLLROutputS4xD(295)(5);
  VNStageIntLLRInputS4xD(15)(5) <= CNStageIntLLROutputS4xD(296)(0);
  VNStageIntLLRInputS4xD(108)(5) <= CNStageIntLLROutputS4xD(296)(1);
  VNStageIntLLRInputS4xD(153)(5) <= CNStageIntLLROutputS4xD(296)(2);
  VNStageIntLLRInputS4xD(212)(4) <= CNStageIntLLROutputS4xD(296)(3);
  VNStageIntLLRInputS4xD(256)(4) <= CNStageIntLLROutputS4xD(296)(4);
  VNStageIntLLRInputS4xD(341)(5) <= CNStageIntLLROutputS4xD(296)(5);
  VNStageIntLLRInputS4xD(14)(5) <= CNStageIntLLROutputS4xD(297)(0);
  VNStageIntLLRInputS4xD(88)(5) <= CNStageIntLLROutputS4xD(297)(1);
  VNStageIntLLRInputS4xD(147)(5) <= CNStageIntLLROutputS4xD(297)(2);
  VNStageIntLLRInputS4xD(192)(5) <= CNStageIntLLROutputS4xD(297)(3);
  VNStageIntLLRInputS4xD(276)(5) <= CNStageIntLLROutputS4xD(297)(4);
  VNStageIntLLRInputS4xD(346)(5) <= CNStageIntLLROutputS4xD(297)(5);
  VNStageIntLLRInputS4xD(13)(4) <= CNStageIntLLROutputS4xD(298)(0);
  VNStageIntLLRInputS4xD(82)(5) <= CNStageIntLLROutputS4xD(298)(1);
  VNStageIntLLRInputS4xD(128)(5) <= CNStageIntLLROutputS4xD(298)(2);
  VNStageIntLLRInputS4xD(211)(5) <= CNStageIntLLROutputS4xD(298)(3);
  VNStageIntLLRInputS4xD(281)(5) <= CNStageIntLLROutputS4xD(298)(4);
  VNStageIntLLRInputS4xD(365)(5) <= CNStageIntLLROutputS4xD(298)(5);
  VNStageIntLLRInputS4xD(12)(5) <= CNStageIntLLROutputS4xD(299)(0);
  VNStageIntLLRInputS4xD(64)(4) <= CNStageIntLLROutputS4xD(299)(1);
  VNStageIntLLRInputS4xD(146)(4) <= CNStageIntLLROutputS4xD(299)(2);
  VNStageIntLLRInputS4xD(216)(5) <= CNStageIntLLROutputS4xD(299)(3);
  VNStageIntLLRInputS4xD(300)(4) <= CNStageIntLLROutputS4xD(299)(4);
  VNStageIntLLRInputS4xD(356)(4) <= CNStageIntLLROutputS4xD(299)(5);
  VNStageIntLLRInputS4xD(9)(5) <= CNStageIntLLROutputS4xD(300)(0);
  VNStageIntLLRInputS4xD(105)(4) <= CNStageIntLLROutputS4xD(300)(1);
  VNStageIntLLRInputS4xD(161)(5) <= CNStageIntLLROutputS4xD(300)(2);
  VNStageIntLLRInputS4xD(200)(5) <= CNStageIntLLROutputS4xD(300)(3);
  VNStageIntLLRInputS4xD(266)(4) <= CNStageIntLLROutputS4xD(300)(4);
  VNStageIntLLRInputS4xD(355)(5) <= CNStageIntLLROutputS4xD(300)(5);
  VNStageIntLLRInputS4xD(7)(5) <= CNStageIntLLROutputS4xD(301)(0);
  VNStageIntLLRInputS4xD(70)(5) <= CNStageIntLLROutputS4xD(301)(1);
  VNStageIntLLRInputS4xD(136)(5) <= CNStageIntLLROutputS4xD(301)(2);
  VNStageIntLLRInputS4xD(225)(5) <= CNStageIntLLROutputS4xD(301)(3);
  VNStageIntLLRInputS4xD(311)(4) <= CNStageIntLLROutputS4xD(301)(4);
  VNStageIntLLRInputS4xD(372)(4) <= CNStageIntLLROutputS4xD(301)(5);
  VNStageIntLLRInputS4xD(6)(5) <= CNStageIntLLROutputS4xD(302)(0);
  VNStageIntLLRInputS4xD(71)(4) <= CNStageIntLLROutputS4xD(302)(1);
  VNStageIntLLRInputS4xD(160)(5) <= CNStageIntLLROutputS4xD(302)(2);
  VNStageIntLLRInputS4xD(246)(5) <= CNStageIntLLROutputS4xD(302)(3);
  VNStageIntLLRInputS4xD(307)(5) <= CNStageIntLLROutputS4xD(302)(4);
  VNStageIntLLRInputS4xD(324)(5) <= CNStageIntLLROutputS4xD(302)(5);
  VNStageIntLLRInputS4xD(5)(5) <= CNStageIntLLROutputS4xD(303)(0);
  VNStageIntLLRInputS4xD(95)(5) <= CNStageIntLLROutputS4xD(303)(1);
  VNStageIntLLRInputS4xD(181)(5) <= CNStageIntLLROutputS4xD(303)(2);
  VNStageIntLLRInputS4xD(242)(5) <= CNStageIntLLROutputS4xD(303)(3);
  VNStageIntLLRInputS4xD(259)(3) <= CNStageIntLLROutputS4xD(303)(4);
  VNStageIntLLRInputS4xD(350)(5) <= CNStageIntLLROutputS4xD(303)(5);
  VNStageIntLLRInputS4xD(4)(4) <= CNStageIntLLROutputS4xD(304)(0);
  VNStageIntLLRInputS4xD(116)(4) <= CNStageIntLLROutputS4xD(304)(1);
  VNStageIntLLRInputS4xD(177)(5) <= CNStageIntLLROutputS4xD(304)(2);
  VNStageIntLLRInputS4xD(194)(5) <= CNStageIntLLROutputS4xD(304)(3);
  VNStageIntLLRInputS4xD(285)(5) <= CNStageIntLLROutputS4xD(304)(4);
  VNStageIntLLRInputS4xD(326)(4) <= CNStageIntLLROutputS4xD(304)(5);
  VNStageIntLLRInputS4xD(3)(4) <= CNStageIntLLROutputS4xD(305)(0);
  VNStageIntLLRInputS4xD(112)(5) <= CNStageIntLLROutputS4xD(305)(1);
  VNStageIntLLRInputS4xD(129)(5) <= CNStageIntLLROutputS4xD(305)(2);
  VNStageIntLLRInputS4xD(220)(5) <= CNStageIntLLROutputS4xD(305)(3);
  VNStageIntLLRInputS4xD(261)(4) <= CNStageIntLLROutputS4xD(305)(4);
  VNStageIntLLRInputS4xD(358)(4) <= CNStageIntLLROutputS4xD(305)(5);
  VNStageIntLLRInputS4xD(2)(5) <= CNStageIntLLROutputS4xD(306)(0);
  VNStageIntLLRInputS4xD(127)(5) <= CNStageIntLLROutputS4xD(306)(1);
  VNStageIntLLRInputS4xD(155)(5) <= CNStageIntLLROutputS4xD(306)(2);
  VNStageIntLLRInputS4xD(196)(5) <= CNStageIntLLROutputS4xD(306)(3);
  VNStageIntLLRInputS4xD(293)(4) <= CNStageIntLLROutputS4xD(306)(4);
  VNStageIntLLRInputS4xD(374)(5) <= CNStageIntLLROutputS4xD(306)(5);
  VNStageIntLLRInputS4xD(1)(4) <= CNStageIntLLROutputS4xD(307)(0);
  VNStageIntLLRInputS4xD(90)(5) <= CNStageIntLLROutputS4xD(307)(1);
  VNStageIntLLRInputS4xD(131)(4) <= CNStageIntLLROutputS4xD(307)(2);
  VNStageIntLLRInputS4xD(228)(5) <= CNStageIntLLROutputS4xD(307)(3);
  VNStageIntLLRInputS4xD(309)(5) <= CNStageIntLLROutputS4xD(307)(4);
  VNStageIntLLRInputS4xD(344)(5) <= CNStageIntLLROutputS4xD(307)(5);
  VNStageIntLLRInputS4xD(62)(4) <= CNStageIntLLROutputS4xD(308)(0);
  VNStageIntLLRInputS4xD(98)(4) <= CNStageIntLLROutputS4xD(308)(1);
  VNStageIntLLRInputS4xD(179)(5) <= CNStageIntLLROutputS4xD(308)(2);
  VNStageIntLLRInputS4xD(214)(5) <= CNStageIntLLROutputS4xD(308)(3);
  VNStageIntLLRInputS4xD(288)(5) <= CNStageIntLLROutputS4xD(308)(4);
  VNStageIntLLRInputS4xD(366)(5) <= CNStageIntLLROutputS4xD(308)(5);
  VNStageIntLLRInputS4xD(61)(4) <= CNStageIntLLROutputS4xD(309)(0);
  VNStageIntLLRInputS4xD(114)(5) <= CNStageIntLLROutputS4xD(309)(1);
  VNStageIntLLRInputS4xD(149)(5) <= CNStageIntLLROutputS4xD(309)(2);
  VNStageIntLLRInputS4xD(223)(5) <= CNStageIntLLROutputS4xD(309)(3);
  VNStageIntLLRInputS4xD(301)(5) <= CNStageIntLLROutputS4xD(309)(4);
  VNStageIntLLRInputS4xD(345)(4) <= CNStageIntLLROutputS4xD(309)(5);
  VNStageIntLLRInputS4xD(60)(4) <= CNStageIntLLROutputS4xD(310)(0);
  VNStageIntLLRInputS4xD(84)(4) <= CNStageIntLLROutputS4xD(310)(1);
  VNStageIntLLRInputS4xD(158)(5) <= CNStageIntLLROutputS4xD(310)(2);
  VNStageIntLLRInputS4xD(236)(5) <= CNStageIntLLROutputS4xD(310)(3);
  VNStageIntLLRInputS4xD(280)(5) <= CNStageIntLLROutputS4xD(310)(4);
  VNStageIntLLRInputS4xD(373)(3) <= CNStageIntLLROutputS4xD(310)(5);
  VNStageIntLLRInputS4xD(59)(3) <= CNStageIntLLROutputS4xD(311)(0);
  VNStageIntLLRInputS4xD(93)(5) <= CNStageIntLLROutputS4xD(311)(1);
  VNStageIntLLRInputS4xD(171)(3) <= CNStageIntLLROutputS4xD(311)(2);
  VNStageIntLLRInputS4xD(215)(5) <= CNStageIntLLROutputS4xD(311)(3);
  VNStageIntLLRInputS4xD(308)(3) <= CNStageIntLLROutputS4xD(311)(4);
  VNStageIntLLRInputS4xD(375)(4) <= CNStageIntLLROutputS4xD(311)(5);
  VNStageIntLLRInputS4xD(58)(3) <= CNStageIntLLROutputS4xD(312)(0);
  VNStageIntLLRInputS4xD(106)(4) <= CNStageIntLLROutputS4xD(312)(1);
  VNStageIntLLRInputS4xD(150)(4) <= CNStageIntLLROutputS4xD(312)(2);
  VNStageIntLLRInputS4xD(243)(5) <= CNStageIntLLROutputS4xD(312)(3);
  VNStageIntLLRInputS4xD(310)(4) <= CNStageIntLLROutputS4xD(312)(4);
  VNStageIntLLRInputS4xD(357)(5) <= CNStageIntLLROutputS4xD(312)(5);
  VNStageIntLLRInputS4xD(57)(4) <= CNStageIntLLROutputS4xD(313)(0);
  VNStageIntLLRInputS4xD(85)(4) <= CNStageIntLLROutputS4xD(313)(1);
  VNStageIntLLRInputS4xD(178)(4) <= CNStageIntLLROutputS4xD(313)(2);
  VNStageIntLLRInputS4xD(245)(5) <= CNStageIntLLROutputS4xD(313)(3);
  VNStageIntLLRInputS4xD(292)(5) <= CNStageIntLLROutputS4xD(313)(4);
  VNStageIntLLRInputS4xD(364)(5) <= CNStageIntLLROutputS4xD(313)(5);
  VNStageIntLLRInputS4xD(56)(5) <= CNStageIntLLROutputS4xD(314)(0);
  VNStageIntLLRInputS4xD(113)(5) <= CNStageIntLLROutputS4xD(314)(1);
  VNStageIntLLRInputS4xD(180)(3) <= CNStageIntLLROutputS4xD(314)(2);
  VNStageIntLLRInputS4xD(227)(5) <= CNStageIntLLROutputS4xD(314)(3);
  VNStageIntLLRInputS4xD(299)(4) <= CNStageIntLLROutputS4xD(314)(4);
  VNStageIntLLRInputS4xD(328)(3) <= CNStageIntLLROutputS4xD(314)(5);
  VNStageIntLLRInputS4xD(55)(5) <= CNStageIntLLROutputS4xD(315)(0);
  VNStageIntLLRInputS4xD(115)(5) <= CNStageIntLLROutputS4xD(315)(1);
  VNStageIntLLRInputS4xD(162)(5) <= CNStageIntLLROutputS4xD(315)(2);
  VNStageIntLLRInputS4xD(234)(5) <= CNStageIntLLROutputS4xD(315)(3);
  VNStageIntLLRInputS4xD(263)(5) <= CNStageIntLLROutputS4xD(315)(4);
  VNStageIntLLRInputS4xD(379)(3) <= CNStageIntLLROutputS4xD(315)(5);
  VNStageIntLLRInputS4xD(54)(4) <= CNStageIntLLROutputS4xD(316)(0);
  VNStageIntLLRInputS4xD(97)(5) <= CNStageIntLLROutputS4xD(316)(1);
  VNStageIntLLRInputS4xD(169)(5) <= CNStageIntLLROutputS4xD(316)(2);
  VNStageIntLLRInputS4xD(198)(5) <= CNStageIntLLROutputS4xD(316)(3);
  VNStageIntLLRInputS4xD(314)(2) <= CNStageIntLLROutputS4xD(316)(4);
  VNStageIntLLRInputS4xD(322)(4) <= CNStageIntLLROutputS4xD(316)(5);
  VNStageIntLLRInputS4xD(53)(4) <= CNStageIntLLROutputS4xD(317)(0);
  VNStageIntLLRInputS4xD(104)(5) <= CNStageIntLLROutputS4xD(317)(1);
  VNStageIntLLRInputS4xD(133)(3) <= CNStageIntLLROutputS4xD(317)(2);
  VNStageIntLLRInputS4xD(249)(3) <= CNStageIntLLROutputS4xD(317)(3);
  VNStageIntLLRInputS4xD(257)(5) <= CNStageIntLLROutputS4xD(317)(4);
  VNStageIntLLRInputS4xD(380)(4) <= CNStageIntLLROutputS4xD(317)(5);
  VNStageIntLLRInputS4xD(52)(3) <= CNStageIntLLROutputS4xD(318)(0);
  VNStageIntLLRInputS4xD(68)(4) <= CNStageIntLLROutputS4xD(318)(1);
  VNStageIntLLRInputS4xD(184)(5) <= CNStageIntLLROutputS4xD(318)(2);
  VNStageIntLLRInputS4xD(255)(5) <= CNStageIntLLROutputS4xD(318)(3);
  VNStageIntLLRInputS4xD(315)(4) <= CNStageIntLLROutputS4xD(318)(4);
  VNStageIntLLRInputS4xD(327)(5) <= CNStageIntLLROutputS4xD(318)(5);
  VNStageIntLLRInputS4xD(51)(4) <= CNStageIntLLROutputS4xD(319)(0);
  VNStageIntLLRInputS4xD(119)(4) <= CNStageIntLLROutputS4xD(319)(1);
  VNStageIntLLRInputS4xD(190)(3) <= CNStageIntLLROutputS4xD(319)(2);
  VNStageIntLLRInputS4xD(250)(3) <= CNStageIntLLROutputS4xD(319)(3);
  VNStageIntLLRInputS4xD(262)(4) <= CNStageIntLLROutputS4xD(319)(4);
  VNStageIntLLRInputS4xD(349)(4) <= CNStageIntLLROutputS4xD(319)(5);
  VNStageIntLLRInputS4xD(50)(5) <= CNStageIntLLROutputS4xD(320)(0);
  VNStageIntLLRInputS4xD(125)(2) <= CNStageIntLLROutputS4xD(320)(1);
  VNStageIntLLRInputS4xD(185)(2) <= CNStageIntLLROutputS4xD(320)(2);
  VNStageIntLLRInputS4xD(197)(5) <= CNStageIntLLROutputS4xD(320)(3);
  VNStageIntLLRInputS4xD(284)(5) <= CNStageIntLLROutputS4xD(320)(4);
  VNStageIntLLRInputS4xD(367)(5) <= CNStageIntLLROutputS4xD(320)(5);
  VNStageIntLLRInputS4xD(49)(5) <= CNStageIntLLROutputS4xD(321)(0);
  VNStageIntLLRInputS4xD(120)(2) <= CNStageIntLLROutputS4xD(321)(1);
  VNStageIntLLRInputS4xD(132)(4) <= CNStageIntLLROutputS4xD(321)(2);
  VNStageIntLLRInputS4xD(219)(4) <= CNStageIntLLROutputS4xD(321)(3);
  VNStageIntLLRInputS4xD(302)(5) <= CNStageIntLLROutputS4xD(321)(4);
  VNStageIntLLRInputS4xD(352)(5) <= CNStageIntLLROutputS4xD(321)(5);
  VNStageIntLLRInputS4xD(48)(2) <= CNStageIntLLROutputS4xD(322)(0);
  VNStageIntLLRInputS4xD(67)(2) <= CNStageIntLLROutputS4xD(322)(1);
  VNStageIntLLRInputS4xD(154)(4) <= CNStageIntLLROutputS4xD(322)(2);
  VNStageIntLLRInputS4xD(237)(4) <= CNStageIntLLROutputS4xD(322)(3);
  VNStageIntLLRInputS4xD(287)(5) <= CNStageIntLLROutputS4xD(322)(4);
  VNStageIntLLRInputS4xD(339)(5) <= CNStageIntLLROutputS4xD(322)(5);
  VNStageIntLLRInputS4xD(46)(5) <= CNStageIntLLROutputS4xD(323)(0);
  VNStageIntLLRInputS4xD(107)(4) <= CNStageIntLLROutputS4xD(323)(1);
  VNStageIntLLRInputS4xD(157)(4) <= CNStageIntLLROutputS4xD(323)(2);
  VNStageIntLLRInputS4xD(209)(4) <= CNStageIntLLROutputS4xD(323)(3);
  VNStageIntLLRInputS4xD(305)(5) <= CNStageIntLLROutputS4xD(323)(4);
  VNStageIntLLRInputS4xD(382)(4) <= CNStageIntLLROutputS4xD(323)(5);
  VNStageIntLLRInputS4xD(45)(5) <= CNStageIntLLROutputS4xD(324)(0);
  VNStageIntLLRInputS4xD(92)(5) <= CNStageIntLLROutputS4xD(324)(1);
  VNStageIntLLRInputS4xD(144)(5) <= CNStageIntLLROutputS4xD(324)(2);
  VNStageIntLLRInputS4xD(240)(5) <= CNStageIntLLROutputS4xD(324)(3);
  VNStageIntLLRInputS4xD(317)(2) <= CNStageIntLLROutputS4xD(324)(4);
  VNStageIntLLRInputS4xD(333)(4) <= CNStageIntLLROutputS4xD(324)(5);
  VNStageIntLLRInputS4xD(44)(5) <= CNStageIntLLROutputS4xD(325)(0);
  VNStageIntLLRInputS4xD(79)(4) <= CNStageIntLLROutputS4xD(325)(1);
  VNStageIntLLRInputS4xD(175)(5) <= CNStageIntLLROutputS4xD(325)(2);
  VNStageIntLLRInputS4xD(252)(4) <= CNStageIntLLROutputS4xD(325)(3);
  VNStageIntLLRInputS4xD(268)(5) <= CNStageIntLLROutputS4xD(325)(4);
  VNStageIntLLRInputS4xD(377)(3) <= CNStageIntLLROutputS4xD(325)(5);
  VNStageIntLLRInputS4xD(43)(4) <= CNStageIntLLROutputS4xD(326)(0);
  VNStageIntLLRInputS4xD(110)(5) <= CNStageIntLLROutputS4xD(326)(1);
  VNStageIntLLRInputS4xD(187)(4) <= CNStageIntLLROutputS4xD(326)(2);
  VNStageIntLLRInputS4xD(203)(5) <= CNStageIntLLROutputS4xD(326)(3);
  VNStageIntLLRInputS4xD(312)(4) <= CNStageIntLLROutputS4xD(326)(4);
  VNStageIntLLRInputS4xD(354)(4) <= CNStageIntLLROutputS4xD(326)(5);
  VNStageIntLLRInputS4xD(42)(5) <= CNStageIntLLROutputS4xD(327)(0);
  VNStageIntLLRInputS4xD(122)(4) <= CNStageIntLLROutputS4xD(327)(1);
  VNStageIntLLRInputS4xD(138)(5) <= CNStageIntLLROutputS4xD(327)(2);
  VNStageIntLLRInputS4xD(247)(5) <= CNStageIntLLROutputS4xD(327)(3);
  VNStageIntLLRInputS4xD(289)(5) <= CNStageIntLLROutputS4xD(327)(4);
  VNStageIntLLRInputS4xD(343)(5) <= CNStageIntLLROutputS4xD(327)(5);
  VNStageIntLLRInputS4xD(41)(5) <= CNStageIntLLROutputS4xD(328)(0);
  VNStageIntLLRInputS4xD(73)(4) <= CNStageIntLLROutputS4xD(328)(1);
  VNStageIntLLRInputS4xD(182)(5) <= CNStageIntLLROutputS4xD(328)(2);
  VNStageIntLLRInputS4xD(224)(5) <= CNStageIntLLROutputS4xD(328)(3);
  VNStageIntLLRInputS4xD(278)(4) <= CNStageIntLLROutputS4xD(328)(4);
  VNStageIntLLRInputS4xD(347)(5) <= CNStageIntLLROutputS4xD(328)(5);
  VNStageIntLLRInputS4xD(39)(5) <= CNStageIntLLROutputS4xD(329)(0);
  VNStageIntLLRInputS4xD(94)(3) <= CNStageIntLLROutputS4xD(329)(1);
  VNStageIntLLRInputS4xD(148)(5) <= CNStageIntLLROutputS4xD(329)(2);
  VNStageIntLLRInputS4xD(217)(5) <= CNStageIntLLROutputS4xD(329)(3);
  VNStageIntLLRInputS4xD(275)(4) <= CNStageIntLLROutputS4xD(329)(4);
  VNStageIntLLRInputS4xD(351)(4) <= CNStageIntLLROutputS4xD(329)(5);
  VNStageIntLLRInputS4xD(38)(5) <= CNStageIntLLROutputS4xD(330)(0);
  VNStageIntLLRInputS4xD(83)(5) <= CNStageIntLLROutputS4xD(330)(1);
  VNStageIntLLRInputS4xD(152)(5) <= CNStageIntLLROutputS4xD(330)(2);
  VNStageIntLLRInputS4xD(210)(5) <= CNStageIntLLROutputS4xD(330)(3);
  VNStageIntLLRInputS4xD(286)(5) <= CNStageIntLLROutputS4xD(330)(4);
  VNStageIntLLRInputS4xD(323)(4) <= CNStageIntLLROutputS4xD(330)(5);
  VNStageIntLLRInputS4xD(37)(5) <= CNStageIntLLROutputS4xD(331)(0);
  VNStageIntLLRInputS4xD(87)(5) <= CNStageIntLLROutputS4xD(331)(1);
  VNStageIntLLRInputS4xD(145)(5) <= CNStageIntLLROutputS4xD(331)(2);
  VNStageIntLLRInputS4xD(221)(5) <= CNStageIntLLROutputS4xD(331)(3);
  VNStageIntLLRInputS4xD(258)(2) <= CNStageIntLLROutputS4xD(331)(4);
  VNStageIntLLRInputS4xD(378)(4) <= CNStageIntLLROutputS4xD(331)(5);
  VNStageIntLLRInputS4xD(0)(5) <= CNStageIntLLROutputS4xD(332)(0);
  VNStageIntLLRInputS4xD(76)(5) <= CNStageIntLLROutputS4xD(332)(1);
  VNStageIntLLRInputS4xD(141)(3) <= CNStageIntLLROutputS4xD(332)(2);
  VNStageIntLLRInputS4xD(206)(3) <= CNStageIntLLROutputS4xD(332)(3);
  VNStageIntLLRInputS4xD(271)(4) <= CNStageIntLLROutputS4xD(332)(4);
  VNStageIntLLRInputS4xD(336)(4) <= CNStageIntLLROutputS4xD(332)(5);
  VNStageIntLLRInputS4xD(28)(5) <= CNStageIntLLROutputS4xD(333)(0);
  VNStageIntLLRInputS4xD(106)(5) <= CNStageIntLLROutputS4xD(333)(1);
  VNStageIntLLRInputS4xD(144)(6) <= CNStageIntLLROutputS4xD(333)(2);
  VNStageIntLLRInputS4xD(193)(4) <= CNStageIntLLROutputS4xD(333)(3);
  VNStageIntLLRInputS4xD(261)(5) <= CNStageIntLLROutputS4xD(333)(4);
  VNStageIntLLRInputS4xD(367)(6) <= CNStageIntLLROutputS4xD(333)(5);
  VNStageIntLLRInputS4xD(26)(6) <= CNStageIntLLROutputS4xD(334)(0);
  VNStageIntLLRInputS4xD(126)(5) <= CNStageIntLLROutputS4xD(334)(1);
  VNStageIntLLRInputS4xD(131)(5) <= CNStageIntLLROutputS4xD(334)(2);
  VNStageIntLLRInputS4xD(237)(5) <= CNStageIntLLROutputS4xD(334)(3);
  VNStageIntLLRInputS4xD(277)(6) <= CNStageIntLLROutputS4xD(334)(4);
  VNStageIntLLRInputS4xD(340)(5) <= CNStageIntLLROutputS4xD(334)(5);
  VNStageIntLLRInputS4xD(24)(6) <= CNStageIntLLROutputS4xD(335)(0);
  VNStageIntLLRInputS4xD(107)(5) <= CNStageIntLLROutputS4xD(335)(1);
  VNStageIntLLRInputS4xD(147)(6) <= CNStageIntLLROutputS4xD(335)(2);
  VNStageIntLLRInputS4xD(210)(6) <= CNStageIntLLROutputS4xD(335)(3);
  VNStageIntLLRInputS4xD(300)(5) <= CNStageIntLLROutputS4xD(335)(4);
  VNStageIntLLRInputS4xD(373)(4) <= CNStageIntLLROutputS4xD(335)(5);
  VNStageIntLLRInputS4xD(23)(6) <= CNStageIntLLROutputS4xD(336)(0);
  VNStageIntLLRInputS4xD(82)(6) <= CNStageIntLLROutputS4xD(336)(1);
  VNStageIntLLRInputS4xD(145)(6) <= CNStageIntLLROutputS4xD(336)(2);
  VNStageIntLLRInputS4xD(235)(4) <= CNStageIntLLROutputS4xD(336)(3);
  VNStageIntLLRInputS4xD(308)(4) <= CNStageIntLLROutputS4xD(336)(4);
  VNStageIntLLRInputS4xD(353)(5) <= CNStageIntLLROutputS4xD(336)(5);
  VNStageIntLLRInputS4xD(22)(6) <= CNStageIntLLROutputS4xD(337)(0);
  VNStageIntLLRInputS4xD(80)(5) <= CNStageIntLLROutputS4xD(337)(1);
  VNStageIntLLRInputS4xD(170)(4) <= CNStageIntLLROutputS4xD(337)(2);
  VNStageIntLLRInputS4xD(243)(6) <= CNStageIntLLROutputS4xD(337)(3);
  VNStageIntLLRInputS4xD(288)(6) <= CNStageIntLLROutputS4xD(337)(4);
  VNStageIntLLRInputS4xD(347)(6) <= CNStageIntLLROutputS4xD(337)(5);
  VNStageIntLLRInputS4xD(21)(6) <= CNStageIntLLROutputS4xD(338)(0);
  VNStageIntLLRInputS4xD(105)(5) <= CNStageIntLLROutputS4xD(338)(1);
  VNStageIntLLRInputS4xD(178)(5) <= CNStageIntLLROutputS4xD(338)(2);
  VNStageIntLLRInputS4xD(223)(6) <= CNStageIntLLROutputS4xD(338)(3);
  VNStageIntLLRInputS4xD(282)(5) <= CNStageIntLLROutputS4xD(338)(4);
  VNStageIntLLRInputS4xD(320)(4) <= CNStageIntLLROutputS4xD(338)(5);
  VNStageIntLLRInputS4xD(20)(4) <= CNStageIntLLROutputS4xD(339)(0);
  VNStageIntLLRInputS4xD(113)(6) <= CNStageIntLLROutputS4xD(339)(1);
  VNStageIntLLRInputS4xD(158)(6) <= CNStageIntLLROutputS4xD(339)(2);
  VNStageIntLLRInputS4xD(217)(6) <= CNStageIntLLROutputS4xD(339)(3);
  VNStageIntLLRInputS4xD(256)(5) <= CNStageIntLLROutputS4xD(339)(4);
  VNStageIntLLRInputS4xD(346)(6) <= CNStageIntLLROutputS4xD(339)(5);
  VNStageIntLLRInputS4xD(19)(4) <= CNStageIntLLROutputS4xD(340)(0);
  VNStageIntLLRInputS4xD(93)(6) <= CNStageIntLLROutputS4xD(340)(1);
  VNStageIntLLRInputS4xD(152)(6) <= CNStageIntLLROutputS4xD(340)(2);
  VNStageIntLLRInputS4xD(192)(6) <= CNStageIntLLROutputS4xD(340)(3);
  VNStageIntLLRInputS4xD(281)(6) <= CNStageIntLLROutputS4xD(340)(4);
  VNStageIntLLRInputS4xD(351)(5) <= CNStageIntLLROutputS4xD(340)(5);
  VNStageIntLLRInputS4xD(18)(6) <= CNStageIntLLROutputS4xD(341)(0);
  VNStageIntLLRInputS4xD(87)(6) <= CNStageIntLLROutputS4xD(341)(1);
  VNStageIntLLRInputS4xD(128)(6) <= CNStageIntLLROutputS4xD(341)(2);
  VNStageIntLLRInputS4xD(216)(6) <= CNStageIntLLROutputS4xD(341)(3);
  VNStageIntLLRInputS4xD(286)(6) <= CNStageIntLLROutputS4xD(341)(4);
  VNStageIntLLRInputS4xD(370)(4) <= CNStageIntLLROutputS4xD(341)(5);
  VNStageIntLLRInputS4xD(17)(6) <= CNStageIntLLROutputS4xD(342)(0);
  VNStageIntLLRInputS4xD(64)(5) <= CNStageIntLLROutputS4xD(342)(1);
  VNStageIntLLRInputS4xD(151)(5) <= CNStageIntLLROutputS4xD(342)(2);
  VNStageIntLLRInputS4xD(221)(6) <= CNStageIntLLROutputS4xD(342)(3);
  VNStageIntLLRInputS4xD(305)(6) <= CNStageIntLLROutputS4xD(342)(4);
  VNStageIntLLRInputS4xD(361)(6) <= CNStageIntLLROutputS4xD(342)(5);
  VNStageIntLLRInputS4xD(16)(5) <= CNStageIntLLROutputS4xD(343)(0);
  VNStageIntLLRInputS4xD(86)(3) <= CNStageIntLLROutputS4xD(343)(1);
  VNStageIntLLRInputS4xD(156)(3) <= CNStageIntLLROutputS4xD(343)(2);
  VNStageIntLLRInputS4xD(240)(6) <= CNStageIntLLROutputS4xD(343)(3);
  VNStageIntLLRInputS4xD(296)(5) <= CNStageIntLLROutputS4xD(343)(4);
  VNStageIntLLRInputS4xD(335)(6) <= CNStageIntLLROutputS4xD(343)(5);
  VNStageIntLLRInputS4xD(15)(6) <= CNStageIntLLROutputS4xD(344)(0);
  VNStageIntLLRInputS4xD(91)(6) <= CNStageIntLLROutputS4xD(344)(1);
  VNStageIntLLRInputS4xD(175)(6) <= CNStageIntLLROutputS4xD(344)(2);
  VNStageIntLLRInputS4xD(231)(5) <= CNStageIntLLROutputS4xD(344)(3);
  VNStageIntLLRInputS4xD(270)(6) <= CNStageIntLLROutputS4xD(344)(4);
  VNStageIntLLRInputS4xD(336)(5) <= CNStageIntLLROutputS4xD(344)(5);
  VNStageIntLLRInputS4xD(14)(6) <= CNStageIntLLROutputS4xD(345)(0);
  VNStageIntLLRInputS4xD(110)(6) <= CNStageIntLLROutputS4xD(345)(1);
  VNStageIntLLRInputS4xD(166)(5) <= CNStageIntLLROutputS4xD(345)(2);
  VNStageIntLLRInputS4xD(205)(2) <= CNStageIntLLROutputS4xD(345)(3);
  VNStageIntLLRInputS4xD(271)(5) <= CNStageIntLLROutputS4xD(345)(4);
  VNStageIntLLRInputS4xD(360)(6) <= CNStageIntLLROutputS4xD(345)(5);
  VNStageIntLLRInputS4xD(13)(5) <= CNStageIntLLROutputS4xD(346)(0);
  VNStageIntLLRInputS4xD(101)(6) <= CNStageIntLLROutputS4xD(346)(1);
  VNStageIntLLRInputS4xD(140)(6) <= CNStageIntLLROutputS4xD(346)(2);
  VNStageIntLLRInputS4xD(206)(4) <= CNStageIntLLROutputS4xD(346)(3);
  VNStageIntLLRInputS4xD(295)(4) <= CNStageIntLLROutputS4xD(346)(4);
  VNStageIntLLRInputS4xD(381)(5) <= CNStageIntLLROutputS4xD(346)(5);
  VNStageIntLLRInputS4xD(12)(6) <= CNStageIntLLROutputS4xD(347)(0);
  VNStageIntLLRInputS4xD(75)(6) <= CNStageIntLLROutputS4xD(347)(1);
  VNStageIntLLRInputS4xD(141)(4) <= CNStageIntLLROutputS4xD(347)(2);
  VNStageIntLLRInputS4xD(230)(5) <= CNStageIntLLROutputS4xD(347)(3);
  VNStageIntLLRInputS4xD(316)(4) <= CNStageIntLLROutputS4xD(347)(4);
  VNStageIntLLRInputS4xD(377)(4) <= CNStageIntLLROutputS4xD(347)(5);
  VNStageIntLLRInputS4xD(11)(5) <= CNStageIntLLROutputS4xD(348)(0);
  VNStageIntLLRInputS4xD(76)(6) <= CNStageIntLLROutputS4xD(348)(1);
  VNStageIntLLRInputS4xD(165)(5) <= CNStageIntLLROutputS4xD(348)(2);
  VNStageIntLLRInputS4xD(251)(4) <= CNStageIntLLROutputS4xD(348)(3);
  VNStageIntLLRInputS4xD(312)(5) <= CNStageIntLLROutputS4xD(348)(4);
  VNStageIntLLRInputS4xD(329)(6) <= CNStageIntLLROutputS4xD(348)(5);
  VNStageIntLLRInputS4xD(10)(4) <= CNStageIntLLROutputS4xD(349)(0);
  VNStageIntLLRInputS4xD(100)(6) <= CNStageIntLLROutputS4xD(349)(1);
  VNStageIntLLRInputS4xD(186)(5) <= CNStageIntLLROutputS4xD(349)(2);
  VNStageIntLLRInputS4xD(247)(6) <= CNStageIntLLROutputS4xD(349)(3);
  VNStageIntLLRInputS4xD(264)(6) <= CNStageIntLLROutputS4xD(349)(4);
  VNStageIntLLRInputS4xD(355)(6) <= CNStageIntLLROutputS4xD(349)(5);
  VNStageIntLLRInputS4xD(9)(6) <= CNStageIntLLROutputS4xD(350)(0);
  VNStageIntLLRInputS4xD(121)(5) <= CNStageIntLLROutputS4xD(350)(1);
  VNStageIntLLRInputS4xD(182)(6) <= CNStageIntLLROutputS4xD(350)(2);
  VNStageIntLLRInputS4xD(199)(6) <= CNStageIntLLROutputS4xD(350)(3);
  VNStageIntLLRInputS4xD(290)(5) <= CNStageIntLLROutputS4xD(350)(4);
  VNStageIntLLRInputS4xD(331)(4) <= CNStageIntLLROutputS4xD(350)(5);
  VNStageIntLLRInputS4xD(7)(6) <= CNStageIntLLROutputS4xD(351)(0);
  VNStageIntLLRInputS4xD(69)(6) <= CNStageIntLLROutputS4xD(351)(1);
  VNStageIntLLRInputS4xD(160)(6) <= CNStageIntLLROutputS4xD(351)(2);
  VNStageIntLLRInputS4xD(201)(5) <= CNStageIntLLROutputS4xD(351)(3);
  VNStageIntLLRInputS4xD(298)(6) <= CNStageIntLLROutputS4xD(351)(4);
  VNStageIntLLRInputS4xD(379)(4) <= CNStageIntLLROutputS4xD(351)(5);
  VNStageIntLLRInputS4xD(6)(6) <= CNStageIntLLROutputS4xD(352)(0);
  VNStageIntLLRInputS4xD(95)(6) <= CNStageIntLLROutputS4xD(352)(1);
  VNStageIntLLRInputS4xD(136)(6) <= CNStageIntLLROutputS4xD(352)(2);
  VNStageIntLLRInputS4xD(233)(4) <= CNStageIntLLROutputS4xD(352)(3);
  VNStageIntLLRInputS4xD(314)(3) <= CNStageIntLLROutputS4xD(352)(4);
  VNStageIntLLRInputS4xD(349)(5) <= CNStageIntLLROutputS4xD(352)(5);
  VNStageIntLLRInputS4xD(5)(6) <= CNStageIntLLROutputS4xD(353)(0);
  VNStageIntLLRInputS4xD(71)(5) <= CNStageIntLLROutputS4xD(353)(1);
  VNStageIntLLRInputS4xD(168)(5) <= CNStageIntLLROutputS4xD(353)(2);
  VNStageIntLLRInputS4xD(249)(4) <= CNStageIntLLROutputS4xD(353)(3);
  VNStageIntLLRInputS4xD(284)(6) <= CNStageIntLLROutputS4xD(353)(4);
  VNStageIntLLRInputS4xD(358)(5) <= CNStageIntLLROutputS4xD(353)(5);
  VNStageIntLLRInputS4xD(4)(5) <= CNStageIntLLROutputS4xD(354)(0);
  VNStageIntLLRInputS4xD(103)(6) <= CNStageIntLLROutputS4xD(354)(1);
  VNStageIntLLRInputS4xD(184)(6) <= CNStageIntLLROutputS4xD(354)(2);
  VNStageIntLLRInputS4xD(219)(5) <= CNStageIntLLROutputS4xD(354)(3);
  VNStageIntLLRInputS4xD(293)(5) <= CNStageIntLLROutputS4xD(354)(4);
  VNStageIntLLRInputS4xD(371)(4) <= CNStageIntLLROutputS4xD(354)(5);
  VNStageIntLLRInputS4xD(2)(6) <= CNStageIntLLROutputS4xD(355)(0);
  VNStageIntLLRInputS4xD(89)(5) <= CNStageIntLLROutputS4xD(355)(1);
  VNStageIntLLRInputS4xD(163)(4) <= CNStageIntLLROutputS4xD(355)(2);
  VNStageIntLLRInputS4xD(241)(5) <= CNStageIntLLROutputS4xD(355)(3);
  VNStageIntLLRInputS4xD(285)(6) <= CNStageIntLLROutputS4xD(355)(4);
  VNStageIntLLRInputS4xD(378)(5) <= CNStageIntLLROutputS4xD(355)(5);
  VNStageIntLLRInputS4xD(1)(5) <= CNStageIntLLROutputS4xD(356)(0);
  VNStageIntLLRInputS4xD(98)(5) <= CNStageIntLLROutputS4xD(356)(1);
  VNStageIntLLRInputS4xD(176)(6) <= CNStageIntLLROutputS4xD(356)(2);
  VNStageIntLLRInputS4xD(220)(6) <= CNStageIntLLROutputS4xD(356)(3);
  VNStageIntLLRInputS4xD(313)(3) <= CNStageIntLLROutputS4xD(356)(4);
  VNStageIntLLRInputS4xD(380)(5) <= CNStageIntLLROutputS4xD(356)(5);
  VNStageIntLLRInputS4xD(63)(3) <= CNStageIntLLROutputS4xD(357)(0);
  VNStageIntLLRInputS4xD(111)(6) <= CNStageIntLLROutputS4xD(357)(1);
  VNStageIntLLRInputS4xD(155)(6) <= CNStageIntLLROutputS4xD(357)(2);
  VNStageIntLLRInputS4xD(248)(6) <= CNStageIntLLROutputS4xD(357)(3);
  VNStageIntLLRInputS4xD(315)(5) <= CNStageIntLLROutputS4xD(357)(4);
  VNStageIntLLRInputS4xD(362)(6) <= CNStageIntLLROutputS4xD(357)(5);
  VNStageIntLLRInputS4xD(62)(5) <= CNStageIntLLROutputS4xD(358)(0);
  VNStageIntLLRInputS4xD(90)(6) <= CNStageIntLLROutputS4xD(358)(1);
  VNStageIntLLRInputS4xD(183)(4) <= CNStageIntLLROutputS4xD(358)(2);
  VNStageIntLLRInputS4xD(250)(4) <= CNStageIntLLROutputS4xD(358)(3);
  VNStageIntLLRInputS4xD(297)(6) <= CNStageIntLLROutputS4xD(358)(4);
  VNStageIntLLRInputS4xD(369)(4) <= CNStageIntLLROutputS4xD(358)(5);
  VNStageIntLLRInputS4xD(61)(5) <= CNStageIntLLROutputS4xD(359)(0);
  VNStageIntLLRInputS4xD(118)(5) <= CNStageIntLLROutputS4xD(359)(1);
  VNStageIntLLRInputS4xD(185)(3) <= CNStageIntLLROutputS4xD(359)(2);
  VNStageIntLLRInputS4xD(232)(5) <= CNStageIntLLROutputS4xD(359)(3);
  VNStageIntLLRInputS4xD(304)(6) <= CNStageIntLLROutputS4xD(359)(4);
  VNStageIntLLRInputS4xD(333)(5) <= CNStageIntLLROutputS4xD(359)(5);
  VNStageIntLLRInputS4xD(60)(5) <= CNStageIntLLROutputS4xD(360)(0);
  VNStageIntLLRInputS4xD(120)(3) <= CNStageIntLLROutputS4xD(360)(1);
  VNStageIntLLRInputS4xD(167)(6) <= CNStageIntLLROutputS4xD(360)(2);
  VNStageIntLLRInputS4xD(239)(6) <= CNStageIntLLROutputS4xD(360)(3);
  VNStageIntLLRInputS4xD(268)(6) <= CNStageIntLLROutputS4xD(360)(4);
  VNStageIntLLRInputS4xD(321)(6) <= CNStageIntLLROutputS4xD(360)(5);
  VNStageIntLLRInputS4xD(59)(4) <= CNStageIntLLROutputS4xD(361)(0);
  VNStageIntLLRInputS4xD(102)(5) <= CNStageIntLLROutputS4xD(361)(1);
  VNStageIntLLRInputS4xD(174)(4) <= CNStageIntLLROutputS4xD(361)(2);
  VNStageIntLLRInputS4xD(203)(6) <= CNStageIntLLROutputS4xD(361)(3);
  VNStageIntLLRInputS4xD(319)(6) <= CNStageIntLLROutputS4xD(361)(4);
  VNStageIntLLRInputS4xD(327)(6) <= CNStageIntLLROutputS4xD(361)(5);
  VNStageIntLLRInputS4xD(58)(4) <= CNStageIntLLROutputS4xD(362)(0);
  VNStageIntLLRInputS4xD(109)(5) <= CNStageIntLLROutputS4xD(362)(1);
  VNStageIntLLRInputS4xD(138)(6) <= CNStageIntLLROutputS4xD(362)(2);
  VNStageIntLLRInputS4xD(254)(4) <= CNStageIntLLROutputS4xD(362)(3);
  VNStageIntLLRInputS4xD(262)(5) <= CNStageIntLLROutputS4xD(362)(4);
  VNStageIntLLRInputS4xD(322)(5) <= CNStageIntLLROutputS4xD(362)(5);
  VNStageIntLLRInputS4xD(57)(5) <= CNStageIntLLROutputS4xD(363)(0);
  VNStageIntLLRInputS4xD(73)(5) <= CNStageIntLLROutputS4xD(363)(1);
  VNStageIntLLRInputS4xD(189)(5) <= CNStageIntLLROutputS4xD(363)(2);
  VNStageIntLLRInputS4xD(197)(6) <= CNStageIntLLROutputS4xD(363)(3);
  VNStageIntLLRInputS4xD(257)(6) <= CNStageIntLLROutputS4xD(363)(4);
  VNStageIntLLRInputS4xD(332)(5) <= CNStageIntLLROutputS4xD(363)(5);
  VNStageIntLLRInputS4xD(56)(6) <= CNStageIntLLROutputS4xD(364)(0);
  VNStageIntLLRInputS4xD(124)(4) <= CNStageIntLLROutputS4xD(364)(1);
  VNStageIntLLRInputS4xD(132)(5) <= CNStageIntLLROutputS4xD(364)(2);
  VNStageIntLLRInputS4xD(255)(6) <= CNStageIntLLROutputS4xD(364)(3);
  VNStageIntLLRInputS4xD(267)(6) <= CNStageIntLLROutputS4xD(364)(4);
  VNStageIntLLRInputS4xD(354)(5) <= CNStageIntLLROutputS4xD(364)(5);
  VNStageIntLLRInputS4xD(55)(6) <= CNStageIntLLROutputS4xD(365)(0);
  VNStageIntLLRInputS4xD(67)(3) <= CNStageIntLLROutputS4xD(365)(1);
  VNStageIntLLRInputS4xD(190)(4) <= CNStageIntLLROutputS4xD(365)(2);
  VNStageIntLLRInputS4xD(202)(5) <= CNStageIntLLROutputS4xD(365)(3);
  VNStageIntLLRInputS4xD(289)(6) <= CNStageIntLLROutputS4xD(365)(4);
  VNStageIntLLRInputS4xD(372)(5) <= CNStageIntLLROutputS4xD(365)(5);
  VNStageIntLLRInputS4xD(54)(5) <= CNStageIntLLROutputS4xD(366)(0);
  VNStageIntLLRInputS4xD(125)(3) <= CNStageIntLLROutputS4xD(366)(1);
  VNStageIntLLRInputS4xD(137)(6) <= CNStageIntLLROutputS4xD(366)(2);
  VNStageIntLLRInputS4xD(224)(6) <= CNStageIntLLROutputS4xD(366)(3);
  VNStageIntLLRInputS4xD(307)(6) <= CNStageIntLLROutputS4xD(366)(4);
  VNStageIntLLRInputS4xD(357)(6) <= CNStageIntLLROutputS4xD(366)(5);
  VNStageIntLLRInputS4xD(53)(5) <= CNStageIntLLROutputS4xD(367)(0);
  VNStageIntLLRInputS4xD(72)(5) <= CNStageIntLLROutputS4xD(367)(1);
  VNStageIntLLRInputS4xD(159)(4) <= CNStageIntLLROutputS4xD(367)(2);
  VNStageIntLLRInputS4xD(242)(6) <= CNStageIntLLROutputS4xD(367)(3);
  VNStageIntLLRInputS4xD(292)(6) <= CNStageIntLLROutputS4xD(367)(4);
  VNStageIntLLRInputS4xD(344)(6) <= CNStageIntLLROutputS4xD(367)(5);
  VNStageIntLLRInputS4xD(52)(4) <= CNStageIntLLROutputS4xD(368)(0);
  VNStageIntLLRInputS4xD(94)(4) <= CNStageIntLLROutputS4xD(368)(1);
  VNStageIntLLRInputS4xD(177)(6) <= CNStageIntLLROutputS4xD(368)(2);
  VNStageIntLLRInputS4xD(227)(6) <= CNStageIntLLROutputS4xD(368)(3);
  VNStageIntLLRInputS4xD(279)(5) <= CNStageIntLLROutputS4xD(368)(4);
  VNStageIntLLRInputS4xD(375)(5) <= CNStageIntLLROutputS4xD(368)(5);
  VNStageIntLLRInputS4xD(51)(5) <= CNStageIntLLROutputS4xD(369)(0);
  VNStageIntLLRInputS4xD(112)(6) <= CNStageIntLLROutputS4xD(369)(1);
  VNStageIntLLRInputS4xD(162)(6) <= CNStageIntLLROutputS4xD(369)(2);
  VNStageIntLLRInputS4xD(214)(6) <= CNStageIntLLROutputS4xD(369)(3);
  VNStageIntLLRInputS4xD(310)(5) <= CNStageIntLLROutputS4xD(369)(4);
  VNStageIntLLRInputS4xD(324)(6) <= CNStageIntLLROutputS4xD(369)(5);
  VNStageIntLLRInputS4xD(50)(6) <= CNStageIntLLROutputS4xD(370)(0);
  VNStageIntLLRInputS4xD(97)(6) <= CNStageIntLLROutputS4xD(370)(1);
  VNStageIntLLRInputS4xD(149)(6) <= CNStageIntLLROutputS4xD(370)(2);
  VNStageIntLLRInputS4xD(245)(6) <= CNStageIntLLROutputS4xD(370)(3);
  VNStageIntLLRInputS4xD(259)(4) <= CNStageIntLLROutputS4xD(370)(4);
  VNStageIntLLRInputS4xD(338)(4) <= CNStageIntLLROutputS4xD(370)(5);
  VNStageIntLLRInputS4xD(49)(6) <= CNStageIntLLROutputS4xD(371)(0);
  VNStageIntLLRInputS4xD(84)(5) <= CNStageIntLLROutputS4xD(371)(1);
  VNStageIntLLRInputS4xD(180)(4) <= CNStageIntLLROutputS4xD(371)(2);
  VNStageIntLLRInputS4xD(194)(6) <= CNStageIntLLROutputS4xD(371)(3);
  VNStageIntLLRInputS4xD(273)(5) <= CNStageIntLLROutputS4xD(371)(4);
  VNStageIntLLRInputS4xD(382)(5) <= CNStageIntLLROutputS4xD(371)(5);
  VNStageIntLLRInputS4xD(48)(3) <= CNStageIntLLROutputS4xD(372)(0);
  VNStageIntLLRInputS4xD(115)(6) <= CNStageIntLLROutputS4xD(372)(1);
  VNStageIntLLRInputS4xD(129)(6) <= CNStageIntLLROutputS4xD(372)(2);
  VNStageIntLLRInputS4xD(208)(5) <= CNStageIntLLROutputS4xD(372)(3);
  VNStageIntLLRInputS4xD(317)(3) <= CNStageIntLLROutputS4xD(372)(4);
  VNStageIntLLRInputS4xD(359)(6) <= CNStageIntLLROutputS4xD(372)(5);
  VNStageIntLLRInputS4xD(47)(3) <= CNStageIntLLROutputS4xD(373)(0);
  VNStageIntLLRInputS4xD(127)(6) <= CNStageIntLLROutputS4xD(373)(1);
  VNStageIntLLRInputS4xD(143)(6) <= CNStageIntLLROutputS4xD(373)(2);
  VNStageIntLLRInputS4xD(252)(5) <= CNStageIntLLROutputS4xD(373)(3);
  VNStageIntLLRInputS4xD(294)(6) <= CNStageIntLLROutputS4xD(373)(4);
  VNStageIntLLRInputS4xD(348)(6) <= CNStageIntLLROutputS4xD(373)(5);
  VNStageIntLLRInputS4xD(46)(6) <= CNStageIntLLROutputS4xD(374)(0);
  VNStageIntLLRInputS4xD(78)(6) <= CNStageIntLLROutputS4xD(374)(1);
  VNStageIntLLRInputS4xD(187)(5) <= CNStageIntLLROutputS4xD(374)(2);
  VNStageIntLLRInputS4xD(229)(4) <= CNStageIntLLROutputS4xD(374)(3);
  VNStageIntLLRInputS4xD(283)(6) <= CNStageIntLLROutputS4xD(374)(4);
  VNStageIntLLRInputS4xD(352)(6) <= CNStageIntLLROutputS4xD(374)(5);
  VNStageIntLLRInputS4xD(45)(6) <= CNStageIntLLROutputS4xD(375)(0);
  VNStageIntLLRInputS4xD(122)(5) <= CNStageIntLLROutputS4xD(375)(1);
  VNStageIntLLRInputS4xD(164)(5) <= CNStageIntLLROutputS4xD(375)(2);
  VNStageIntLLRInputS4xD(218)(6) <= CNStageIntLLROutputS4xD(375)(3);
  VNStageIntLLRInputS4xD(287)(6) <= CNStageIntLLROutputS4xD(375)(4);
  VNStageIntLLRInputS4xD(345)(5) <= CNStageIntLLROutputS4xD(375)(5);
  VNStageIntLLRInputS4xD(44)(6) <= CNStageIntLLROutputS4xD(376)(0);
  VNStageIntLLRInputS4xD(99)(6) <= CNStageIntLLROutputS4xD(376)(1);
  VNStageIntLLRInputS4xD(153)(6) <= CNStageIntLLROutputS4xD(376)(2);
  VNStageIntLLRInputS4xD(222)(3) <= CNStageIntLLROutputS4xD(376)(3);
  VNStageIntLLRInputS4xD(280)(6) <= CNStageIntLLROutputS4xD(376)(4);
  VNStageIntLLRInputS4xD(356)(5) <= CNStageIntLLROutputS4xD(376)(5);
  VNStageIntLLRInputS4xD(43)(5) <= CNStageIntLLROutputS4xD(377)(0);
  VNStageIntLLRInputS4xD(88)(6) <= CNStageIntLLROutputS4xD(377)(1);
  VNStageIntLLRInputS4xD(157)(5) <= CNStageIntLLROutputS4xD(377)(2);
  VNStageIntLLRInputS4xD(215)(6) <= CNStageIntLLROutputS4xD(377)(3);
  VNStageIntLLRInputS4xD(291)(5) <= CNStageIntLLROutputS4xD(377)(4);
  VNStageIntLLRInputS4xD(328)(4) <= CNStageIntLLROutputS4xD(377)(5);
  VNStageIntLLRInputS4xD(42)(6) <= CNStageIntLLROutputS4xD(378)(0);
  VNStageIntLLRInputS4xD(92)(6) <= CNStageIntLLROutputS4xD(378)(1);
  VNStageIntLLRInputS4xD(150)(5) <= CNStageIntLLROutputS4xD(378)(2);
  VNStageIntLLRInputS4xD(226)(2) <= CNStageIntLLROutputS4xD(378)(3);
  VNStageIntLLRInputS4xD(263)(6) <= CNStageIntLLROutputS4xD(378)(4);
  VNStageIntLLRInputS4xD(383)(6) <= CNStageIntLLROutputS4xD(378)(5);
  VNStageIntLLRInputS4xD(41)(6) <= CNStageIntLLROutputS4xD(379)(0);
  VNStageIntLLRInputS4xD(85)(5) <= CNStageIntLLROutputS4xD(379)(1);
  VNStageIntLLRInputS4xD(161)(6) <= CNStageIntLLROutputS4xD(379)(2);
  VNStageIntLLRInputS4xD(198)(6) <= CNStageIntLLROutputS4xD(379)(3);
  VNStageIntLLRInputS4xD(318)(3) <= CNStageIntLLROutputS4xD(379)(4);
  VNStageIntLLRInputS4xD(337)(6) <= CNStageIntLLROutputS4xD(379)(5);
  VNStageIntLLRInputS4xD(40)(4) <= CNStageIntLLROutputS4xD(380)(0);
  VNStageIntLLRInputS4xD(96)(5) <= CNStageIntLLROutputS4xD(380)(1);
  VNStageIntLLRInputS4xD(133)(4) <= CNStageIntLLROutputS4xD(380)(2);
  VNStageIntLLRInputS4xD(253)(5) <= CNStageIntLLROutputS4xD(380)(3);
  VNStageIntLLRInputS4xD(272)(6) <= CNStageIntLLROutputS4xD(380)(4);
  VNStageIntLLRInputS4xD(334)(4) <= CNStageIntLLROutputS4xD(380)(5);
  VNStageIntLLRInputS4xD(39)(6) <= CNStageIntLLROutputS4xD(381)(0);
  VNStageIntLLRInputS4xD(68)(5) <= CNStageIntLLROutputS4xD(381)(1);
  VNStageIntLLRInputS4xD(188)(4) <= CNStageIntLLROutputS4xD(381)(2);
  VNStageIntLLRInputS4xD(207)(5) <= CNStageIntLLROutputS4xD(381)(3);
  VNStageIntLLRInputS4xD(269)(5) <= CNStageIntLLROutputS4xD(381)(4);
  VNStageIntLLRInputS4xD(368)(2) <= CNStageIntLLROutputS4xD(381)(5);
  VNStageIntLLRInputS4xD(38)(6) <= CNStageIntLLROutputS4xD(382)(0);
  VNStageIntLLRInputS4xD(123)(4) <= CNStageIntLLROutputS4xD(382)(1);
  VNStageIntLLRInputS4xD(142)(4) <= CNStageIntLLROutputS4xD(382)(2);
  VNStageIntLLRInputS4xD(204)(6) <= CNStageIntLLROutputS4xD(382)(3);
  VNStageIntLLRInputS4xD(303)(6) <= CNStageIntLLROutputS4xD(382)(4);
  VNStageIntLLRInputS4xD(325)(6) <= CNStageIntLLROutputS4xD(382)(5);
  VNStageIntLLRInputS4xD(37)(6) <= CNStageIntLLROutputS4xD(383)(0);
  VNStageIntLLRInputS4xD(77)(4) <= CNStageIntLLROutputS4xD(383)(1);
  VNStageIntLLRInputS4xD(139)(6) <= CNStageIntLLROutputS4xD(383)(2);
  VNStageIntLLRInputS4xD(238)(6) <= CNStageIntLLROutputS4xD(383)(3);
  VNStageIntLLRInputS4xD(260)(5) <= CNStageIntLLROutputS4xD(383)(4);
  VNStageIntLLRInputS4xD(374)(6) <= CNStageIntLLROutputS4xD(383)(5);

  -- Check Nodes (Iteration 5)
  CNStageIntLLRInputS5xD(53)(0) <= VNStageIntLLROutputS4xD(0)(0);
  CNStageIntLLRInputS5xD(110)(0) <= VNStageIntLLROutputS4xD(0)(1);
  CNStageIntLLRInputS5xD(170)(0) <= VNStageIntLLROutputS4xD(0)(2);
  CNStageIntLLRInputS5xD(224)(0) <= VNStageIntLLROutputS4xD(0)(3);
  CNStageIntLLRInputS5xD(279)(0) <= VNStageIntLLROutputS4xD(0)(4);
  CNStageIntLLRInputS5xD(332)(0) <= VNStageIntLLROutputS4xD(0)(5);
  CNStageIntLLRInputS5xD(51)(0) <= VNStageIntLLROutputS4xD(1)(0);
  CNStageIntLLRInputS5xD(139)(0) <= VNStageIntLLROutputS4xD(1)(1);
  CNStageIntLLRInputS5xD(223)(0) <= VNStageIntLLROutputS4xD(1)(2);
  CNStageIntLLRInputS5xD(241)(0) <= VNStageIntLLROutputS4xD(1)(3);
  CNStageIntLLRInputS5xD(307)(0) <= VNStageIntLLROutputS4xD(1)(4);
  CNStageIntLLRInputS5xD(356)(0) <= VNStageIntLLROutputS4xD(1)(5);
  CNStageIntLLRInputS5xD(50)(0) <= VNStageIntLLROutputS4xD(2)(0);
  CNStageIntLLRInputS5xD(92)(0) <= VNStageIntLLROutputS4xD(2)(1);
  CNStageIntLLRInputS5xD(138)(0) <= VNStageIntLLROutputS4xD(2)(2);
  CNStageIntLLRInputS5xD(222)(0) <= VNStageIntLLROutputS4xD(2)(3);
  CNStageIntLLRInputS5xD(240)(0) <= VNStageIntLLROutputS4xD(2)(4);
  CNStageIntLLRInputS5xD(306)(0) <= VNStageIntLLROutputS4xD(2)(5);
  CNStageIntLLRInputS5xD(355)(0) <= VNStageIntLLROutputS4xD(2)(6);
  CNStageIntLLRInputS5xD(91)(0) <= VNStageIntLLROutputS4xD(3)(0);
  CNStageIntLLRInputS5xD(137)(0) <= VNStageIntLLROutputS4xD(3)(1);
  CNStageIntLLRInputS5xD(221)(0) <= VNStageIntLLROutputS4xD(3)(2);
  CNStageIntLLRInputS5xD(239)(0) <= VNStageIntLLROutputS4xD(3)(3);
  CNStageIntLLRInputS5xD(305)(0) <= VNStageIntLLROutputS4xD(3)(4);
  CNStageIntLLRInputS5xD(49)(0) <= VNStageIntLLROutputS4xD(4)(0);
  CNStageIntLLRInputS5xD(90)(0) <= VNStageIntLLROutputS4xD(4)(1);
  CNStageIntLLRInputS5xD(220)(0) <= VNStageIntLLROutputS4xD(4)(2);
  CNStageIntLLRInputS5xD(238)(0) <= VNStageIntLLROutputS4xD(4)(3);
  CNStageIntLLRInputS5xD(304)(0) <= VNStageIntLLROutputS4xD(4)(4);
  CNStageIntLLRInputS5xD(354)(0) <= VNStageIntLLROutputS4xD(4)(5);
  CNStageIntLLRInputS5xD(48)(0) <= VNStageIntLLROutputS4xD(5)(0);
  CNStageIntLLRInputS5xD(89)(0) <= VNStageIntLLROutputS4xD(5)(1);
  CNStageIntLLRInputS5xD(136)(0) <= VNStageIntLLROutputS4xD(5)(2);
  CNStageIntLLRInputS5xD(219)(0) <= VNStageIntLLROutputS4xD(5)(3);
  CNStageIntLLRInputS5xD(237)(0) <= VNStageIntLLROutputS4xD(5)(4);
  CNStageIntLLRInputS5xD(303)(0) <= VNStageIntLLROutputS4xD(5)(5);
  CNStageIntLLRInputS5xD(353)(0) <= VNStageIntLLROutputS4xD(5)(6);
  CNStageIntLLRInputS5xD(47)(0) <= VNStageIntLLROutputS4xD(6)(0);
  CNStageIntLLRInputS5xD(88)(0) <= VNStageIntLLROutputS4xD(6)(1);
  CNStageIntLLRInputS5xD(135)(0) <= VNStageIntLLROutputS4xD(6)(2);
  CNStageIntLLRInputS5xD(218)(0) <= VNStageIntLLROutputS4xD(6)(3);
  CNStageIntLLRInputS5xD(236)(0) <= VNStageIntLLROutputS4xD(6)(4);
  CNStageIntLLRInputS5xD(302)(0) <= VNStageIntLLROutputS4xD(6)(5);
  CNStageIntLLRInputS5xD(352)(0) <= VNStageIntLLROutputS4xD(6)(6);
  CNStageIntLLRInputS5xD(46)(0) <= VNStageIntLLROutputS4xD(7)(0);
  CNStageIntLLRInputS5xD(87)(0) <= VNStageIntLLROutputS4xD(7)(1);
  CNStageIntLLRInputS5xD(134)(0) <= VNStageIntLLROutputS4xD(7)(2);
  CNStageIntLLRInputS5xD(217)(0) <= VNStageIntLLROutputS4xD(7)(3);
  CNStageIntLLRInputS5xD(235)(0) <= VNStageIntLLROutputS4xD(7)(4);
  CNStageIntLLRInputS5xD(301)(0) <= VNStageIntLLROutputS4xD(7)(5);
  CNStageIntLLRInputS5xD(351)(0) <= VNStageIntLLROutputS4xD(7)(6);
  CNStageIntLLRInputS5xD(45)(0) <= VNStageIntLLROutputS4xD(8)(0);
  CNStageIntLLRInputS5xD(133)(0) <= VNStageIntLLROutputS4xD(8)(1);
  CNStageIntLLRInputS5xD(216)(0) <= VNStageIntLLROutputS4xD(8)(2);
  CNStageIntLLRInputS5xD(44)(0) <= VNStageIntLLROutputS4xD(9)(0);
  CNStageIntLLRInputS5xD(86)(0) <= VNStageIntLLROutputS4xD(9)(1);
  CNStageIntLLRInputS5xD(132)(0) <= VNStageIntLLROutputS4xD(9)(2);
  CNStageIntLLRInputS5xD(215)(0) <= VNStageIntLLROutputS4xD(9)(3);
  CNStageIntLLRInputS5xD(234)(0) <= VNStageIntLLROutputS4xD(9)(4);
  CNStageIntLLRInputS5xD(300)(0) <= VNStageIntLLROutputS4xD(9)(5);
  CNStageIntLLRInputS5xD(350)(0) <= VNStageIntLLROutputS4xD(9)(6);
  CNStageIntLLRInputS5xD(43)(0) <= VNStageIntLLROutputS4xD(10)(0);
  CNStageIntLLRInputS5xD(85)(0) <= VNStageIntLLROutputS4xD(10)(1);
  CNStageIntLLRInputS5xD(131)(0) <= VNStageIntLLROutputS4xD(10)(2);
  CNStageIntLLRInputS5xD(233)(0) <= VNStageIntLLROutputS4xD(10)(3);
  CNStageIntLLRInputS5xD(349)(0) <= VNStageIntLLROutputS4xD(10)(4);
  CNStageIntLLRInputS5xD(42)(0) <= VNStageIntLLROutputS4xD(11)(0);
  CNStageIntLLRInputS5xD(84)(0) <= VNStageIntLLROutputS4xD(11)(1);
  CNStageIntLLRInputS5xD(130)(0) <= VNStageIntLLROutputS4xD(11)(2);
  CNStageIntLLRInputS5xD(214)(0) <= VNStageIntLLROutputS4xD(11)(3);
  CNStageIntLLRInputS5xD(232)(0) <= VNStageIntLLROutputS4xD(11)(4);
  CNStageIntLLRInputS5xD(348)(0) <= VNStageIntLLROutputS4xD(11)(5);
  CNStageIntLLRInputS5xD(41)(0) <= VNStageIntLLROutputS4xD(12)(0);
  CNStageIntLLRInputS5xD(83)(0) <= VNStageIntLLROutputS4xD(12)(1);
  CNStageIntLLRInputS5xD(129)(0) <= VNStageIntLLROutputS4xD(12)(2);
  CNStageIntLLRInputS5xD(213)(0) <= VNStageIntLLROutputS4xD(12)(3);
  CNStageIntLLRInputS5xD(231)(0) <= VNStageIntLLROutputS4xD(12)(4);
  CNStageIntLLRInputS5xD(299)(0) <= VNStageIntLLROutputS4xD(12)(5);
  CNStageIntLLRInputS5xD(347)(0) <= VNStageIntLLROutputS4xD(12)(6);
  CNStageIntLLRInputS5xD(82)(0) <= VNStageIntLLROutputS4xD(13)(0);
  CNStageIntLLRInputS5xD(128)(0) <= VNStageIntLLROutputS4xD(13)(1);
  CNStageIntLLRInputS5xD(212)(0) <= VNStageIntLLROutputS4xD(13)(2);
  CNStageIntLLRInputS5xD(230)(0) <= VNStageIntLLROutputS4xD(13)(3);
  CNStageIntLLRInputS5xD(298)(0) <= VNStageIntLLROutputS4xD(13)(4);
  CNStageIntLLRInputS5xD(346)(0) <= VNStageIntLLROutputS4xD(13)(5);
  CNStageIntLLRInputS5xD(40)(0) <= VNStageIntLLROutputS4xD(14)(0);
  CNStageIntLLRInputS5xD(81)(0) <= VNStageIntLLROutputS4xD(14)(1);
  CNStageIntLLRInputS5xD(127)(0) <= VNStageIntLLROutputS4xD(14)(2);
  CNStageIntLLRInputS5xD(211)(0) <= VNStageIntLLROutputS4xD(14)(3);
  CNStageIntLLRInputS5xD(229)(0) <= VNStageIntLLROutputS4xD(14)(4);
  CNStageIntLLRInputS5xD(297)(0) <= VNStageIntLLROutputS4xD(14)(5);
  CNStageIntLLRInputS5xD(345)(0) <= VNStageIntLLROutputS4xD(14)(6);
  CNStageIntLLRInputS5xD(39)(0) <= VNStageIntLLROutputS4xD(15)(0);
  CNStageIntLLRInputS5xD(80)(0) <= VNStageIntLLROutputS4xD(15)(1);
  CNStageIntLLRInputS5xD(126)(0) <= VNStageIntLLROutputS4xD(15)(2);
  CNStageIntLLRInputS5xD(210)(0) <= VNStageIntLLROutputS4xD(15)(3);
  CNStageIntLLRInputS5xD(228)(0) <= VNStageIntLLROutputS4xD(15)(4);
  CNStageIntLLRInputS5xD(296)(0) <= VNStageIntLLROutputS4xD(15)(5);
  CNStageIntLLRInputS5xD(344)(0) <= VNStageIntLLROutputS4xD(15)(6);
  CNStageIntLLRInputS5xD(38)(0) <= VNStageIntLLROutputS4xD(16)(0);
  CNStageIntLLRInputS5xD(125)(0) <= VNStageIntLLROutputS4xD(16)(1);
  CNStageIntLLRInputS5xD(209)(0) <= VNStageIntLLROutputS4xD(16)(2);
  CNStageIntLLRInputS5xD(227)(0) <= VNStageIntLLROutputS4xD(16)(3);
  CNStageIntLLRInputS5xD(295)(0) <= VNStageIntLLROutputS4xD(16)(4);
  CNStageIntLLRInputS5xD(343)(0) <= VNStageIntLLROutputS4xD(16)(5);
  CNStageIntLLRInputS5xD(37)(0) <= VNStageIntLLROutputS4xD(17)(0);
  CNStageIntLLRInputS5xD(79)(0) <= VNStageIntLLROutputS4xD(17)(1);
  CNStageIntLLRInputS5xD(124)(0) <= VNStageIntLLROutputS4xD(17)(2);
  CNStageIntLLRInputS5xD(208)(0) <= VNStageIntLLROutputS4xD(17)(3);
  CNStageIntLLRInputS5xD(226)(0) <= VNStageIntLLROutputS4xD(17)(4);
  CNStageIntLLRInputS5xD(294)(0) <= VNStageIntLLROutputS4xD(17)(5);
  CNStageIntLLRInputS5xD(342)(0) <= VNStageIntLLROutputS4xD(17)(6);
  CNStageIntLLRInputS5xD(36)(0) <= VNStageIntLLROutputS4xD(18)(0);
  CNStageIntLLRInputS5xD(78)(0) <= VNStageIntLLROutputS4xD(18)(1);
  CNStageIntLLRInputS5xD(123)(0) <= VNStageIntLLROutputS4xD(18)(2);
  CNStageIntLLRInputS5xD(207)(0) <= VNStageIntLLROutputS4xD(18)(3);
  CNStageIntLLRInputS5xD(225)(0) <= VNStageIntLLROutputS4xD(18)(4);
  CNStageIntLLRInputS5xD(293)(0) <= VNStageIntLLROutputS4xD(18)(5);
  CNStageIntLLRInputS5xD(341)(0) <= VNStageIntLLROutputS4xD(18)(6);
  CNStageIntLLRInputS5xD(35)(0) <= VNStageIntLLROutputS4xD(19)(0);
  CNStageIntLLRInputS5xD(77)(0) <= VNStageIntLLROutputS4xD(19)(1);
  CNStageIntLLRInputS5xD(122)(0) <= VNStageIntLLROutputS4xD(19)(2);
  CNStageIntLLRInputS5xD(278)(0) <= VNStageIntLLROutputS4xD(19)(3);
  CNStageIntLLRInputS5xD(340)(0) <= VNStageIntLLROutputS4xD(19)(4);
  CNStageIntLLRInputS5xD(34)(0) <= VNStageIntLLROutputS4xD(20)(0);
  CNStageIntLLRInputS5xD(76)(0) <= VNStageIntLLROutputS4xD(20)(1);
  CNStageIntLLRInputS5xD(277)(0) <= VNStageIntLLROutputS4xD(20)(2);
  CNStageIntLLRInputS5xD(292)(0) <= VNStageIntLLROutputS4xD(20)(3);
  CNStageIntLLRInputS5xD(339)(0) <= VNStageIntLLROutputS4xD(20)(4);
  CNStageIntLLRInputS5xD(33)(0) <= VNStageIntLLROutputS4xD(21)(0);
  CNStageIntLLRInputS5xD(75)(0) <= VNStageIntLLROutputS4xD(21)(1);
  CNStageIntLLRInputS5xD(121)(0) <= VNStageIntLLROutputS4xD(21)(2);
  CNStageIntLLRInputS5xD(206)(0) <= VNStageIntLLROutputS4xD(21)(3);
  CNStageIntLLRInputS5xD(276)(0) <= VNStageIntLLROutputS4xD(21)(4);
  CNStageIntLLRInputS5xD(291)(0) <= VNStageIntLLROutputS4xD(21)(5);
  CNStageIntLLRInputS5xD(338)(0) <= VNStageIntLLROutputS4xD(21)(6);
  CNStageIntLLRInputS5xD(32)(0) <= VNStageIntLLROutputS4xD(22)(0);
  CNStageIntLLRInputS5xD(74)(0) <= VNStageIntLLROutputS4xD(22)(1);
  CNStageIntLLRInputS5xD(120)(0) <= VNStageIntLLROutputS4xD(22)(2);
  CNStageIntLLRInputS5xD(205)(0) <= VNStageIntLLROutputS4xD(22)(3);
  CNStageIntLLRInputS5xD(275)(0) <= VNStageIntLLROutputS4xD(22)(4);
  CNStageIntLLRInputS5xD(290)(0) <= VNStageIntLLROutputS4xD(22)(5);
  CNStageIntLLRInputS5xD(337)(0) <= VNStageIntLLROutputS4xD(22)(6);
  CNStageIntLLRInputS5xD(31)(0) <= VNStageIntLLROutputS4xD(23)(0);
  CNStageIntLLRInputS5xD(73)(0) <= VNStageIntLLROutputS4xD(23)(1);
  CNStageIntLLRInputS5xD(119)(0) <= VNStageIntLLROutputS4xD(23)(2);
  CNStageIntLLRInputS5xD(204)(0) <= VNStageIntLLROutputS4xD(23)(3);
  CNStageIntLLRInputS5xD(274)(0) <= VNStageIntLLROutputS4xD(23)(4);
  CNStageIntLLRInputS5xD(289)(0) <= VNStageIntLLROutputS4xD(23)(5);
  CNStageIntLLRInputS5xD(336)(0) <= VNStageIntLLROutputS4xD(23)(6);
  CNStageIntLLRInputS5xD(30)(0) <= VNStageIntLLROutputS4xD(24)(0);
  CNStageIntLLRInputS5xD(72)(0) <= VNStageIntLLROutputS4xD(24)(1);
  CNStageIntLLRInputS5xD(118)(0) <= VNStageIntLLROutputS4xD(24)(2);
  CNStageIntLLRInputS5xD(203)(0) <= VNStageIntLLROutputS4xD(24)(3);
  CNStageIntLLRInputS5xD(273)(0) <= VNStageIntLLROutputS4xD(24)(4);
  CNStageIntLLRInputS5xD(288)(0) <= VNStageIntLLROutputS4xD(24)(5);
  CNStageIntLLRInputS5xD(335)(0) <= VNStageIntLLROutputS4xD(24)(6);
  CNStageIntLLRInputS5xD(29)(0) <= VNStageIntLLROutputS4xD(25)(0);
  CNStageIntLLRInputS5xD(71)(0) <= VNStageIntLLROutputS4xD(25)(1);
  CNStageIntLLRInputS5xD(117)(0) <= VNStageIntLLROutputS4xD(25)(2);
  CNStageIntLLRInputS5xD(202)(0) <= VNStageIntLLROutputS4xD(25)(3);
  CNStageIntLLRInputS5xD(287)(0) <= VNStageIntLLROutputS4xD(25)(4);
  CNStageIntLLRInputS5xD(28)(0) <= VNStageIntLLROutputS4xD(26)(0);
  CNStageIntLLRInputS5xD(70)(0) <= VNStageIntLLROutputS4xD(26)(1);
  CNStageIntLLRInputS5xD(116)(0) <= VNStageIntLLROutputS4xD(26)(2);
  CNStageIntLLRInputS5xD(201)(0) <= VNStageIntLLROutputS4xD(26)(3);
  CNStageIntLLRInputS5xD(272)(0) <= VNStageIntLLROutputS4xD(26)(4);
  CNStageIntLLRInputS5xD(286)(0) <= VNStageIntLLROutputS4xD(26)(5);
  CNStageIntLLRInputS5xD(334)(0) <= VNStageIntLLROutputS4xD(26)(6);
  CNStageIntLLRInputS5xD(27)(0) <= VNStageIntLLROutputS4xD(27)(0);
  CNStageIntLLRInputS5xD(69)(0) <= VNStageIntLLROutputS4xD(27)(1);
  CNStageIntLLRInputS5xD(115)(0) <= VNStageIntLLROutputS4xD(27)(2);
  CNStageIntLLRInputS5xD(200)(0) <= VNStageIntLLROutputS4xD(27)(3);
  CNStageIntLLRInputS5xD(285)(0) <= VNStageIntLLROutputS4xD(27)(4);
  CNStageIntLLRInputS5xD(26)(0) <= VNStageIntLLROutputS4xD(28)(0);
  CNStageIntLLRInputS5xD(68)(0) <= VNStageIntLLROutputS4xD(28)(1);
  CNStageIntLLRInputS5xD(114)(0) <= VNStageIntLLROutputS4xD(28)(2);
  CNStageIntLLRInputS5xD(199)(0) <= VNStageIntLLROutputS4xD(28)(3);
  CNStageIntLLRInputS5xD(271)(0) <= VNStageIntLLROutputS4xD(28)(4);
  CNStageIntLLRInputS5xD(333)(0) <= VNStageIntLLROutputS4xD(28)(5);
  CNStageIntLLRInputS5xD(25)(0) <= VNStageIntLLROutputS4xD(29)(0);
  CNStageIntLLRInputS5xD(67)(0) <= VNStageIntLLROutputS4xD(29)(1);
  CNStageIntLLRInputS5xD(113)(0) <= VNStageIntLLROutputS4xD(29)(2);
  CNStageIntLLRInputS5xD(270)(0) <= VNStageIntLLROutputS4xD(29)(3);
  CNStageIntLLRInputS5xD(24)(0) <= VNStageIntLLROutputS4xD(30)(0);
  CNStageIntLLRInputS5xD(66)(0) <= VNStageIntLLROutputS4xD(30)(1);
  CNStageIntLLRInputS5xD(112)(0) <= VNStageIntLLROutputS4xD(30)(2);
  CNStageIntLLRInputS5xD(198)(0) <= VNStageIntLLROutputS4xD(30)(3);
  CNStageIntLLRInputS5xD(269)(0) <= VNStageIntLLROutputS4xD(30)(4);
  CNStageIntLLRInputS5xD(284)(0) <= VNStageIntLLROutputS4xD(30)(5);
  CNStageIntLLRInputS5xD(23)(0) <= VNStageIntLLROutputS4xD(31)(0);
  CNStageIntLLRInputS5xD(65)(0) <= VNStageIntLLROutputS4xD(31)(1);
  CNStageIntLLRInputS5xD(197)(0) <= VNStageIntLLROutputS4xD(31)(2);
  CNStageIntLLRInputS5xD(283)(0) <= VNStageIntLLROutputS4xD(31)(3);
  CNStageIntLLRInputS5xD(22)(0) <= VNStageIntLLROutputS4xD(32)(0);
  CNStageIntLLRInputS5xD(64)(0) <= VNStageIntLLROutputS4xD(32)(1);
  CNStageIntLLRInputS5xD(111)(0) <= VNStageIntLLROutputS4xD(32)(2);
  CNStageIntLLRInputS5xD(268)(0) <= VNStageIntLLROutputS4xD(32)(3);
  CNStageIntLLRInputS5xD(21)(0) <= VNStageIntLLROutputS4xD(33)(0);
  CNStageIntLLRInputS5xD(63)(0) <= VNStageIntLLROutputS4xD(33)(1);
  CNStageIntLLRInputS5xD(169)(0) <= VNStageIntLLROutputS4xD(33)(2);
  CNStageIntLLRInputS5xD(196)(0) <= VNStageIntLLROutputS4xD(33)(3);
  CNStageIntLLRInputS5xD(267)(0) <= VNStageIntLLROutputS4xD(33)(4);
  CNStageIntLLRInputS5xD(282)(0) <= VNStageIntLLROutputS4xD(33)(5);
  CNStageIntLLRInputS5xD(20)(0) <= VNStageIntLLROutputS4xD(34)(0);
  CNStageIntLLRInputS5xD(62)(0) <= VNStageIntLLROutputS4xD(34)(1);
  CNStageIntLLRInputS5xD(168)(0) <= VNStageIntLLROutputS4xD(34)(2);
  CNStageIntLLRInputS5xD(195)(0) <= VNStageIntLLROutputS4xD(34)(3);
  CNStageIntLLRInputS5xD(266)(0) <= VNStageIntLLROutputS4xD(34)(4);
  CNStageIntLLRInputS5xD(281)(0) <= VNStageIntLLROutputS4xD(34)(5);
  CNStageIntLLRInputS5xD(19)(0) <= VNStageIntLLROutputS4xD(35)(0);
  CNStageIntLLRInputS5xD(61)(0) <= VNStageIntLLROutputS4xD(35)(1);
  CNStageIntLLRInputS5xD(167)(0) <= VNStageIntLLROutputS4xD(35)(2);
  CNStageIntLLRInputS5xD(194)(0) <= VNStageIntLLROutputS4xD(35)(3);
  CNStageIntLLRInputS5xD(265)(0) <= VNStageIntLLROutputS4xD(35)(4);
  CNStageIntLLRInputS5xD(280)(0) <= VNStageIntLLROutputS4xD(35)(5);
  CNStageIntLLRInputS5xD(18)(0) <= VNStageIntLLROutputS4xD(36)(0);
  CNStageIntLLRInputS5xD(60)(0) <= VNStageIntLLROutputS4xD(36)(1);
  CNStageIntLLRInputS5xD(166)(0) <= VNStageIntLLROutputS4xD(36)(2);
  CNStageIntLLRInputS5xD(264)(0) <= VNStageIntLLROutputS4xD(36)(3);
  CNStageIntLLRInputS5xD(17)(0) <= VNStageIntLLROutputS4xD(37)(0);
  CNStageIntLLRInputS5xD(59)(0) <= VNStageIntLLROutputS4xD(37)(1);
  CNStageIntLLRInputS5xD(165)(0) <= VNStageIntLLROutputS4xD(37)(2);
  CNStageIntLLRInputS5xD(193)(0) <= VNStageIntLLROutputS4xD(37)(3);
  CNStageIntLLRInputS5xD(263)(0) <= VNStageIntLLROutputS4xD(37)(4);
  CNStageIntLLRInputS5xD(331)(0) <= VNStageIntLLROutputS4xD(37)(5);
  CNStageIntLLRInputS5xD(383)(0) <= VNStageIntLLROutputS4xD(37)(6);
  CNStageIntLLRInputS5xD(16)(0) <= VNStageIntLLROutputS4xD(38)(0);
  CNStageIntLLRInputS5xD(58)(0) <= VNStageIntLLROutputS4xD(38)(1);
  CNStageIntLLRInputS5xD(164)(0) <= VNStageIntLLROutputS4xD(38)(2);
  CNStageIntLLRInputS5xD(192)(0) <= VNStageIntLLROutputS4xD(38)(3);
  CNStageIntLLRInputS5xD(262)(0) <= VNStageIntLLROutputS4xD(38)(4);
  CNStageIntLLRInputS5xD(330)(0) <= VNStageIntLLROutputS4xD(38)(5);
  CNStageIntLLRInputS5xD(382)(0) <= VNStageIntLLROutputS4xD(38)(6);
  CNStageIntLLRInputS5xD(15)(0) <= VNStageIntLLROutputS4xD(39)(0);
  CNStageIntLLRInputS5xD(57)(0) <= VNStageIntLLROutputS4xD(39)(1);
  CNStageIntLLRInputS5xD(163)(0) <= VNStageIntLLROutputS4xD(39)(2);
  CNStageIntLLRInputS5xD(191)(0) <= VNStageIntLLROutputS4xD(39)(3);
  CNStageIntLLRInputS5xD(261)(0) <= VNStageIntLLROutputS4xD(39)(4);
  CNStageIntLLRInputS5xD(329)(0) <= VNStageIntLLROutputS4xD(39)(5);
  CNStageIntLLRInputS5xD(381)(0) <= VNStageIntLLROutputS4xD(39)(6);
  CNStageIntLLRInputS5xD(14)(0) <= VNStageIntLLROutputS4xD(40)(0);
  CNStageIntLLRInputS5xD(56)(0) <= VNStageIntLLROutputS4xD(40)(1);
  CNStageIntLLRInputS5xD(162)(0) <= VNStageIntLLROutputS4xD(40)(2);
  CNStageIntLLRInputS5xD(260)(0) <= VNStageIntLLROutputS4xD(40)(3);
  CNStageIntLLRInputS5xD(380)(0) <= VNStageIntLLROutputS4xD(40)(4);
  CNStageIntLLRInputS5xD(13)(0) <= VNStageIntLLROutputS4xD(41)(0);
  CNStageIntLLRInputS5xD(55)(0) <= VNStageIntLLROutputS4xD(41)(1);
  CNStageIntLLRInputS5xD(161)(0) <= VNStageIntLLROutputS4xD(41)(2);
  CNStageIntLLRInputS5xD(190)(0) <= VNStageIntLLROutputS4xD(41)(3);
  CNStageIntLLRInputS5xD(259)(0) <= VNStageIntLLROutputS4xD(41)(4);
  CNStageIntLLRInputS5xD(328)(0) <= VNStageIntLLROutputS4xD(41)(5);
  CNStageIntLLRInputS5xD(379)(0) <= VNStageIntLLROutputS4xD(41)(6);
  CNStageIntLLRInputS5xD(12)(0) <= VNStageIntLLROutputS4xD(42)(0);
  CNStageIntLLRInputS5xD(54)(0) <= VNStageIntLLROutputS4xD(42)(1);
  CNStageIntLLRInputS5xD(160)(0) <= VNStageIntLLROutputS4xD(42)(2);
  CNStageIntLLRInputS5xD(189)(0) <= VNStageIntLLROutputS4xD(42)(3);
  CNStageIntLLRInputS5xD(258)(0) <= VNStageIntLLROutputS4xD(42)(4);
  CNStageIntLLRInputS5xD(327)(0) <= VNStageIntLLROutputS4xD(42)(5);
  CNStageIntLLRInputS5xD(378)(0) <= VNStageIntLLROutputS4xD(42)(6);
  CNStageIntLLRInputS5xD(109)(0) <= VNStageIntLLROutputS4xD(43)(0);
  CNStageIntLLRInputS5xD(159)(0) <= VNStageIntLLROutputS4xD(43)(1);
  CNStageIntLLRInputS5xD(188)(0) <= VNStageIntLLROutputS4xD(43)(2);
  CNStageIntLLRInputS5xD(257)(0) <= VNStageIntLLROutputS4xD(43)(3);
  CNStageIntLLRInputS5xD(326)(0) <= VNStageIntLLROutputS4xD(43)(4);
  CNStageIntLLRInputS5xD(377)(0) <= VNStageIntLLROutputS4xD(43)(5);
  CNStageIntLLRInputS5xD(11)(0) <= VNStageIntLLROutputS4xD(44)(0);
  CNStageIntLLRInputS5xD(108)(0) <= VNStageIntLLROutputS4xD(44)(1);
  CNStageIntLLRInputS5xD(158)(0) <= VNStageIntLLROutputS4xD(44)(2);
  CNStageIntLLRInputS5xD(187)(0) <= VNStageIntLLROutputS4xD(44)(3);
  CNStageIntLLRInputS5xD(256)(0) <= VNStageIntLLROutputS4xD(44)(4);
  CNStageIntLLRInputS5xD(325)(0) <= VNStageIntLLROutputS4xD(44)(5);
  CNStageIntLLRInputS5xD(376)(0) <= VNStageIntLLROutputS4xD(44)(6);
  CNStageIntLLRInputS5xD(10)(0) <= VNStageIntLLROutputS4xD(45)(0);
  CNStageIntLLRInputS5xD(107)(0) <= VNStageIntLLROutputS4xD(45)(1);
  CNStageIntLLRInputS5xD(157)(0) <= VNStageIntLLROutputS4xD(45)(2);
  CNStageIntLLRInputS5xD(186)(0) <= VNStageIntLLROutputS4xD(45)(3);
  CNStageIntLLRInputS5xD(255)(0) <= VNStageIntLLROutputS4xD(45)(4);
  CNStageIntLLRInputS5xD(324)(0) <= VNStageIntLLROutputS4xD(45)(5);
  CNStageIntLLRInputS5xD(375)(0) <= VNStageIntLLROutputS4xD(45)(6);
  CNStageIntLLRInputS5xD(9)(0) <= VNStageIntLLROutputS4xD(46)(0);
  CNStageIntLLRInputS5xD(106)(0) <= VNStageIntLLROutputS4xD(46)(1);
  CNStageIntLLRInputS5xD(156)(0) <= VNStageIntLLROutputS4xD(46)(2);
  CNStageIntLLRInputS5xD(185)(0) <= VNStageIntLLROutputS4xD(46)(3);
  CNStageIntLLRInputS5xD(254)(0) <= VNStageIntLLROutputS4xD(46)(4);
  CNStageIntLLRInputS5xD(323)(0) <= VNStageIntLLROutputS4xD(46)(5);
  CNStageIntLLRInputS5xD(374)(0) <= VNStageIntLLROutputS4xD(46)(6);
  CNStageIntLLRInputS5xD(8)(0) <= VNStageIntLLROutputS4xD(47)(0);
  CNStageIntLLRInputS5xD(155)(0) <= VNStageIntLLROutputS4xD(47)(1);
  CNStageIntLLRInputS5xD(253)(0) <= VNStageIntLLROutputS4xD(47)(2);
  CNStageIntLLRInputS5xD(373)(0) <= VNStageIntLLROutputS4xD(47)(3);
  CNStageIntLLRInputS5xD(7)(0) <= VNStageIntLLROutputS4xD(48)(0);
  CNStageIntLLRInputS5xD(154)(0) <= VNStageIntLLROutputS4xD(48)(1);
  CNStageIntLLRInputS5xD(322)(0) <= VNStageIntLLROutputS4xD(48)(2);
  CNStageIntLLRInputS5xD(372)(0) <= VNStageIntLLROutputS4xD(48)(3);
  CNStageIntLLRInputS5xD(6)(0) <= VNStageIntLLROutputS4xD(49)(0);
  CNStageIntLLRInputS5xD(105)(0) <= VNStageIntLLROutputS4xD(49)(1);
  CNStageIntLLRInputS5xD(153)(0) <= VNStageIntLLROutputS4xD(49)(2);
  CNStageIntLLRInputS5xD(184)(0) <= VNStageIntLLROutputS4xD(49)(3);
  CNStageIntLLRInputS5xD(252)(0) <= VNStageIntLLROutputS4xD(49)(4);
  CNStageIntLLRInputS5xD(321)(0) <= VNStageIntLLROutputS4xD(49)(5);
  CNStageIntLLRInputS5xD(371)(0) <= VNStageIntLLROutputS4xD(49)(6);
  CNStageIntLLRInputS5xD(5)(0) <= VNStageIntLLROutputS4xD(50)(0);
  CNStageIntLLRInputS5xD(104)(0) <= VNStageIntLLROutputS4xD(50)(1);
  CNStageIntLLRInputS5xD(152)(0) <= VNStageIntLLROutputS4xD(50)(2);
  CNStageIntLLRInputS5xD(183)(0) <= VNStageIntLLROutputS4xD(50)(3);
  CNStageIntLLRInputS5xD(251)(0) <= VNStageIntLLROutputS4xD(50)(4);
  CNStageIntLLRInputS5xD(320)(0) <= VNStageIntLLROutputS4xD(50)(5);
  CNStageIntLLRInputS5xD(370)(0) <= VNStageIntLLROutputS4xD(50)(6);
  CNStageIntLLRInputS5xD(4)(0) <= VNStageIntLLROutputS4xD(51)(0);
  CNStageIntLLRInputS5xD(103)(0) <= VNStageIntLLROutputS4xD(51)(1);
  CNStageIntLLRInputS5xD(182)(0) <= VNStageIntLLROutputS4xD(51)(2);
  CNStageIntLLRInputS5xD(250)(0) <= VNStageIntLLROutputS4xD(51)(3);
  CNStageIntLLRInputS5xD(319)(0) <= VNStageIntLLROutputS4xD(51)(4);
  CNStageIntLLRInputS5xD(369)(0) <= VNStageIntLLROutputS4xD(51)(5);
  CNStageIntLLRInputS5xD(102)(0) <= VNStageIntLLROutputS4xD(52)(0);
  CNStageIntLLRInputS5xD(151)(0) <= VNStageIntLLROutputS4xD(52)(1);
  CNStageIntLLRInputS5xD(181)(0) <= VNStageIntLLROutputS4xD(52)(2);
  CNStageIntLLRInputS5xD(318)(0) <= VNStageIntLLROutputS4xD(52)(3);
  CNStageIntLLRInputS5xD(368)(0) <= VNStageIntLLROutputS4xD(52)(4);
  CNStageIntLLRInputS5xD(3)(0) <= VNStageIntLLROutputS4xD(53)(0);
  CNStageIntLLRInputS5xD(150)(0) <= VNStageIntLLROutputS4xD(53)(1);
  CNStageIntLLRInputS5xD(180)(0) <= VNStageIntLLROutputS4xD(53)(2);
  CNStageIntLLRInputS5xD(249)(0) <= VNStageIntLLROutputS4xD(53)(3);
  CNStageIntLLRInputS5xD(317)(0) <= VNStageIntLLROutputS4xD(53)(4);
  CNStageIntLLRInputS5xD(367)(0) <= VNStageIntLLROutputS4xD(53)(5);
  CNStageIntLLRInputS5xD(2)(0) <= VNStageIntLLROutputS4xD(54)(0);
  CNStageIntLLRInputS5xD(101)(0) <= VNStageIntLLROutputS4xD(54)(1);
  CNStageIntLLRInputS5xD(149)(0) <= VNStageIntLLROutputS4xD(54)(2);
  CNStageIntLLRInputS5xD(179)(0) <= VNStageIntLLROutputS4xD(54)(3);
  CNStageIntLLRInputS5xD(316)(0) <= VNStageIntLLROutputS4xD(54)(4);
  CNStageIntLLRInputS5xD(366)(0) <= VNStageIntLLROutputS4xD(54)(5);
  CNStageIntLLRInputS5xD(1)(0) <= VNStageIntLLROutputS4xD(55)(0);
  CNStageIntLLRInputS5xD(100)(0) <= VNStageIntLLROutputS4xD(55)(1);
  CNStageIntLLRInputS5xD(148)(0) <= VNStageIntLLROutputS4xD(55)(2);
  CNStageIntLLRInputS5xD(178)(0) <= VNStageIntLLROutputS4xD(55)(3);
  CNStageIntLLRInputS5xD(248)(0) <= VNStageIntLLROutputS4xD(55)(4);
  CNStageIntLLRInputS5xD(315)(0) <= VNStageIntLLROutputS4xD(55)(5);
  CNStageIntLLRInputS5xD(365)(0) <= VNStageIntLLROutputS4xD(55)(6);
  CNStageIntLLRInputS5xD(0)(0) <= VNStageIntLLROutputS4xD(56)(0);
  CNStageIntLLRInputS5xD(99)(0) <= VNStageIntLLROutputS4xD(56)(1);
  CNStageIntLLRInputS5xD(147)(0) <= VNStageIntLLROutputS4xD(56)(2);
  CNStageIntLLRInputS5xD(177)(0) <= VNStageIntLLROutputS4xD(56)(3);
  CNStageIntLLRInputS5xD(247)(0) <= VNStageIntLLROutputS4xD(56)(4);
  CNStageIntLLRInputS5xD(314)(0) <= VNStageIntLLROutputS4xD(56)(5);
  CNStageIntLLRInputS5xD(364)(0) <= VNStageIntLLROutputS4xD(56)(6);
  CNStageIntLLRInputS5xD(98)(0) <= VNStageIntLLROutputS4xD(57)(0);
  CNStageIntLLRInputS5xD(146)(0) <= VNStageIntLLROutputS4xD(57)(1);
  CNStageIntLLRInputS5xD(176)(0) <= VNStageIntLLROutputS4xD(57)(2);
  CNStageIntLLRInputS5xD(246)(0) <= VNStageIntLLROutputS4xD(57)(3);
  CNStageIntLLRInputS5xD(313)(0) <= VNStageIntLLROutputS4xD(57)(4);
  CNStageIntLLRInputS5xD(363)(0) <= VNStageIntLLROutputS4xD(57)(5);
  CNStageIntLLRInputS5xD(97)(0) <= VNStageIntLLROutputS4xD(58)(0);
  CNStageIntLLRInputS5xD(145)(0) <= VNStageIntLLROutputS4xD(58)(1);
  CNStageIntLLRInputS5xD(175)(0) <= VNStageIntLLROutputS4xD(58)(2);
  CNStageIntLLRInputS5xD(312)(0) <= VNStageIntLLROutputS4xD(58)(3);
  CNStageIntLLRInputS5xD(362)(0) <= VNStageIntLLROutputS4xD(58)(4);
  CNStageIntLLRInputS5xD(144)(0) <= VNStageIntLLROutputS4xD(59)(0);
  CNStageIntLLRInputS5xD(174)(0) <= VNStageIntLLROutputS4xD(59)(1);
  CNStageIntLLRInputS5xD(245)(0) <= VNStageIntLLROutputS4xD(59)(2);
  CNStageIntLLRInputS5xD(311)(0) <= VNStageIntLLROutputS4xD(59)(3);
  CNStageIntLLRInputS5xD(361)(0) <= VNStageIntLLROutputS4xD(59)(4);
  CNStageIntLLRInputS5xD(96)(0) <= VNStageIntLLROutputS4xD(60)(0);
  CNStageIntLLRInputS5xD(143)(0) <= VNStageIntLLROutputS4xD(60)(1);
  CNStageIntLLRInputS5xD(173)(0) <= VNStageIntLLROutputS4xD(60)(2);
  CNStageIntLLRInputS5xD(244)(0) <= VNStageIntLLROutputS4xD(60)(3);
  CNStageIntLLRInputS5xD(310)(0) <= VNStageIntLLROutputS4xD(60)(4);
  CNStageIntLLRInputS5xD(360)(0) <= VNStageIntLLROutputS4xD(60)(5);
  CNStageIntLLRInputS5xD(95)(0) <= VNStageIntLLROutputS4xD(61)(0);
  CNStageIntLLRInputS5xD(142)(0) <= VNStageIntLLROutputS4xD(61)(1);
  CNStageIntLLRInputS5xD(172)(0) <= VNStageIntLLROutputS4xD(61)(2);
  CNStageIntLLRInputS5xD(243)(0) <= VNStageIntLLROutputS4xD(61)(3);
  CNStageIntLLRInputS5xD(309)(0) <= VNStageIntLLROutputS4xD(61)(4);
  CNStageIntLLRInputS5xD(359)(0) <= VNStageIntLLROutputS4xD(61)(5);
  CNStageIntLLRInputS5xD(94)(0) <= VNStageIntLLROutputS4xD(62)(0);
  CNStageIntLLRInputS5xD(141)(0) <= VNStageIntLLROutputS4xD(62)(1);
  CNStageIntLLRInputS5xD(171)(0) <= VNStageIntLLROutputS4xD(62)(2);
  CNStageIntLLRInputS5xD(242)(0) <= VNStageIntLLROutputS4xD(62)(3);
  CNStageIntLLRInputS5xD(308)(0) <= VNStageIntLLROutputS4xD(62)(4);
  CNStageIntLLRInputS5xD(358)(0) <= VNStageIntLLROutputS4xD(62)(5);
  CNStageIntLLRInputS5xD(52)(0) <= VNStageIntLLROutputS4xD(63)(0);
  CNStageIntLLRInputS5xD(93)(0) <= VNStageIntLLROutputS4xD(63)(1);
  CNStageIntLLRInputS5xD(140)(0) <= VNStageIntLLROutputS4xD(63)(2);
  CNStageIntLLRInputS5xD(357)(0) <= VNStageIntLLROutputS4xD(63)(3);
  CNStageIntLLRInputS5xD(53)(1) <= VNStageIntLLROutputS4xD(64)(0);
  CNStageIntLLRInputS5xD(109)(1) <= VNStageIntLLROutputS4xD(64)(1);
  CNStageIntLLRInputS5xD(130)(1) <= VNStageIntLLROutputS4xD(64)(2);
  CNStageIntLLRInputS5xD(245)(1) <= VNStageIntLLROutputS4xD(64)(3);
  CNStageIntLLRInputS5xD(299)(1) <= VNStageIntLLROutputS4xD(64)(4);
  CNStageIntLLRInputS5xD(342)(1) <= VNStageIntLLROutputS4xD(64)(5);
  CNStageIntLLRInputS5xD(51)(1) <= VNStageIntLLROutputS4xD(65)(0);
  CNStageIntLLRInputS5xD(74)(1) <= VNStageIntLLROutputS4xD(65)(1);
  CNStageIntLLRInputS5xD(141)(1) <= VNStageIntLLROutputS4xD(65)(2);
  CNStageIntLLRInputS5xD(189)(1) <= VNStageIntLLROutputS4xD(65)(3);
  CNStageIntLLRInputS5xD(286)(1) <= VNStageIntLLROutputS4xD(65)(4);
  CNStageIntLLRInputS5xD(50)(1) <= VNStageIntLLROutputS4xD(66)(0);
  CNStageIntLLRInputS5xD(66)(1) <= VNStageIntLLROutputS4xD(66)(1);
  CNStageIntLLRInputS5xD(155)(1) <= VNStageIntLLROutputS4xD(66)(2);
  CNStageIntLLRInputS5xD(244)(1) <= VNStageIntLLROutputS4xD(66)(3);
  CNStageIntLLRInputS5xD(97)(1) <= VNStageIntLLROutputS4xD(67)(0);
  CNStageIntLLRInputS5xD(275)(1) <= VNStageIntLLROutputS4xD(67)(1);
  CNStageIntLLRInputS5xD(322)(1) <= VNStageIntLLROutputS4xD(67)(2);
  CNStageIntLLRInputS5xD(365)(1) <= VNStageIntLLROutputS4xD(67)(3);
  CNStageIntLLRInputS5xD(49)(1) <= VNStageIntLLROutputS4xD(68)(0);
  CNStageIntLLRInputS5xD(112)(1) <= VNStageIntLLROutputS4xD(68)(1);
  CNStageIntLLRInputS5xD(210)(1) <= VNStageIntLLROutputS4xD(68)(2);
  CNStageIntLLRInputS5xD(256)(1) <= VNStageIntLLROutputS4xD(68)(3);
  CNStageIntLLRInputS5xD(318)(1) <= VNStageIntLLROutputS4xD(68)(4);
  CNStageIntLLRInputS5xD(381)(1) <= VNStageIntLLROutputS4xD(68)(5);
  CNStageIntLLRInputS5xD(48)(1) <= VNStageIntLLROutputS4xD(69)(0);
  CNStageIntLLRInputS5xD(101)(1) <= VNStageIntLLROutputS4xD(69)(1);
  CNStageIntLLRInputS5xD(135)(1) <= VNStageIntLLROutputS4xD(69)(2);
  CNStageIntLLRInputS5xD(215)(1) <= VNStageIntLLROutputS4xD(69)(3);
  CNStageIntLLRInputS5xD(259)(1) <= VNStageIntLLROutputS4xD(69)(4);
  CNStageIntLLRInputS5xD(283)(1) <= VNStageIntLLROutputS4xD(69)(5);
  CNStageIntLLRInputS5xD(351)(1) <= VNStageIntLLROutputS4xD(69)(6);
  CNStageIntLLRInputS5xD(47)(1) <= VNStageIntLLROutputS4xD(70)(0);
  CNStageIntLLRInputS5xD(104)(1) <= VNStageIntLLROutputS4xD(70)(1);
  CNStageIntLLRInputS5xD(136)(1) <= VNStageIntLLROutputS4xD(70)(2);
  CNStageIntLLRInputS5xD(206)(1) <= VNStageIntLLROutputS4xD(70)(3);
  CNStageIntLLRInputS5xD(246)(1) <= VNStageIntLLROutputS4xD(70)(4);
  CNStageIntLLRInputS5xD(301)(1) <= VNStageIntLLROutputS4xD(70)(5);
  CNStageIntLLRInputS5xD(46)(1) <= VNStageIntLLROutputS4xD(71)(0);
  CNStageIntLLRInputS5xD(95)(1) <= VNStageIntLLROutputS4xD(71)(1);
  CNStageIntLLRInputS5xD(176)(1) <= VNStageIntLLROutputS4xD(71)(2);
  CNStageIntLLRInputS5xD(276)(1) <= VNStageIntLLROutputS4xD(71)(3);
  CNStageIntLLRInputS5xD(302)(1) <= VNStageIntLLROutputS4xD(71)(4);
  CNStageIntLLRInputS5xD(353)(1) <= VNStageIntLLROutputS4xD(71)(5);
  CNStageIntLLRInputS5xD(45)(1) <= VNStageIntLLROutputS4xD(72)(0);
  CNStageIntLLRInputS5xD(75)(1) <= VNStageIntLLROutputS4xD(72)(1);
  CNStageIntLLRInputS5xD(162)(1) <= VNStageIntLLROutputS4xD(72)(2);
  CNStageIntLLRInputS5xD(183)(1) <= VNStageIntLLROutputS4xD(72)(3);
  CNStageIntLLRInputS5xD(243)(1) <= VNStageIntLLROutputS4xD(72)(4);
  CNStageIntLLRInputS5xD(367)(1) <= VNStageIntLLROutputS4xD(72)(5);
  CNStageIntLLRInputS5xD(44)(1) <= VNStageIntLLROutputS4xD(73)(0);
  CNStageIntLLRInputS5xD(56)(1) <= VNStageIntLLROutputS4xD(73)(1);
  CNStageIntLLRInputS5xD(121)(1) <= VNStageIntLLROutputS4xD(73)(2);
  CNStageIntLLRInputS5xD(219)(1) <= VNStageIntLLROutputS4xD(73)(3);
  CNStageIntLLRInputS5xD(328)(1) <= VNStageIntLLROutputS4xD(73)(4);
  CNStageIntLLRInputS5xD(363)(1) <= VNStageIntLLROutputS4xD(73)(5);
  CNStageIntLLRInputS5xD(43)(1) <= VNStageIntLLROutputS4xD(74)(0);
  CNStageIntLLRInputS5xD(70)(1) <= VNStageIntLLROutputS4xD(74)(1);
  CNStageIntLLRInputS5xD(125)(1) <= VNStageIntLLROutputS4xD(74)(2);
  CNStageIntLLRInputS5xD(221)(1) <= VNStageIntLLROutputS4xD(74)(3);
  CNStageIntLLRInputS5xD(290)(1) <= VNStageIntLLROutputS4xD(74)(4);
  CNStageIntLLRInputS5xD(42)(1) <= VNStageIntLLROutputS4xD(75)(0);
  CNStageIntLLRInputS5xD(81)(1) <= VNStageIntLLROutputS4xD(75)(1);
  CNStageIntLLRInputS5xD(170)(1) <= VNStageIntLLROutputS4xD(75)(2);
  CNStageIntLLRInputS5xD(192)(1) <= VNStageIntLLROutputS4xD(75)(3);
  CNStageIntLLRInputS5xD(278)(1) <= VNStageIntLLROutputS4xD(75)(4);
  CNStageIntLLRInputS5xD(294)(1) <= VNStageIntLLROutputS4xD(75)(5);
  CNStageIntLLRInputS5xD(347)(1) <= VNStageIntLLROutputS4xD(75)(6);
  CNStageIntLLRInputS5xD(41)(1) <= VNStageIntLLROutputS4xD(76)(0);
  CNStageIntLLRInputS5xD(106)(1) <= VNStageIntLLROutputS4xD(76)(1);
  CNStageIntLLRInputS5xD(124)(1) <= VNStageIntLLROutputS4xD(76)(2);
  CNStageIntLLRInputS5xD(174)(1) <= VNStageIntLLROutputS4xD(76)(3);
  CNStageIntLLRInputS5xD(270)(1) <= VNStageIntLLROutputS4xD(76)(4);
  CNStageIntLLRInputS5xD(332)(1) <= VNStageIntLLROutputS4xD(76)(5);
  CNStageIntLLRInputS5xD(348)(1) <= VNStageIntLLROutputS4xD(76)(6);
  CNStageIntLLRInputS5xD(119)(1) <= VNStageIntLLROutputS4xD(77)(0);
  CNStageIntLLRInputS5xD(185)(1) <= VNStageIntLLROutputS4xD(77)(1);
  CNStageIntLLRInputS5xD(257)(1) <= VNStageIntLLROutputS4xD(77)(2);
  CNStageIntLLRInputS5xD(293)(1) <= VNStageIntLLROutputS4xD(77)(3);
  CNStageIntLLRInputS5xD(383)(1) <= VNStageIntLLROutputS4xD(77)(4);
  CNStageIntLLRInputS5xD(40)(1) <= VNStageIntLLROutputS4xD(78)(0);
  CNStageIntLLRInputS5xD(84)(1) <= VNStageIntLLROutputS4xD(78)(1);
  CNStageIntLLRInputS5xD(159)(1) <= VNStageIntLLROutputS4xD(78)(2);
  CNStageIntLLRInputS5xD(193)(1) <= VNStageIntLLROutputS4xD(78)(3);
  CNStageIntLLRInputS5xD(274)(1) <= VNStageIntLLROutputS4xD(78)(4);
  CNStageIntLLRInputS5xD(288)(1) <= VNStageIntLLROutputS4xD(78)(5);
  CNStageIntLLRInputS5xD(374)(1) <= VNStageIntLLROutputS4xD(78)(6);
  CNStageIntLLRInputS5xD(39)(1) <= VNStageIntLLROutputS4xD(79)(0);
  CNStageIntLLRInputS5xD(99)(1) <= VNStageIntLLROutputS4xD(79)(1);
  CNStageIntLLRInputS5xD(167)(1) <= VNStageIntLLROutputS4xD(79)(2);
  CNStageIntLLRInputS5xD(220)(1) <= VNStageIntLLROutputS4xD(79)(3);
  CNStageIntLLRInputS5xD(325)(1) <= VNStageIntLLROutputS4xD(79)(4);
  CNStageIntLLRInputS5xD(38)(1) <= VNStageIntLLROutputS4xD(80)(0);
  CNStageIntLLRInputS5xD(62)(1) <= VNStageIntLLROutputS4xD(80)(1);
  CNStageIntLLRInputS5xD(131)(1) <= VNStageIntLLROutputS4xD(80)(2);
  CNStageIntLLRInputS5xD(182)(1) <= VNStageIntLLROutputS4xD(80)(3);
  CNStageIntLLRInputS5xD(248)(1) <= VNStageIntLLROutputS4xD(80)(4);
  CNStageIntLLRInputS5xD(337)(1) <= VNStageIntLLROutputS4xD(80)(5);
  CNStageIntLLRInputS5xD(37)(1) <= VNStageIntLLROutputS4xD(81)(0);
  CNStageIntLLRInputS5xD(72)(1) <= VNStageIntLLROutputS4xD(81)(1);
  CNStageIntLLRInputS5xD(129)(1) <= VNStageIntLLROutputS4xD(81)(2);
  CNStageIntLLRInputS5xD(262)(1) <= VNStageIntLLROutputS4xD(81)(3);
  CNStageIntLLRInputS5xD(36)(1) <= VNStageIntLLROutputS4xD(82)(0);
  CNStageIntLLRInputS5xD(67)(1) <= VNStageIntLLROutputS4xD(82)(1);
  CNStageIntLLRInputS5xD(165)(1) <= VNStageIntLLROutputS4xD(82)(2);
  CNStageIntLLRInputS5xD(188)(1) <= VNStageIntLLROutputS4xD(82)(3);
  CNStageIntLLRInputS5xD(254)(1) <= VNStageIntLLROutputS4xD(82)(4);
  CNStageIntLLRInputS5xD(298)(1) <= VNStageIntLLROutputS4xD(82)(5);
  CNStageIntLLRInputS5xD(336)(1) <= VNStageIntLLROutputS4xD(82)(6);
  CNStageIntLLRInputS5xD(35)(1) <= VNStageIntLLROutputS4xD(83)(0);
  CNStageIntLLRInputS5xD(73)(1) <= VNStageIntLLROutputS4xD(83)(1);
  CNStageIntLLRInputS5xD(144)(1) <= VNStageIntLLROutputS4xD(83)(2);
  CNStageIntLLRInputS5xD(208)(1) <= VNStageIntLLROutputS4xD(83)(3);
  CNStageIntLLRInputS5xD(232)(1) <= VNStageIntLLROutputS4xD(83)(4);
  CNStageIntLLRInputS5xD(330)(1) <= VNStageIntLLROutputS4xD(83)(5);
  CNStageIntLLRInputS5xD(34)(1) <= VNStageIntLLROutputS4xD(84)(0);
  CNStageIntLLRInputS5xD(61)(1) <= VNStageIntLLROutputS4xD(84)(1);
  CNStageIntLLRInputS5xD(147)(1) <= VNStageIntLLROutputS4xD(84)(2);
  CNStageIntLLRInputS5xD(222)(1) <= VNStageIntLLROutputS4xD(84)(3);
  CNStageIntLLRInputS5xD(310)(1) <= VNStageIntLLROutputS4xD(84)(4);
  CNStageIntLLRInputS5xD(371)(1) <= VNStageIntLLROutputS4xD(84)(5);
  CNStageIntLLRInputS5xD(33)(1) <= VNStageIntLLROutputS4xD(85)(0);
  CNStageIntLLRInputS5xD(132)(1) <= VNStageIntLLROutputS4xD(85)(1);
  CNStageIntLLRInputS5xD(218)(1) <= VNStageIntLLROutputS4xD(85)(2);
  CNStageIntLLRInputS5xD(235)(1) <= VNStageIntLLROutputS4xD(85)(3);
  CNStageIntLLRInputS5xD(313)(1) <= VNStageIntLLROutputS4xD(85)(4);
  CNStageIntLLRInputS5xD(379)(1) <= VNStageIntLLROutputS4xD(85)(5);
  CNStageIntLLRInputS5xD(32)(1) <= VNStageIntLLROutputS4xD(86)(0);
  CNStageIntLLRInputS5xD(166)(1) <= VNStageIntLLROutputS4xD(86)(1);
  CNStageIntLLRInputS5xD(239)(1) <= VNStageIntLLROutputS4xD(86)(2);
  CNStageIntLLRInputS5xD(343)(1) <= VNStageIntLLROutputS4xD(86)(3);
  CNStageIntLLRInputS5xD(31)(1) <= VNStageIntLLROutputS4xD(87)(0);
  CNStageIntLLRInputS5xD(77)(1) <= VNStageIntLLROutputS4xD(87)(1);
  CNStageIntLLRInputS5xD(128)(1) <= VNStageIntLLROutputS4xD(87)(2);
  CNStageIntLLRInputS5xD(203)(1) <= VNStageIntLLROutputS4xD(87)(3);
  CNStageIntLLRInputS5xD(229)(1) <= VNStageIntLLROutputS4xD(87)(4);
  CNStageIntLLRInputS5xD(331)(1) <= VNStageIntLLROutputS4xD(87)(5);
  CNStageIntLLRInputS5xD(341)(1) <= VNStageIntLLROutputS4xD(87)(6);
  CNStageIntLLRInputS5xD(30)(1) <= VNStageIntLLROutputS4xD(88)(0);
  CNStageIntLLRInputS5xD(79)(1) <= VNStageIntLLROutputS4xD(88)(1);
  CNStageIntLLRInputS5xD(156)(1) <= VNStageIntLLROutputS4xD(88)(2);
  CNStageIntLLRInputS5xD(204)(1) <= VNStageIntLLROutputS4xD(88)(3);
  CNStageIntLLRInputS5xD(263)(1) <= VNStageIntLLROutputS4xD(88)(4);
  CNStageIntLLRInputS5xD(297)(1) <= VNStageIntLLROutputS4xD(88)(5);
  CNStageIntLLRInputS5xD(377)(1) <= VNStageIntLLROutputS4xD(88)(6);
  CNStageIntLLRInputS5xD(29)(1) <= VNStageIntLLROutputS4xD(89)(0);
  CNStageIntLLRInputS5xD(102)(1) <= VNStageIntLLROutputS4xD(89)(1);
  CNStageIntLLRInputS5xD(140)(1) <= VNStageIntLLROutputS4xD(89)(2);
  CNStageIntLLRInputS5xD(184)(1) <= VNStageIntLLROutputS4xD(89)(3);
  CNStageIntLLRInputS5xD(247)(1) <= VNStageIntLLROutputS4xD(89)(4);
  CNStageIntLLRInputS5xD(355)(1) <= VNStageIntLLROutputS4xD(89)(5);
  CNStageIntLLRInputS5xD(28)(1) <= VNStageIntLLROutputS4xD(90)(0);
  CNStageIntLLRInputS5xD(85)(1) <= VNStageIntLLROutputS4xD(90)(1);
  CNStageIntLLRInputS5xD(168)(1) <= VNStageIntLLROutputS4xD(90)(2);
  CNStageIntLLRInputS5xD(175)(1) <= VNStageIntLLROutputS4xD(90)(3);
  CNStageIntLLRInputS5xD(258)(1) <= VNStageIntLLROutputS4xD(90)(4);
  CNStageIntLLRInputS5xD(307)(1) <= VNStageIntLLROutputS4xD(90)(5);
  CNStageIntLLRInputS5xD(358)(1) <= VNStageIntLLROutputS4xD(90)(6);
  CNStageIntLLRInputS5xD(27)(1) <= VNStageIntLLROutputS4xD(91)(0);
  CNStageIntLLRInputS5xD(96)(1) <= VNStageIntLLROutputS4xD(91)(1);
  CNStageIntLLRInputS5xD(158)(1) <= VNStageIntLLROutputS4xD(91)(2);
  CNStageIntLLRInputS5xD(191)(1) <= VNStageIntLLROutputS4xD(91)(3);
  CNStageIntLLRInputS5xD(269)(1) <= VNStageIntLLROutputS4xD(91)(4);
  CNStageIntLLRInputS5xD(280)(1) <= VNStageIntLLROutputS4xD(91)(5);
  CNStageIntLLRInputS5xD(344)(1) <= VNStageIntLLROutputS4xD(91)(6);
  CNStageIntLLRInputS5xD(26)(1) <= VNStageIntLLROutputS4xD(92)(0);
  CNStageIntLLRInputS5xD(103)(1) <= VNStageIntLLROutputS4xD(92)(1);
  CNStageIntLLRInputS5xD(145)(1) <= VNStageIntLLROutputS4xD(92)(2);
  CNStageIntLLRInputS5xD(195)(1) <= VNStageIntLLROutputS4xD(92)(3);
  CNStageIntLLRInputS5xD(242)(1) <= VNStageIntLLROutputS4xD(92)(4);
  CNStageIntLLRInputS5xD(324)(1) <= VNStageIntLLROutputS4xD(92)(5);
  CNStageIntLLRInputS5xD(378)(1) <= VNStageIntLLROutputS4xD(92)(6);
  CNStageIntLLRInputS5xD(25)(1) <= VNStageIntLLROutputS4xD(93)(0);
  CNStageIntLLRInputS5xD(78)(1) <= VNStageIntLLROutputS4xD(93)(1);
  CNStageIntLLRInputS5xD(164)(1) <= VNStageIntLLROutputS4xD(93)(2);
  CNStageIntLLRInputS5xD(224)(1) <= VNStageIntLLROutputS4xD(93)(3);
  CNStageIntLLRInputS5xD(231)(1) <= VNStageIntLLROutputS4xD(93)(4);
  CNStageIntLLRInputS5xD(311)(1) <= VNStageIntLLROutputS4xD(93)(5);
  CNStageIntLLRInputS5xD(340)(1) <= VNStageIntLLROutputS4xD(93)(6);
  CNStageIntLLRInputS5xD(24)(1) <= VNStageIntLLROutputS4xD(94)(0);
  CNStageIntLLRInputS5xD(92)(1) <= VNStageIntLLROutputS4xD(94)(1);
  CNStageIntLLRInputS5xD(194)(1) <= VNStageIntLLROutputS4xD(94)(2);
  CNStageIntLLRInputS5xD(329)(1) <= VNStageIntLLROutputS4xD(94)(3);
  CNStageIntLLRInputS5xD(368)(1) <= VNStageIntLLROutputS4xD(94)(4);
  CNStageIntLLRInputS5xD(23)(1) <= VNStageIntLLROutputS4xD(95)(0);
  CNStageIntLLRInputS5xD(63)(1) <= VNStageIntLLROutputS4xD(95)(1);
  CNStageIntLLRInputS5xD(134)(1) <= VNStageIntLLROutputS4xD(95)(2);
  CNStageIntLLRInputS5xD(190)(1) <= VNStageIntLLROutputS4xD(95)(3);
  CNStageIntLLRInputS5xD(234)(1) <= VNStageIntLLROutputS4xD(95)(4);
  CNStageIntLLRInputS5xD(303)(1) <= VNStageIntLLROutputS4xD(95)(5);
  CNStageIntLLRInputS5xD(352)(1) <= VNStageIntLLROutputS4xD(95)(6);
  CNStageIntLLRInputS5xD(22)(1) <= VNStageIntLLROutputS4xD(96)(0);
  CNStageIntLLRInputS5xD(98)(1) <= VNStageIntLLROutputS4xD(96)(1);
  CNStageIntLLRInputS5xD(150)(1) <= VNStageIntLLROutputS4xD(96)(2);
  CNStageIntLLRInputS5xD(172)(1) <= VNStageIntLLROutputS4xD(96)(3);
  CNStageIntLLRInputS5xD(251)(1) <= VNStageIntLLROutputS4xD(96)(4);
  CNStageIntLLRInputS5xD(380)(1) <= VNStageIntLLROutputS4xD(96)(5);
  CNStageIntLLRInputS5xD(21)(1) <= VNStageIntLLROutputS4xD(97)(0);
  CNStageIntLLRInputS5xD(65)(1) <= VNStageIntLLROutputS4xD(97)(1);
  CNStageIntLLRInputS5xD(142)(1) <= VNStageIntLLROutputS4xD(97)(2);
  CNStageIntLLRInputS5xD(180)(1) <= VNStageIntLLROutputS4xD(97)(3);
  CNStageIntLLRInputS5xD(260)(1) <= VNStageIntLLROutputS4xD(97)(4);
  CNStageIntLLRInputS5xD(316)(1) <= VNStageIntLLROutputS4xD(97)(5);
  CNStageIntLLRInputS5xD(370)(1) <= VNStageIntLLROutputS4xD(97)(6);
  CNStageIntLLRInputS5xD(20)(1) <= VNStageIntLLROutputS4xD(98)(0);
  CNStageIntLLRInputS5xD(116)(1) <= VNStageIntLLROutputS4xD(98)(1);
  CNStageIntLLRInputS5xD(199)(1) <= VNStageIntLLROutputS4xD(98)(2);
  CNStageIntLLRInputS5xD(255)(1) <= VNStageIntLLROutputS4xD(98)(3);
  CNStageIntLLRInputS5xD(308)(1) <= VNStageIntLLROutputS4xD(98)(4);
  CNStageIntLLRInputS5xD(356)(1) <= VNStageIntLLROutputS4xD(98)(5);
  CNStageIntLLRInputS5xD(19)(1) <= VNStageIntLLROutputS4xD(99)(0);
  CNStageIntLLRInputS5xD(76)(1) <= VNStageIntLLROutputS4xD(99)(1);
  CNStageIntLLRInputS5xD(126)(1) <= VNStageIntLLROutputS4xD(99)(2);
  CNStageIntLLRInputS5xD(198)(1) <= VNStageIntLLROutputS4xD(99)(3);
  CNStageIntLLRInputS5xD(261)(1) <= VNStageIntLLROutputS4xD(99)(4);
  CNStageIntLLRInputS5xD(285)(1) <= VNStageIntLLROutputS4xD(99)(5);
  CNStageIntLLRInputS5xD(376)(1) <= VNStageIntLLROutputS4xD(99)(6);
  CNStageIntLLRInputS5xD(18)(1) <= VNStageIntLLROutputS4xD(100)(0);
  CNStageIntLLRInputS5xD(94)(1) <= VNStageIntLLROutputS4xD(100)(1);
  CNStageIntLLRInputS5xD(120)(1) <= VNStageIntLLROutputS4xD(100)(2);
  CNStageIntLLRInputS5xD(178)(1) <= VNStageIntLLROutputS4xD(100)(3);
  CNStageIntLLRInputS5xD(250)(1) <= VNStageIntLLROutputS4xD(100)(4);
  CNStageIntLLRInputS5xD(295)(1) <= VNStageIntLLROutputS4xD(100)(5);
  CNStageIntLLRInputS5xD(349)(1) <= VNStageIntLLROutputS4xD(100)(6);
  CNStageIntLLRInputS5xD(17)(1) <= VNStageIntLLROutputS4xD(101)(0);
  CNStageIntLLRInputS5xD(58)(1) <= VNStageIntLLROutputS4xD(101)(1);
  CNStageIntLLRInputS5xD(123)(1) <= VNStageIntLLROutputS4xD(101)(2);
  CNStageIntLLRInputS5xD(211)(1) <= VNStageIntLLROutputS4xD(101)(3);
  CNStageIntLLRInputS5xD(273)(1) <= VNStageIntLLROutputS4xD(101)(4);
  CNStageIntLLRInputS5xD(289)(1) <= VNStageIntLLROutputS4xD(101)(5);
  CNStageIntLLRInputS5xD(346)(1) <= VNStageIntLLROutputS4xD(101)(6);
  CNStageIntLLRInputS5xD(16)(1) <= VNStageIntLLROutputS4xD(102)(0);
  CNStageIntLLRInputS5xD(59)(1) <= VNStageIntLLROutputS4xD(102)(1);
  CNStageIntLLRInputS5xD(113)(1) <= VNStageIntLLROutputS4xD(102)(2);
  CNStageIntLLRInputS5xD(214)(1) <= VNStageIntLLROutputS4xD(102)(3);
  CNStageIntLLRInputS5xD(226)(1) <= VNStageIntLLROutputS4xD(102)(4);
  CNStageIntLLRInputS5xD(361)(1) <= VNStageIntLLROutputS4xD(102)(5);
  CNStageIntLLRInputS5xD(15)(1) <= VNStageIntLLROutputS4xD(103)(0);
  CNStageIntLLRInputS5xD(93)(1) <= VNStageIntLLROutputS4xD(103)(1);
  CNStageIntLLRInputS5xD(151)(1) <= VNStageIntLLROutputS4xD(103)(2);
  CNStageIntLLRInputS5xD(200)(1) <= VNStageIntLLROutputS4xD(103)(3);
  CNStageIntLLRInputS5xD(265)(1) <= VNStageIntLLROutputS4xD(103)(4);
  CNStageIntLLRInputS5xD(284)(1) <= VNStageIntLLROutputS4xD(103)(5);
  CNStageIntLLRInputS5xD(354)(1) <= VNStageIntLLROutputS4xD(103)(6);
  CNStageIntLLRInputS5xD(14)(1) <= VNStageIntLLROutputS4xD(104)(0);
  CNStageIntLLRInputS5xD(86)(1) <= VNStageIntLLROutputS4xD(104)(1);
  CNStageIntLLRInputS5xD(133)(1) <= VNStageIntLLROutputS4xD(104)(2);
  CNStageIntLLRInputS5xD(179)(1) <= VNStageIntLLROutputS4xD(104)(3);
  CNStageIntLLRInputS5xD(267)(1) <= VNStageIntLLROutputS4xD(104)(4);
  CNStageIntLLRInputS5xD(317)(1) <= VNStageIntLLROutputS4xD(104)(5);
  CNStageIntLLRInputS5xD(13)(1) <= VNStageIntLLROutputS4xD(105)(0);
  CNStageIntLLRInputS5xD(146)(1) <= VNStageIntLLROutputS4xD(105)(1);
  CNStageIntLLRInputS5xD(197)(1) <= VNStageIntLLROutputS4xD(105)(2);
  CNStageIntLLRInputS5xD(237)(1) <= VNStageIntLLROutputS4xD(105)(3);
  CNStageIntLLRInputS5xD(300)(1) <= VNStageIntLLROutputS4xD(105)(4);
  CNStageIntLLRInputS5xD(338)(1) <= VNStageIntLLROutputS4xD(105)(5);
  CNStageIntLLRInputS5xD(12)(1) <= VNStageIntLLROutputS4xD(106)(0);
  CNStageIntLLRInputS5xD(157)(1) <= VNStageIntLLROutputS4xD(106)(1);
  CNStageIntLLRInputS5xD(223)(1) <= VNStageIntLLROutputS4xD(106)(2);
  CNStageIntLLRInputS5xD(272)(1) <= VNStageIntLLROutputS4xD(106)(3);
  CNStageIntLLRInputS5xD(312)(1) <= VNStageIntLLROutputS4xD(106)(4);
  CNStageIntLLRInputS5xD(333)(1) <= VNStageIntLLROutputS4xD(106)(5);
  CNStageIntLLRInputS5xD(110)(1) <= VNStageIntLLROutputS4xD(107)(0);
  CNStageIntLLRInputS5xD(127)(1) <= VNStageIntLLROutputS4xD(107)(1);
  CNStageIntLLRInputS5xD(207)(1) <= VNStageIntLLROutputS4xD(107)(2);
  CNStageIntLLRInputS5xD(230)(1) <= VNStageIntLLROutputS4xD(107)(3);
  CNStageIntLLRInputS5xD(323)(1) <= VNStageIntLLROutputS4xD(107)(4);
  CNStageIntLLRInputS5xD(335)(1) <= VNStageIntLLROutputS4xD(107)(5);
  CNStageIntLLRInputS5xD(11)(1) <= VNStageIntLLROutputS4xD(108)(0);
  CNStageIntLLRInputS5xD(105)(1) <= VNStageIntLLROutputS4xD(108)(1);
  CNStageIntLLRInputS5xD(115)(1) <= VNStageIntLLROutputS4xD(108)(2);
  CNStageIntLLRInputS5xD(181)(1) <= VNStageIntLLROutputS4xD(108)(3);
  CNStageIntLLRInputS5xD(238)(1) <= VNStageIntLLROutputS4xD(108)(4);
  CNStageIntLLRInputS5xD(296)(1) <= VNStageIntLLROutputS4xD(108)(5);
  CNStageIntLLRInputS5xD(10)(1) <= VNStageIntLLROutputS4xD(109)(0);
  CNStageIntLLRInputS5xD(100)(1) <= VNStageIntLLROutputS4xD(109)(1);
  CNStageIntLLRInputS5xD(160)(1) <= VNStageIntLLROutputS4xD(109)(2);
  CNStageIntLLRInputS5xD(171)(1) <= VNStageIntLLROutputS4xD(109)(3);
  CNStageIntLLRInputS5xD(266)(1) <= VNStageIntLLROutputS4xD(109)(4);
  CNStageIntLLRInputS5xD(362)(1) <= VNStageIntLLROutputS4xD(109)(5);
  CNStageIntLLRInputS5xD(9)(1) <= VNStageIntLLROutputS4xD(110)(0);
  CNStageIntLLRInputS5xD(83)(1) <= VNStageIntLLROutputS4xD(110)(1);
  CNStageIntLLRInputS5xD(118)(1) <= VNStageIntLLROutputS4xD(110)(2);
  CNStageIntLLRInputS5xD(212)(1) <= VNStageIntLLROutputS4xD(110)(3);
  CNStageIntLLRInputS5xD(225)(1) <= VNStageIntLLROutputS4xD(110)(4);
  CNStageIntLLRInputS5xD(326)(1) <= VNStageIntLLROutputS4xD(110)(5);
  CNStageIntLLRInputS5xD(345)(1) <= VNStageIntLLROutputS4xD(110)(6);
  CNStageIntLLRInputS5xD(8)(1) <= VNStageIntLLROutputS4xD(111)(0);
  CNStageIntLLRInputS5xD(90)(1) <= VNStageIntLLROutputS4xD(111)(1);
  CNStageIntLLRInputS5xD(138)(1) <= VNStageIntLLROutputS4xD(111)(2);
  CNStageIntLLRInputS5xD(177)(1) <= VNStageIntLLROutputS4xD(111)(3);
  CNStageIntLLRInputS5xD(252)(1) <= VNStageIntLLROutputS4xD(111)(4);
  CNStageIntLLRInputS5xD(287)(1) <= VNStageIntLLROutputS4xD(111)(5);
  CNStageIntLLRInputS5xD(357)(1) <= VNStageIntLLROutputS4xD(111)(6);
  CNStageIntLLRInputS5xD(7)(1) <= VNStageIntLLROutputS4xD(112)(0);
  CNStageIntLLRInputS5xD(54)(1) <= VNStageIntLLROutputS4xD(112)(1);
  CNStageIntLLRInputS5xD(148)(1) <= VNStageIntLLROutputS4xD(112)(2);
  CNStageIntLLRInputS5xD(205)(1) <= VNStageIntLLROutputS4xD(112)(3);
  CNStageIntLLRInputS5xD(233)(1) <= VNStageIntLLROutputS4xD(112)(4);
  CNStageIntLLRInputS5xD(305)(1) <= VNStageIntLLROutputS4xD(112)(5);
  CNStageIntLLRInputS5xD(369)(1) <= VNStageIntLLROutputS4xD(112)(6);
  CNStageIntLLRInputS5xD(6)(1) <= VNStageIntLLROutputS4xD(113)(0);
  CNStageIntLLRInputS5xD(108)(1) <= VNStageIntLLROutputS4xD(113)(1);
  CNStageIntLLRInputS5xD(143)(1) <= VNStageIntLLROutputS4xD(113)(2);
  CNStageIntLLRInputS5xD(202)(1) <= VNStageIntLLROutputS4xD(113)(3);
  CNStageIntLLRInputS5xD(253)(1) <= VNStageIntLLROutputS4xD(113)(4);
  CNStageIntLLRInputS5xD(314)(1) <= VNStageIntLLROutputS4xD(113)(5);
  CNStageIntLLRInputS5xD(339)(1) <= VNStageIntLLROutputS4xD(113)(6);
  CNStageIntLLRInputS5xD(5)(1) <= VNStageIntLLROutputS4xD(114)(0);
  CNStageIntLLRInputS5xD(88)(1) <= VNStageIntLLROutputS4xD(114)(1);
  CNStageIntLLRInputS5xD(149)(1) <= VNStageIntLLROutputS4xD(114)(2);
  CNStageIntLLRInputS5xD(216)(1) <= VNStageIntLLROutputS4xD(114)(3);
  CNStageIntLLRInputS5xD(268)(1) <= VNStageIntLLROutputS4xD(114)(4);
  CNStageIntLLRInputS5xD(309)(1) <= VNStageIntLLROutputS4xD(114)(5);
  CNStageIntLLRInputS5xD(4)(1) <= VNStageIntLLROutputS4xD(115)(0);
  CNStageIntLLRInputS5xD(68)(1) <= VNStageIntLLROutputS4xD(115)(1);
  CNStageIntLLRInputS5xD(137)(1) <= VNStageIntLLROutputS4xD(115)(2);
  CNStageIntLLRInputS5xD(209)(1) <= VNStageIntLLROutputS4xD(115)(3);
  CNStageIntLLRInputS5xD(264)(1) <= VNStageIntLLROutputS4xD(115)(4);
  CNStageIntLLRInputS5xD(315)(1) <= VNStageIntLLROutputS4xD(115)(5);
  CNStageIntLLRInputS5xD(372)(1) <= VNStageIntLLROutputS4xD(115)(6);
  CNStageIntLLRInputS5xD(71)(1) <= VNStageIntLLROutputS4xD(116)(0);
  CNStageIntLLRInputS5xD(163)(1) <= VNStageIntLLROutputS4xD(116)(1);
  CNStageIntLLRInputS5xD(187)(1) <= VNStageIntLLROutputS4xD(116)(2);
  CNStageIntLLRInputS5xD(228)(1) <= VNStageIntLLROutputS4xD(116)(3);
  CNStageIntLLRInputS5xD(304)(1) <= VNStageIntLLROutputS4xD(116)(4);
  CNStageIntLLRInputS5xD(3)(1) <= VNStageIntLLROutputS4xD(117)(0);
  CNStageIntLLRInputS5xD(55)(1) <= VNStageIntLLROutputS4xD(117)(1);
  CNStageIntLLRInputS5xD(111)(1) <= VNStageIntLLROutputS4xD(117)(2);
  CNStageIntLLRInputS5xD(196)(1) <= VNStageIntLLROutputS4xD(117)(3);
  CNStageIntLLRInputS5xD(2)(1) <= VNStageIntLLROutputS4xD(118)(0);
  CNStageIntLLRInputS5xD(89)(1) <= VNStageIntLLROutputS4xD(118)(1);
  CNStageIntLLRInputS5xD(152)(1) <= VNStageIntLLROutputS4xD(118)(2);
  CNStageIntLLRInputS5xD(249)(1) <= VNStageIntLLROutputS4xD(118)(3);
  CNStageIntLLRInputS5xD(282)(1) <= VNStageIntLLROutputS4xD(118)(4);
  CNStageIntLLRInputS5xD(359)(1) <= VNStageIntLLROutputS4xD(118)(5);
  CNStageIntLLRInputS5xD(1)(1) <= VNStageIntLLROutputS4xD(119)(0);
  CNStageIntLLRInputS5xD(107)(1) <= VNStageIntLLROutputS4xD(119)(1);
  CNStageIntLLRInputS5xD(154)(1) <= VNStageIntLLROutputS4xD(119)(2);
  CNStageIntLLRInputS5xD(227)(1) <= VNStageIntLLROutputS4xD(119)(3);
  CNStageIntLLRInputS5xD(319)(1) <= VNStageIntLLROutputS4xD(119)(4);
  CNStageIntLLRInputS5xD(0)(1) <= VNStageIntLLROutputS4xD(120)(0);
  CNStageIntLLRInputS5xD(80)(1) <= VNStageIntLLROutputS4xD(120)(1);
  CNStageIntLLRInputS5xD(321)(1) <= VNStageIntLLROutputS4xD(120)(2);
  CNStageIntLLRInputS5xD(360)(1) <= VNStageIntLLROutputS4xD(120)(3);
  CNStageIntLLRInputS5xD(64)(1) <= VNStageIntLLROutputS4xD(121)(0);
  CNStageIntLLRInputS5xD(161)(1) <= VNStageIntLLROutputS4xD(121)(1);
  CNStageIntLLRInputS5xD(217)(1) <= VNStageIntLLROutputS4xD(121)(2);
  CNStageIntLLRInputS5xD(236)(1) <= VNStageIntLLROutputS4xD(121)(3);
  CNStageIntLLRInputS5xD(291)(1) <= VNStageIntLLROutputS4xD(121)(4);
  CNStageIntLLRInputS5xD(350)(1) <= VNStageIntLLROutputS4xD(121)(5);
  CNStageIntLLRInputS5xD(91)(1) <= VNStageIntLLROutputS4xD(122)(0);
  CNStageIntLLRInputS5xD(114)(1) <= VNStageIntLLROutputS4xD(122)(1);
  CNStageIntLLRInputS5xD(201)(1) <= VNStageIntLLROutputS4xD(122)(2);
  CNStageIntLLRInputS5xD(241)(1) <= VNStageIntLLROutputS4xD(122)(3);
  CNStageIntLLRInputS5xD(327)(1) <= VNStageIntLLROutputS4xD(122)(4);
  CNStageIntLLRInputS5xD(375)(1) <= VNStageIntLLROutputS4xD(122)(5);
  CNStageIntLLRInputS5xD(82)(1) <= VNStageIntLLROutputS4xD(123)(0);
  CNStageIntLLRInputS5xD(122)(1) <= VNStageIntLLROutputS4xD(123)(1);
  CNStageIntLLRInputS5xD(213)(1) <= VNStageIntLLROutputS4xD(123)(2);
  CNStageIntLLRInputS5xD(279)(1) <= VNStageIntLLROutputS4xD(123)(3);
  CNStageIntLLRInputS5xD(382)(1) <= VNStageIntLLROutputS4xD(123)(4);
  CNStageIntLLRInputS5xD(69)(1) <= VNStageIntLLROutputS4xD(124)(0);
  CNStageIntLLRInputS5xD(153)(1) <= VNStageIntLLROutputS4xD(124)(1);
  CNStageIntLLRInputS5xD(240)(1) <= VNStageIntLLROutputS4xD(124)(2);
  CNStageIntLLRInputS5xD(292)(1) <= VNStageIntLLROutputS4xD(124)(3);
  CNStageIntLLRInputS5xD(364)(1) <= VNStageIntLLROutputS4xD(124)(4);
  CNStageIntLLRInputS5xD(87)(1) <= VNStageIntLLROutputS4xD(125)(0);
  CNStageIntLLRInputS5xD(169)(1) <= VNStageIntLLROutputS4xD(125)(1);
  CNStageIntLLRInputS5xD(320)(1) <= VNStageIntLLROutputS4xD(125)(2);
  CNStageIntLLRInputS5xD(366)(1) <= VNStageIntLLROutputS4xD(125)(3);
  CNStageIntLLRInputS5xD(60)(1) <= VNStageIntLLROutputS4xD(126)(0);
  CNStageIntLLRInputS5xD(139)(1) <= VNStageIntLLROutputS4xD(126)(1);
  CNStageIntLLRInputS5xD(186)(1) <= VNStageIntLLROutputS4xD(126)(2);
  CNStageIntLLRInputS5xD(271)(1) <= VNStageIntLLROutputS4xD(126)(3);
  CNStageIntLLRInputS5xD(281)(1) <= VNStageIntLLROutputS4xD(126)(4);
  CNStageIntLLRInputS5xD(334)(1) <= VNStageIntLLROutputS4xD(126)(5);
  CNStageIntLLRInputS5xD(52)(1) <= VNStageIntLLROutputS4xD(127)(0);
  CNStageIntLLRInputS5xD(57)(1) <= VNStageIntLLROutputS4xD(127)(1);
  CNStageIntLLRInputS5xD(117)(1) <= VNStageIntLLROutputS4xD(127)(2);
  CNStageIntLLRInputS5xD(173)(1) <= VNStageIntLLROutputS4xD(127)(3);
  CNStageIntLLRInputS5xD(277)(1) <= VNStageIntLLROutputS4xD(127)(4);
  CNStageIntLLRInputS5xD(306)(1) <= VNStageIntLLROutputS4xD(127)(5);
  CNStageIntLLRInputS5xD(373)(1) <= VNStageIntLLROutputS4xD(127)(6);
  CNStageIntLLRInputS5xD(53)(2) <= VNStageIntLLROutputS4xD(128)(0);
  CNStageIntLLRInputS5xD(108)(2) <= VNStageIntLLROutputS4xD(128)(1);
  CNStageIntLLRInputS5xD(129)(2) <= VNStageIntLLROutputS4xD(128)(2);
  CNStageIntLLRInputS5xD(198)(2) <= VNStageIntLLROutputS4xD(128)(3);
  CNStageIntLLRInputS5xD(244)(2) <= VNStageIntLLROutputS4xD(128)(4);
  CNStageIntLLRInputS5xD(298)(2) <= VNStageIntLLROutputS4xD(128)(5);
  CNStageIntLLRInputS5xD(341)(2) <= VNStageIntLLROutputS4xD(128)(6);
  CNStageIntLLRInputS5xD(51)(2) <= VNStageIntLLROutputS4xD(129)(0);
  CNStageIntLLRInputS5xD(56)(2) <= VNStageIntLLROutputS4xD(129)(1);
  CNStageIntLLRInputS5xD(116)(2) <= VNStageIntLLROutputS4xD(129)(2);
  CNStageIntLLRInputS5xD(172)(2) <= VNStageIntLLROutputS4xD(129)(3);
  CNStageIntLLRInputS5xD(276)(2) <= VNStageIntLLROutputS4xD(129)(4);
  CNStageIntLLRInputS5xD(305)(2) <= VNStageIntLLROutputS4xD(129)(5);
  CNStageIntLLRInputS5xD(372)(2) <= VNStageIntLLROutputS4xD(129)(6);
  CNStageIntLLRInputS5xD(50)(2) <= VNStageIntLLROutputS4xD(130)(0);
  CNStageIntLLRInputS5xD(73)(2) <= VNStageIntLLROutputS4xD(130)(1);
  CNStageIntLLRInputS5xD(140)(2) <= VNStageIntLLROutputS4xD(130)(2);
  CNStageIntLLRInputS5xD(188)(2) <= VNStageIntLLROutputS4xD(130)(3);
  CNStageIntLLRInputS5xD(245)(2) <= VNStageIntLLROutputS4xD(130)(4);
  CNStageIntLLRInputS5xD(285)(2) <= VNStageIntLLROutputS4xD(130)(5);
  CNStageIntLLRInputS5xD(65)(2) <= VNStageIntLLROutputS4xD(131)(0);
  CNStageIntLLRInputS5xD(154)(2) <= VNStageIntLLROutputS4xD(131)(1);
  CNStageIntLLRInputS5xD(206)(2) <= VNStageIntLLROutputS4xD(131)(2);
  CNStageIntLLRInputS5xD(243)(2) <= VNStageIntLLROutputS4xD(131)(3);
  CNStageIntLLRInputS5xD(307)(2) <= VNStageIntLLROutputS4xD(131)(4);
  CNStageIntLLRInputS5xD(334)(2) <= VNStageIntLLROutputS4xD(131)(5);
  CNStageIntLLRInputS5xD(49)(2) <= VNStageIntLLROutputS4xD(132)(0);
  CNStageIntLLRInputS5xD(151)(2) <= VNStageIntLLROutputS4xD(132)(1);
  CNStageIntLLRInputS5xD(214)(2) <= VNStageIntLLROutputS4xD(132)(2);
  CNStageIntLLRInputS5xD(274)(2) <= VNStageIntLLROutputS4xD(132)(3);
  CNStageIntLLRInputS5xD(321)(2) <= VNStageIntLLROutputS4xD(132)(4);
  CNStageIntLLRInputS5xD(364)(2) <= VNStageIntLLROutputS4xD(132)(5);
  CNStageIntLLRInputS5xD(48)(2) <= VNStageIntLLROutputS4xD(133)(0);
  CNStageIntLLRInputS5xD(209)(2) <= VNStageIntLLROutputS4xD(133)(1);
  CNStageIntLLRInputS5xD(255)(2) <= VNStageIntLLROutputS4xD(133)(2);
  CNStageIntLLRInputS5xD(317)(2) <= VNStageIntLLROutputS4xD(133)(3);
  CNStageIntLLRInputS5xD(380)(2) <= VNStageIntLLROutputS4xD(133)(4);
  CNStageIntLLRInputS5xD(47)(2) <= VNStageIntLLROutputS4xD(134)(0);
  CNStageIntLLRInputS5xD(100)(2) <= VNStageIntLLROutputS4xD(134)(1);
  CNStageIntLLRInputS5xD(134)(2) <= VNStageIntLLROutputS4xD(134)(2);
  CNStageIntLLRInputS5xD(258)(2) <= VNStageIntLLROutputS4xD(134)(3);
  CNStageIntLLRInputS5xD(46)(2) <= VNStageIntLLROutputS4xD(135)(0);
  CNStageIntLLRInputS5xD(103)(2) <= VNStageIntLLROutputS4xD(135)(1);
  CNStageIntLLRInputS5xD(135)(2) <= VNStageIntLLROutputS4xD(135)(2);
  CNStageIntLLRInputS5xD(205)(2) <= VNStageIntLLROutputS4xD(135)(3);
  CNStageIntLLRInputS5xD(45)(2) <= VNStageIntLLROutputS4xD(136)(0);
  CNStageIntLLRInputS5xD(94)(2) <= VNStageIntLLROutputS4xD(136)(1);
  CNStageIntLLRInputS5xD(111)(2) <= VNStageIntLLROutputS4xD(136)(2);
  CNStageIntLLRInputS5xD(175)(2) <= VNStageIntLLROutputS4xD(136)(3);
  CNStageIntLLRInputS5xD(275)(2) <= VNStageIntLLROutputS4xD(136)(4);
  CNStageIntLLRInputS5xD(301)(2) <= VNStageIntLLROutputS4xD(136)(5);
  CNStageIntLLRInputS5xD(352)(2) <= VNStageIntLLROutputS4xD(136)(6);
  CNStageIntLLRInputS5xD(44)(2) <= VNStageIntLLROutputS4xD(137)(0);
  CNStageIntLLRInputS5xD(74)(2) <= VNStageIntLLROutputS4xD(137)(1);
  CNStageIntLLRInputS5xD(161)(2) <= VNStageIntLLROutputS4xD(137)(2);
  CNStageIntLLRInputS5xD(182)(2) <= VNStageIntLLROutputS4xD(137)(3);
  CNStageIntLLRInputS5xD(242)(2) <= VNStageIntLLROutputS4xD(137)(4);
  CNStageIntLLRInputS5xD(282)(2) <= VNStageIntLLROutputS4xD(137)(5);
  CNStageIntLLRInputS5xD(366)(2) <= VNStageIntLLROutputS4xD(137)(6);
  CNStageIntLLRInputS5xD(43)(2) <= VNStageIntLLROutputS4xD(138)(0);
  CNStageIntLLRInputS5xD(55)(2) <= VNStageIntLLROutputS4xD(138)(1);
  CNStageIntLLRInputS5xD(120)(2) <= VNStageIntLLROutputS4xD(138)(2);
  CNStageIntLLRInputS5xD(218)(2) <= VNStageIntLLROutputS4xD(138)(3);
  CNStageIntLLRInputS5xD(268)(2) <= VNStageIntLLROutputS4xD(138)(4);
  CNStageIntLLRInputS5xD(327)(2) <= VNStageIntLLROutputS4xD(138)(5);
  CNStageIntLLRInputS5xD(362)(2) <= VNStageIntLLROutputS4xD(138)(6);
  CNStageIntLLRInputS5xD(42)(2) <= VNStageIntLLROutputS4xD(139)(0);
  CNStageIntLLRInputS5xD(69)(2) <= VNStageIntLLROutputS4xD(139)(1);
  CNStageIntLLRInputS5xD(124)(2) <= VNStageIntLLROutputS4xD(139)(2);
  CNStageIntLLRInputS5xD(220)(2) <= VNStageIntLLROutputS4xD(139)(3);
  CNStageIntLLRInputS5xD(252)(2) <= VNStageIntLLROutputS4xD(139)(4);
  CNStageIntLLRInputS5xD(289)(2) <= VNStageIntLLROutputS4xD(139)(5);
  CNStageIntLLRInputS5xD(383)(2) <= VNStageIntLLROutputS4xD(139)(6);
  CNStageIntLLRInputS5xD(41)(2) <= VNStageIntLLROutputS4xD(140)(0);
  CNStageIntLLRInputS5xD(80)(2) <= VNStageIntLLROutputS4xD(140)(1);
  CNStageIntLLRInputS5xD(170)(2) <= VNStageIntLLROutputS4xD(140)(2);
  CNStageIntLLRInputS5xD(191)(2) <= VNStageIntLLROutputS4xD(140)(3);
  CNStageIntLLRInputS5xD(277)(2) <= VNStageIntLLROutputS4xD(140)(4);
  CNStageIntLLRInputS5xD(293)(2) <= VNStageIntLLROutputS4xD(140)(5);
  CNStageIntLLRInputS5xD(346)(2) <= VNStageIntLLROutputS4xD(140)(6);
  CNStageIntLLRInputS5xD(123)(2) <= VNStageIntLLROutputS4xD(141)(0);
  CNStageIntLLRInputS5xD(173)(2) <= VNStageIntLLROutputS4xD(141)(1);
  CNStageIntLLRInputS5xD(269)(2) <= VNStageIntLLROutputS4xD(141)(2);
  CNStageIntLLRInputS5xD(332)(2) <= VNStageIntLLROutputS4xD(141)(3);
  CNStageIntLLRInputS5xD(347)(2) <= VNStageIntLLROutputS4xD(141)(4);
  CNStageIntLLRInputS5xD(40)(2) <= VNStageIntLLROutputS4xD(142)(0);
  CNStageIntLLRInputS5xD(96)(2) <= VNStageIntLLROutputS4xD(142)(1);
  CNStageIntLLRInputS5xD(118)(2) <= VNStageIntLLROutputS4xD(142)(2);
  CNStageIntLLRInputS5xD(256)(2) <= VNStageIntLLROutputS4xD(142)(3);
  CNStageIntLLRInputS5xD(382)(2) <= VNStageIntLLROutputS4xD(142)(4);
  CNStageIntLLRInputS5xD(39)(2) <= VNStageIntLLROutputS4xD(143)(0);
  CNStageIntLLRInputS5xD(83)(2) <= VNStageIntLLROutputS4xD(143)(1);
  CNStageIntLLRInputS5xD(158)(2) <= VNStageIntLLROutputS4xD(143)(2);
  CNStageIntLLRInputS5xD(192)(2) <= VNStageIntLLROutputS4xD(143)(3);
  CNStageIntLLRInputS5xD(273)(2) <= VNStageIntLLROutputS4xD(143)(4);
  CNStageIntLLRInputS5xD(287)(2) <= VNStageIntLLROutputS4xD(143)(5);
  CNStageIntLLRInputS5xD(373)(2) <= VNStageIntLLROutputS4xD(143)(6);
  CNStageIntLLRInputS5xD(38)(2) <= VNStageIntLLROutputS4xD(144)(0);
  CNStageIntLLRInputS5xD(98)(2) <= VNStageIntLLROutputS4xD(144)(1);
  CNStageIntLLRInputS5xD(166)(2) <= VNStageIntLLROutputS4xD(144)(2);
  CNStageIntLLRInputS5xD(219)(2) <= VNStageIntLLROutputS4xD(144)(3);
  CNStageIntLLRInputS5xD(249)(2) <= VNStageIntLLROutputS4xD(144)(4);
  CNStageIntLLRInputS5xD(324)(2) <= VNStageIntLLROutputS4xD(144)(5);
  CNStageIntLLRInputS5xD(333)(2) <= VNStageIntLLROutputS4xD(144)(6);
  CNStageIntLLRInputS5xD(37)(2) <= VNStageIntLLROutputS4xD(145)(0);
  CNStageIntLLRInputS5xD(61)(2) <= VNStageIntLLROutputS4xD(145)(1);
  CNStageIntLLRInputS5xD(130)(2) <= VNStageIntLLROutputS4xD(145)(2);
  CNStageIntLLRInputS5xD(181)(2) <= VNStageIntLLROutputS4xD(145)(3);
  CNStageIntLLRInputS5xD(247)(2) <= VNStageIntLLROutputS4xD(145)(4);
  CNStageIntLLRInputS5xD(331)(2) <= VNStageIntLLROutputS4xD(145)(5);
  CNStageIntLLRInputS5xD(336)(2) <= VNStageIntLLROutputS4xD(145)(6);
  CNStageIntLLRInputS5xD(36)(2) <= VNStageIntLLROutputS4xD(146)(0);
  CNStageIntLLRInputS5xD(71)(2) <= VNStageIntLLROutputS4xD(146)(1);
  CNStageIntLLRInputS5xD(128)(2) <= VNStageIntLLROutputS4xD(146)(2);
  CNStageIntLLRInputS5xD(261)(2) <= VNStageIntLLROutputS4xD(146)(3);
  CNStageIntLLRInputS5xD(299)(2) <= VNStageIntLLROutputS4xD(146)(4);
  CNStageIntLLRInputS5xD(35)(2) <= VNStageIntLLROutputS4xD(147)(0);
  CNStageIntLLRInputS5xD(66)(2) <= VNStageIntLLROutputS4xD(147)(1);
  CNStageIntLLRInputS5xD(164)(2) <= VNStageIntLLROutputS4xD(147)(2);
  CNStageIntLLRInputS5xD(187)(2) <= VNStageIntLLROutputS4xD(147)(3);
  CNStageIntLLRInputS5xD(253)(2) <= VNStageIntLLROutputS4xD(147)(4);
  CNStageIntLLRInputS5xD(297)(2) <= VNStageIntLLROutputS4xD(147)(5);
  CNStageIntLLRInputS5xD(335)(2) <= VNStageIntLLROutputS4xD(147)(6);
  CNStageIntLLRInputS5xD(34)(2) <= VNStageIntLLROutputS4xD(148)(0);
  CNStageIntLLRInputS5xD(72)(2) <= VNStageIntLLROutputS4xD(148)(1);
  CNStageIntLLRInputS5xD(143)(2) <= VNStageIntLLROutputS4xD(148)(2);
  CNStageIntLLRInputS5xD(207)(2) <= VNStageIntLLROutputS4xD(148)(3);
  CNStageIntLLRInputS5xD(231)(2) <= VNStageIntLLROutputS4xD(148)(4);
  CNStageIntLLRInputS5xD(329)(2) <= VNStageIntLLROutputS4xD(148)(5);
  CNStageIntLLRInputS5xD(33)(2) <= VNStageIntLLROutputS4xD(149)(0);
  CNStageIntLLRInputS5xD(60)(2) <= VNStageIntLLROutputS4xD(149)(1);
  CNStageIntLLRInputS5xD(146)(2) <= VNStageIntLLROutputS4xD(149)(2);
  CNStageIntLLRInputS5xD(221)(2) <= VNStageIntLLROutputS4xD(149)(3);
  CNStageIntLLRInputS5xD(241)(2) <= VNStageIntLLROutputS4xD(149)(4);
  CNStageIntLLRInputS5xD(309)(2) <= VNStageIntLLROutputS4xD(149)(5);
  CNStageIntLLRInputS5xD(370)(2) <= VNStageIntLLROutputS4xD(149)(6);
  CNStageIntLLRInputS5xD(32)(2) <= VNStageIntLLROutputS4xD(150)(0);
  CNStageIntLLRInputS5xD(86)(2) <= VNStageIntLLROutputS4xD(150)(1);
  CNStageIntLLRInputS5xD(131)(2) <= VNStageIntLLROutputS4xD(150)(2);
  CNStageIntLLRInputS5xD(217)(2) <= VNStageIntLLROutputS4xD(150)(3);
  CNStageIntLLRInputS5xD(312)(2) <= VNStageIntLLROutputS4xD(150)(4);
  CNStageIntLLRInputS5xD(378)(2) <= VNStageIntLLROutputS4xD(150)(5);
  CNStageIntLLRInputS5xD(31)(2) <= VNStageIntLLROutputS4xD(151)(0);
  CNStageIntLLRInputS5xD(92)(2) <= VNStageIntLLROutputS4xD(151)(1);
  CNStageIntLLRInputS5xD(165)(2) <= VNStageIntLLROutputS4xD(151)(2);
  CNStageIntLLRInputS5xD(184)(2) <= VNStageIntLLROutputS4xD(151)(3);
  CNStageIntLLRInputS5xD(238)(2) <= VNStageIntLLROutputS4xD(151)(4);
  CNStageIntLLRInputS5xD(342)(2) <= VNStageIntLLROutputS4xD(151)(5);
  CNStageIntLLRInputS5xD(30)(2) <= VNStageIntLLROutputS4xD(152)(0);
  CNStageIntLLRInputS5xD(76)(2) <= VNStageIntLLROutputS4xD(152)(1);
  CNStageIntLLRInputS5xD(127)(2) <= VNStageIntLLROutputS4xD(152)(2);
  CNStageIntLLRInputS5xD(202)(2) <= VNStageIntLLROutputS4xD(152)(3);
  CNStageIntLLRInputS5xD(228)(2) <= VNStageIntLLROutputS4xD(152)(4);
  CNStageIntLLRInputS5xD(330)(2) <= VNStageIntLLROutputS4xD(152)(5);
  CNStageIntLLRInputS5xD(340)(2) <= VNStageIntLLROutputS4xD(152)(6);
  CNStageIntLLRInputS5xD(29)(2) <= VNStageIntLLROutputS4xD(153)(0);
  CNStageIntLLRInputS5xD(78)(2) <= VNStageIntLLROutputS4xD(153)(1);
  CNStageIntLLRInputS5xD(155)(2) <= VNStageIntLLROutputS4xD(153)(2);
  CNStageIntLLRInputS5xD(203)(2) <= VNStageIntLLROutputS4xD(153)(3);
  CNStageIntLLRInputS5xD(262)(2) <= VNStageIntLLROutputS4xD(153)(4);
  CNStageIntLLRInputS5xD(296)(2) <= VNStageIntLLROutputS4xD(153)(5);
  CNStageIntLLRInputS5xD(376)(2) <= VNStageIntLLROutputS4xD(153)(6);
  CNStageIntLLRInputS5xD(28)(2) <= VNStageIntLLROutputS4xD(154)(0);
  CNStageIntLLRInputS5xD(139)(2) <= VNStageIntLLROutputS4xD(154)(1);
  CNStageIntLLRInputS5xD(183)(2) <= VNStageIntLLROutputS4xD(154)(2);
  CNStageIntLLRInputS5xD(246)(2) <= VNStageIntLLROutputS4xD(154)(3);
  CNStageIntLLRInputS5xD(322)(2) <= VNStageIntLLROutputS4xD(154)(4);
  CNStageIntLLRInputS5xD(27)(2) <= VNStageIntLLROutputS4xD(155)(0);
  CNStageIntLLRInputS5xD(84)(2) <= VNStageIntLLROutputS4xD(155)(1);
  CNStageIntLLRInputS5xD(167)(2) <= VNStageIntLLROutputS4xD(155)(2);
  CNStageIntLLRInputS5xD(174)(2) <= VNStageIntLLROutputS4xD(155)(3);
  CNStageIntLLRInputS5xD(257)(2) <= VNStageIntLLROutputS4xD(155)(4);
  CNStageIntLLRInputS5xD(306)(2) <= VNStageIntLLROutputS4xD(155)(5);
  CNStageIntLLRInputS5xD(357)(2) <= VNStageIntLLROutputS4xD(155)(6);
  CNStageIntLLRInputS5xD(26)(2) <= VNStageIntLLROutputS4xD(156)(0);
  CNStageIntLLRInputS5xD(95)(2) <= VNStageIntLLROutputS4xD(156)(1);
  CNStageIntLLRInputS5xD(157)(2) <= VNStageIntLLROutputS4xD(156)(2);
  CNStageIntLLRInputS5xD(343)(2) <= VNStageIntLLROutputS4xD(156)(3);
  CNStageIntLLRInputS5xD(25)(2) <= VNStageIntLLROutputS4xD(157)(0);
  CNStageIntLLRInputS5xD(102)(2) <= VNStageIntLLROutputS4xD(157)(1);
  CNStageIntLLRInputS5xD(144)(2) <= VNStageIntLLROutputS4xD(157)(2);
  CNStageIntLLRInputS5xD(194)(2) <= VNStageIntLLROutputS4xD(157)(3);
  CNStageIntLLRInputS5xD(323)(2) <= VNStageIntLLROutputS4xD(157)(4);
  CNStageIntLLRInputS5xD(377)(2) <= VNStageIntLLROutputS4xD(157)(5);
  CNStageIntLLRInputS5xD(24)(2) <= VNStageIntLLROutputS4xD(158)(0);
  CNStageIntLLRInputS5xD(77)(2) <= VNStageIntLLROutputS4xD(158)(1);
  CNStageIntLLRInputS5xD(163)(2) <= VNStageIntLLROutputS4xD(158)(2);
  CNStageIntLLRInputS5xD(224)(2) <= VNStageIntLLROutputS4xD(158)(3);
  CNStageIntLLRInputS5xD(230)(2) <= VNStageIntLLROutputS4xD(158)(4);
  CNStageIntLLRInputS5xD(310)(2) <= VNStageIntLLROutputS4xD(158)(5);
  CNStageIntLLRInputS5xD(339)(2) <= VNStageIntLLROutputS4xD(158)(6);
  CNStageIntLLRInputS5xD(23)(2) <= VNStageIntLLROutputS4xD(159)(0);
  CNStageIntLLRInputS5xD(91)(2) <= VNStageIntLLROutputS4xD(159)(1);
  CNStageIntLLRInputS5xD(136)(2) <= VNStageIntLLROutputS4xD(159)(2);
  CNStageIntLLRInputS5xD(271)(2) <= VNStageIntLLROutputS4xD(159)(3);
  CNStageIntLLRInputS5xD(367)(2) <= VNStageIntLLROutputS4xD(159)(4);
  CNStageIntLLRInputS5xD(22)(2) <= VNStageIntLLROutputS4xD(160)(0);
  CNStageIntLLRInputS5xD(62)(2) <= VNStageIntLLROutputS4xD(160)(1);
  CNStageIntLLRInputS5xD(133)(2) <= VNStageIntLLROutputS4xD(160)(2);
  CNStageIntLLRInputS5xD(189)(2) <= VNStageIntLLROutputS4xD(160)(3);
  CNStageIntLLRInputS5xD(233)(2) <= VNStageIntLLROutputS4xD(160)(4);
  CNStageIntLLRInputS5xD(302)(2) <= VNStageIntLLROutputS4xD(160)(5);
  CNStageIntLLRInputS5xD(351)(2) <= VNStageIntLLROutputS4xD(160)(6);
  CNStageIntLLRInputS5xD(21)(2) <= VNStageIntLLROutputS4xD(161)(0);
  CNStageIntLLRInputS5xD(97)(2) <= VNStageIntLLROutputS4xD(161)(1);
  CNStageIntLLRInputS5xD(149)(2) <= VNStageIntLLROutputS4xD(161)(2);
  CNStageIntLLRInputS5xD(171)(2) <= VNStageIntLLROutputS4xD(161)(3);
  CNStageIntLLRInputS5xD(250)(2) <= VNStageIntLLROutputS4xD(161)(4);
  CNStageIntLLRInputS5xD(300)(2) <= VNStageIntLLROutputS4xD(161)(5);
  CNStageIntLLRInputS5xD(379)(2) <= VNStageIntLLROutputS4xD(161)(6);
  CNStageIntLLRInputS5xD(20)(2) <= VNStageIntLLROutputS4xD(162)(0);
  CNStageIntLLRInputS5xD(64)(2) <= VNStageIntLLROutputS4xD(162)(1);
  CNStageIntLLRInputS5xD(141)(2) <= VNStageIntLLROutputS4xD(162)(2);
  CNStageIntLLRInputS5xD(179)(2) <= VNStageIntLLROutputS4xD(162)(3);
  CNStageIntLLRInputS5xD(259)(2) <= VNStageIntLLROutputS4xD(162)(4);
  CNStageIntLLRInputS5xD(315)(2) <= VNStageIntLLROutputS4xD(162)(5);
  CNStageIntLLRInputS5xD(369)(2) <= VNStageIntLLROutputS4xD(162)(6);
  CNStageIntLLRInputS5xD(19)(2) <= VNStageIntLLROutputS4xD(163)(0);
  CNStageIntLLRInputS5xD(79)(2) <= VNStageIntLLROutputS4xD(163)(1);
  CNStageIntLLRInputS5xD(115)(2) <= VNStageIntLLROutputS4xD(163)(2);
  CNStageIntLLRInputS5xD(254)(2) <= VNStageIntLLROutputS4xD(163)(3);
  CNStageIntLLRInputS5xD(355)(2) <= VNStageIntLLROutputS4xD(163)(4);
  CNStageIntLLRInputS5xD(18)(2) <= VNStageIntLLROutputS4xD(164)(0);
  CNStageIntLLRInputS5xD(75)(2) <= VNStageIntLLROutputS4xD(164)(1);
  CNStageIntLLRInputS5xD(125)(2) <= VNStageIntLLROutputS4xD(164)(2);
  CNStageIntLLRInputS5xD(197)(2) <= VNStageIntLLROutputS4xD(164)(3);
  CNStageIntLLRInputS5xD(260)(2) <= VNStageIntLLROutputS4xD(164)(4);
  CNStageIntLLRInputS5xD(375)(2) <= VNStageIntLLROutputS4xD(164)(5);
  CNStageIntLLRInputS5xD(17)(2) <= VNStageIntLLROutputS4xD(165)(0);
  CNStageIntLLRInputS5xD(93)(2) <= VNStageIntLLROutputS4xD(165)(1);
  CNStageIntLLRInputS5xD(119)(2) <= VNStageIntLLROutputS4xD(165)(2);
  CNStageIntLLRInputS5xD(177)(2) <= VNStageIntLLROutputS4xD(165)(3);
  CNStageIntLLRInputS5xD(294)(2) <= VNStageIntLLROutputS4xD(165)(4);
  CNStageIntLLRInputS5xD(348)(2) <= VNStageIntLLROutputS4xD(165)(5);
  CNStageIntLLRInputS5xD(16)(2) <= VNStageIntLLROutputS4xD(166)(0);
  CNStageIntLLRInputS5xD(57)(2) <= VNStageIntLLROutputS4xD(166)(1);
  CNStageIntLLRInputS5xD(122)(2) <= VNStageIntLLROutputS4xD(166)(2);
  CNStageIntLLRInputS5xD(210)(2) <= VNStageIntLLROutputS4xD(166)(3);
  CNStageIntLLRInputS5xD(288)(2) <= VNStageIntLLROutputS4xD(166)(4);
  CNStageIntLLRInputS5xD(345)(2) <= VNStageIntLLROutputS4xD(166)(5);
  CNStageIntLLRInputS5xD(15)(2) <= VNStageIntLLROutputS4xD(167)(0);
  CNStageIntLLRInputS5xD(58)(2) <= VNStageIntLLROutputS4xD(167)(1);
  CNStageIntLLRInputS5xD(112)(2) <= VNStageIntLLROutputS4xD(167)(2);
  CNStageIntLLRInputS5xD(213)(2) <= VNStageIntLLROutputS4xD(167)(3);
  CNStageIntLLRInputS5xD(225)(2) <= VNStageIntLLROutputS4xD(167)(4);
  CNStageIntLLRInputS5xD(292)(2) <= VNStageIntLLROutputS4xD(167)(5);
  CNStageIntLLRInputS5xD(360)(2) <= VNStageIntLLROutputS4xD(167)(6);
  CNStageIntLLRInputS5xD(14)(2) <= VNStageIntLLROutputS4xD(168)(0);
  CNStageIntLLRInputS5xD(150)(2) <= VNStageIntLLROutputS4xD(168)(1);
  CNStageIntLLRInputS5xD(199)(2) <= VNStageIntLLROutputS4xD(168)(2);
  CNStageIntLLRInputS5xD(264)(2) <= VNStageIntLLROutputS4xD(168)(3);
  CNStageIntLLRInputS5xD(283)(2) <= VNStageIntLLROutputS4xD(168)(4);
  CNStageIntLLRInputS5xD(353)(2) <= VNStageIntLLROutputS4xD(168)(5);
  CNStageIntLLRInputS5xD(13)(2) <= VNStageIntLLROutputS4xD(169)(0);
  CNStageIntLLRInputS5xD(85)(2) <= VNStageIntLLROutputS4xD(169)(1);
  CNStageIntLLRInputS5xD(132)(2) <= VNStageIntLLROutputS4xD(169)(2);
  CNStageIntLLRInputS5xD(178)(2) <= VNStageIntLLROutputS4xD(169)(3);
  CNStageIntLLRInputS5xD(266)(2) <= VNStageIntLLROutputS4xD(169)(4);
  CNStageIntLLRInputS5xD(316)(2) <= VNStageIntLLROutputS4xD(169)(5);
  CNStageIntLLRInputS5xD(12)(2) <= VNStageIntLLROutputS4xD(170)(0);
  CNStageIntLLRInputS5xD(101)(2) <= VNStageIntLLROutputS4xD(170)(1);
  CNStageIntLLRInputS5xD(145)(2) <= VNStageIntLLROutputS4xD(170)(2);
  CNStageIntLLRInputS5xD(236)(2) <= VNStageIntLLROutputS4xD(170)(3);
  CNStageIntLLRInputS5xD(337)(2) <= VNStageIntLLROutputS4xD(170)(4);
  CNStageIntLLRInputS5xD(105)(2) <= VNStageIntLLROutputS4xD(171)(0);
  CNStageIntLLRInputS5xD(156)(2) <= VNStageIntLLROutputS4xD(171)(1);
  CNStageIntLLRInputS5xD(222)(2) <= VNStageIntLLROutputS4xD(171)(2);
  CNStageIntLLRInputS5xD(311)(2) <= VNStageIntLLROutputS4xD(171)(3);
  CNStageIntLLRInputS5xD(11)(2) <= VNStageIntLLROutputS4xD(172)(0);
  CNStageIntLLRInputS5xD(110)(2) <= VNStageIntLLROutputS4xD(172)(1);
  CNStageIntLLRInputS5xD(126)(2) <= VNStageIntLLROutputS4xD(172)(2);
  CNStageIntLLRInputS5xD(229)(2) <= VNStageIntLLROutputS4xD(172)(3);
  CNStageIntLLRInputS5xD(10)(2) <= VNStageIntLLROutputS4xD(173)(0);
  CNStageIntLLRInputS5xD(104)(2) <= VNStageIntLLROutputS4xD(173)(1);
  CNStageIntLLRInputS5xD(114)(2) <= VNStageIntLLROutputS4xD(173)(2);
  CNStageIntLLRInputS5xD(180)(2) <= VNStageIntLLROutputS4xD(173)(3);
  CNStageIntLLRInputS5xD(237)(2) <= VNStageIntLLROutputS4xD(173)(4);
  CNStageIntLLRInputS5xD(295)(2) <= VNStageIntLLROutputS4xD(173)(5);
  CNStageIntLLRInputS5xD(9)(2) <= VNStageIntLLROutputS4xD(174)(0);
  CNStageIntLLRInputS5xD(99)(2) <= VNStageIntLLROutputS4xD(174)(1);
  CNStageIntLLRInputS5xD(159)(2) <= VNStageIntLLROutputS4xD(174)(2);
  CNStageIntLLRInputS5xD(265)(2) <= VNStageIntLLROutputS4xD(174)(3);
  CNStageIntLLRInputS5xD(361)(2) <= VNStageIntLLROutputS4xD(174)(4);
  CNStageIntLLRInputS5xD(8)(2) <= VNStageIntLLROutputS4xD(175)(0);
  CNStageIntLLRInputS5xD(82)(2) <= VNStageIntLLROutputS4xD(175)(1);
  CNStageIntLLRInputS5xD(117)(2) <= VNStageIntLLROutputS4xD(175)(2);
  CNStageIntLLRInputS5xD(211)(2) <= VNStageIntLLROutputS4xD(175)(3);
  CNStageIntLLRInputS5xD(278)(2) <= VNStageIntLLROutputS4xD(175)(4);
  CNStageIntLLRInputS5xD(325)(2) <= VNStageIntLLROutputS4xD(175)(5);
  CNStageIntLLRInputS5xD(344)(2) <= VNStageIntLLROutputS4xD(175)(6);
  CNStageIntLLRInputS5xD(7)(2) <= VNStageIntLLROutputS4xD(176)(0);
  CNStageIntLLRInputS5xD(89)(2) <= VNStageIntLLROutputS4xD(176)(1);
  CNStageIntLLRInputS5xD(137)(2) <= VNStageIntLLROutputS4xD(176)(2);
  CNStageIntLLRInputS5xD(176)(2) <= VNStageIntLLROutputS4xD(176)(3);
  CNStageIntLLRInputS5xD(251)(2) <= VNStageIntLLROutputS4xD(176)(4);
  CNStageIntLLRInputS5xD(286)(2) <= VNStageIntLLROutputS4xD(176)(5);
  CNStageIntLLRInputS5xD(356)(2) <= VNStageIntLLROutputS4xD(176)(6);
  CNStageIntLLRInputS5xD(6)(2) <= VNStageIntLLROutputS4xD(177)(0);
  CNStageIntLLRInputS5xD(109)(2) <= VNStageIntLLROutputS4xD(177)(1);
  CNStageIntLLRInputS5xD(147)(2) <= VNStageIntLLROutputS4xD(177)(2);
  CNStageIntLLRInputS5xD(204)(2) <= VNStageIntLLROutputS4xD(177)(3);
  CNStageIntLLRInputS5xD(232)(2) <= VNStageIntLLROutputS4xD(177)(4);
  CNStageIntLLRInputS5xD(304)(2) <= VNStageIntLLROutputS4xD(177)(5);
  CNStageIntLLRInputS5xD(368)(2) <= VNStageIntLLROutputS4xD(177)(6);
  CNStageIntLLRInputS5xD(5)(2) <= VNStageIntLLROutputS4xD(178)(0);
  CNStageIntLLRInputS5xD(107)(2) <= VNStageIntLLROutputS4xD(178)(1);
  CNStageIntLLRInputS5xD(142)(2) <= VNStageIntLLROutputS4xD(178)(2);
  CNStageIntLLRInputS5xD(201)(2) <= VNStageIntLLROutputS4xD(178)(3);
  CNStageIntLLRInputS5xD(313)(2) <= VNStageIntLLROutputS4xD(178)(4);
  CNStageIntLLRInputS5xD(338)(2) <= VNStageIntLLROutputS4xD(178)(5);
  CNStageIntLLRInputS5xD(4)(2) <= VNStageIntLLROutputS4xD(179)(0);
  CNStageIntLLRInputS5xD(87)(2) <= VNStageIntLLROutputS4xD(179)(1);
  CNStageIntLLRInputS5xD(148)(2) <= VNStageIntLLROutputS4xD(179)(2);
  CNStageIntLLRInputS5xD(215)(2) <= VNStageIntLLROutputS4xD(179)(3);
  CNStageIntLLRInputS5xD(267)(2) <= VNStageIntLLROutputS4xD(179)(4);
  CNStageIntLLRInputS5xD(308)(2) <= VNStageIntLLROutputS4xD(179)(5);
  CNStageIntLLRInputS5xD(67)(2) <= VNStageIntLLROutputS4xD(180)(0);
  CNStageIntLLRInputS5xD(208)(2) <= VNStageIntLLROutputS4xD(180)(1);
  CNStageIntLLRInputS5xD(263)(2) <= VNStageIntLLROutputS4xD(180)(2);
  CNStageIntLLRInputS5xD(314)(2) <= VNStageIntLLROutputS4xD(180)(3);
  CNStageIntLLRInputS5xD(371)(2) <= VNStageIntLLROutputS4xD(180)(4);
  CNStageIntLLRInputS5xD(3)(2) <= VNStageIntLLROutputS4xD(181)(0);
  CNStageIntLLRInputS5xD(70)(2) <= VNStageIntLLROutputS4xD(181)(1);
  CNStageIntLLRInputS5xD(162)(2) <= VNStageIntLLROutputS4xD(181)(2);
  CNStageIntLLRInputS5xD(186)(2) <= VNStageIntLLROutputS4xD(181)(3);
  CNStageIntLLRInputS5xD(227)(2) <= VNStageIntLLROutputS4xD(181)(4);
  CNStageIntLLRInputS5xD(303)(2) <= VNStageIntLLROutputS4xD(181)(5);
  CNStageIntLLRInputS5xD(2)(2) <= VNStageIntLLROutputS4xD(182)(0);
  CNStageIntLLRInputS5xD(54)(2) <= VNStageIntLLROutputS4xD(182)(1);
  CNStageIntLLRInputS5xD(169)(2) <= VNStageIntLLROutputS4xD(182)(2);
  CNStageIntLLRInputS5xD(195)(2) <= VNStageIntLLROutputS4xD(182)(3);
  CNStageIntLLRInputS5xD(248)(2) <= VNStageIntLLROutputS4xD(182)(4);
  CNStageIntLLRInputS5xD(328)(2) <= VNStageIntLLROutputS4xD(182)(5);
  CNStageIntLLRInputS5xD(350)(2) <= VNStageIntLLROutputS4xD(182)(6);
  CNStageIntLLRInputS5xD(1)(2) <= VNStageIntLLROutputS4xD(183)(0);
  CNStageIntLLRInputS5xD(88)(2) <= VNStageIntLLROutputS4xD(183)(1);
  CNStageIntLLRInputS5xD(190)(2) <= VNStageIntLLROutputS4xD(183)(2);
  CNStageIntLLRInputS5xD(281)(2) <= VNStageIntLLROutputS4xD(183)(3);
  CNStageIntLLRInputS5xD(358)(2) <= VNStageIntLLROutputS4xD(183)(4);
  CNStageIntLLRInputS5xD(0)(2) <= VNStageIntLLROutputS4xD(184)(0);
  CNStageIntLLRInputS5xD(106)(2) <= VNStageIntLLROutputS4xD(184)(1);
  CNStageIntLLRInputS5xD(153)(2) <= VNStageIntLLROutputS4xD(184)(2);
  CNStageIntLLRInputS5xD(193)(2) <= VNStageIntLLROutputS4xD(184)(3);
  CNStageIntLLRInputS5xD(226)(2) <= VNStageIntLLROutputS4xD(184)(4);
  CNStageIntLLRInputS5xD(318)(2) <= VNStageIntLLROutputS4xD(184)(5);
  CNStageIntLLRInputS5xD(354)(2) <= VNStageIntLLROutputS4xD(184)(6);
  CNStageIntLLRInputS5xD(121)(2) <= VNStageIntLLROutputS4xD(185)(0);
  CNStageIntLLRInputS5xD(272)(2) <= VNStageIntLLROutputS4xD(185)(1);
  CNStageIntLLRInputS5xD(320)(2) <= VNStageIntLLROutputS4xD(185)(2);
  CNStageIntLLRInputS5xD(359)(2) <= VNStageIntLLROutputS4xD(185)(3);
  CNStageIntLLRInputS5xD(63)(2) <= VNStageIntLLROutputS4xD(186)(0);
  CNStageIntLLRInputS5xD(160)(2) <= VNStageIntLLROutputS4xD(186)(1);
  CNStageIntLLRInputS5xD(216)(2) <= VNStageIntLLROutputS4xD(186)(2);
  CNStageIntLLRInputS5xD(235)(2) <= VNStageIntLLROutputS4xD(186)(3);
  CNStageIntLLRInputS5xD(290)(2) <= VNStageIntLLROutputS4xD(186)(4);
  CNStageIntLLRInputS5xD(349)(2) <= VNStageIntLLROutputS4xD(186)(5);
  CNStageIntLLRInputS5xD(90)(2) <= VNStageIntLLROutputS4xD(187)(0);
  CNStageIntLLRInputS5xD(113)(2) <= VNStageIntLLROutputS4xD(187)(1);
  CNStageIntLLRInputS5xD(200)(2) <= VNStageIntLLROutputS4xD(187)(2);
  CNStageIntLLRInputS5xD(240)(2) <= VNStageIntLLROutputS4xD(187)(3);
  CNStageIntLLRInputS5xD(326)(2) <= VNStageIntLLROutputS4xD(187)(4);
  CNStageIntLLRInputS5xD(374)(2) <= VNStageIntLLROutputS4xD(187)(5);
  CNStageIntLLRInputS5xD(81)(2) <= VNStageIntLLROutputS4xD(188)(0);
  CNStageIntLLRInputS5xD(212)(2) <= VNStageIntLLROutputS4xD(188)(1);
  CNStageIntLLRInputS5xD(279)(2) <= VNStageIntLLROutputS4xD(188)(2);
  CNStageIntLLRInputS5xD(284)(2) <= VNStageIntLLROutputS4xD(188)(3);
  CNStageIntLLRInputS5xD(381)(2) <= VNStageIntLLROutputS4xD(188)(4);
  CNStageIntLLRInputS5xD(68)(2) <= VNStageIntLLROutputS4xD(189)(0);
  CNStageIntLLRInputS5xD(152)(2) <= VNStageIntLLROutputS4xD(189)(1);
  CNStageIntLLRInputS5xD(223)(2) <= VNStageIntLLROutputS4xD(189)(2);
  CNStageIntLLRInputS5xD(239)(2) <= VNStageIntLLROutputS4xD(189)(3);
  CNStageIntLLRInputS5xD(291)(2) <= VNStageIntLLROutputS4xD(189)(4);
  CNStageIntLLRInputS5xD(363)(2) <= VNStageIntLLROutputS4xD(189)(5);
  CNStageIntLLRInputS5xD(168)(2) <= VNStageIntLLROutputS4xD(190)(0);
  CNStageIntLLRInputS5xD(196)(2) <= VNStageIntLLROutputS4xD(190)(1);
  CNStageIntLLRInputS5xD(234)(2) <= VNStageIntLLROutputS4xD(190)(2);
  CNStageIntLLRInputS5xD(319)(2) <= VNStageIntLLROutputS4xD(190)(3);
  CNStageIntLLRInputS5xD(365)(2) <= VNStageIntLLROutputS4xD(190)(4);
  CNStageIntLLRInputS5xD(52)(2) <= VNStageIntLLROutputS4xD(191)(0);
  CNStageIntLLRInputS5xD(59)(2) <= VNStageIntLLROutputS4xD(191)(1);
  CNStageIntLLRInputS5xD(138)(2) <= VNStageIntLLROutputS4xD(191)(2);
  CNStageIntLLRInputS5xD(185)(2) <= VNStageIntLLROutputS4xD(191)(3);
  CNStageIntLLRInputS5xD(270)(2) <= VNStageIntLLROutputS4xD(191)(4);
  CNStageIntLLRInputS5xD(280)(2) <= VNStageIntLLROutputS4xD(191)(5);
  CNStageIntLLRInputS5xD(53)(3) <= VNStageIntLLROutputS4xD(192)(0);
  CNStageIntLLRInputS5xD(107)(3) <= VNStageIntLLROutputS4xD(192)(1);
  CNStageIntLLRInputS5xD(128)(3) <= VNStageIntLLROutputS4xD(192)(2);
  CNStageIntLLRInputS5xD(197)(3) <= VNStageIntLLROutputS4xD(192)(3);
  CNStageIntLLRInputS5xD(243)(3) <= VNStageIntLLROutputS4xD(192)(4);
  CNStageIntLLRInputS5xD(297)(3) <= VNStageIntLLROutputS4xD(192)(5);
  CNStageIntLLRInputS5xD(340)(3) <= VNStageIntLLROutputS4xD(192)(6);
  CNStageIntLLRInputS5xD(51)(3) <= VNStageIntLLROutputS4xD(193)(0);
  CNStageIntLLRInputS5xD(58)(3) <= VNStageIntLLROutputS4xD(193)(1);
  CNStageIntLLRInputS5xD(137)(3) <= VNStageIntLLROutputS4xD(193)(2);
  CNStageIntLLRInputS5xD(269)(3) <= VNStageIntLLROutputS4xD(193)(3);
  CNStageIntLLRInputS5xD(333)(3) <= VNStageIntLLROutputS4xD(193)(4);
  CNStageIntLLRInputS5xD(50)(3) <= VNStageIntLLROutputS4xD(194)(0);
  CNStageIntLLRInputS5xD(55)(3) <= VNStageIntLLROutputS4xD(194)(1);
  CNStageIntLLRInputS5xD(115)(3) <= VNStageIntLLROutputS4xD(194)(2);
  CNStageIntLLRInputS5xD(171)(3) <= VNStageIntLLROutputS4xD(194)(3);
  CNStageIntLLRInputS5xD(275)(3) <= VNStageIntLLROutputS4xD(194)(4);
  CNStageIntLLRInputS5xD(304)(3) <= VNStageIntLLROutputS4xD(194)(5);
  CNStageIntLLRInputS5xD(371)(3) <= VNStageIntLLROutputS4xD(194)(6);
  CNStageIntLLRInputS5xD(72)(3) <= VNStageIntLLROutputS4xD(195)(0);
  CNStageIntLLRInputS5xD(139)(3) <= VNStageIntLLROutputS4xD(195)(1);
  CNStageIntLLRInputS5xD(187)(3) <= VNStageIntLLROutputS4xD(195)(2);
  CNStageIntLLRInputS5xD(244)(3) <= VNStageIntLLROutputS4xD(195)(3);
  CNStageIntLLRInputS5xD(49)(3) <= VNStageIntLLROutputS4xD(196)(0);
  CNStageIntLLRInputS5xD(64)(3) <= VNStageIntLLROutputS4xD(196)(1);
  CNStageIntLLRInputS5xD(153)(3) <= VNStageIntLLROutputS4xD(196)(2);
  CNStageIntLLRInputS5xD(205)(3) <= VNStageIntLLROutputS4xD(196)(3);
  CNStageIntLLRInputS5xD(242)(3) <= VNStageIntLLROutputS4xD(196)(4);
  CNStageIntLLRInputS5xD(306)(3) <= VNStageIntLLROutputS4xD(196)(5);
  CNStageIntLLRInputS5xD(48)(3) <= VNStageIntLLROutputS4xD(197)(0);
  CNStageIntLLRInputS5xD(96)(3) <= VNStageIntLLROutputS4xD(197)(1);
  CNStageIntLLRInputS5xD(150)(3) <= VNStageIntLLROutputS4xD(197)(2);
  CNStageIntLLRInputS5xD(213)(3) <= VNStageIntLLROutputS4xD(197)(3);
  CNStageIntLLRInputS5xD(273)(3) <= VNStageIntLLROutputS4xD(197)(4);
  CNStageIntLLRInputS5xD(320)(3) <= VNStageIntLLROutputS4xD(197)(5);
  CNStageIntLLRInputS5xD(363)(3) <= VNStageIntLLROutputS4xD(197)(6);
  CNStageIntLLRInputS5xD(47)(3) <= VNStageIntLLROutputS4xD(198)(0);
  CNStageIntLLRInputS5xD(105)(3) <= VNStageIntLLROutputS4xD(198)(1);
  CNStageIntLLRInputS5xD(111)(3) <= VNStageIntLLROutputS4xD(198)(2);
  CNStageIntLLRInputS5xD(208)(3) <= VNStageIntLLROutputS4xD(198)(3);
  CNStageIntLLRInputS5xD(254)(3) <= VNStageIntLLROutputS4xD(198)(4);
  CNStageIntLLRInputS5xD(316)(3) <= VNStageIntLLROutputS4xD(198)(5);
  CNStageIntLLRInputS5xD(379)(3) <= VNStageIntLLROutputS4xD(198)(6);
  CNStageIntLLRInputS5xD(46)(3) <= VNStageIntLLROutputS4xD(199)(0);
  CNStageIntLLRInputS5xD(99)(3) <= VNStageIntLLROutputS4xD(199)(1);
  CNStageIntLLRInputS5xD(133)(3) <= VNStageIntLLROutputS4xD(199)(2);
  CNStageIntLLRInputS5xD(214)(3) <= VNStageIntLLROutputS4xD(199)(3);
  CNStageIntLLRInputS5xD(257)(3) <= VNStageIntLLROutputS4xD(199)(4);
  CNStageIntLLRInputS5xD(282)(3) <= VNStageIntLLROutputS4xD(199)(5);
  CNStageIntLLRInputS5xD(350)(3) <= VNStageIntLLROutputS4xD(199)(6);
  CNStageIntLLRInputS5xD(45)(3) <= VNStageIntLLROutputS4xD(200)(0);
  CNStageIntLLRInputS5xD(102)(3) <= VNStageIntLLROutputS4xD(200)(1);
  CNStageIntLLRInputS5xD(134)(3) <= VNStageIntLLROutputS4xD(200)(2);
  CNStageIntLLRInputS5xD(204)(3) <= VNStageIntLLROutputS4xD(200)(3);
  CNStageIntLLRInputS5xD(245)(3) <= VNStageIntLLROutputS4xD(200)(4);
  CNStageIntLLRInputS5xD(300)(3) <= VNStageIntLLROutputS4xD(200)(5);
  CNStageIntLLRInputS5xD(44)(3) <= VNStageIntLLROutputS4xD(201)(0);
  CNStageIntLLRInputS5xD(93)(3) <= VNStageIntLLROutputS4xD(201)(1);
  CNStageIntLLRInputS5xD(169)(3) <= VNStageIntLLROutputS4xD(201)(2);
  CNStageIntLLRInputS5xD(174)(3) <= VNStageIntLLROutputS4xD(201)(3);
  CNStageIntLLRInputS5xD(274)(3) <= VNStageIntLLROutputS4xD(201)(4);
  CNStageIntLLRInputS5xD(351)(3) <= VNStageIntLLROutputS4xD(201)(5);
  CNStageIntLLRInputS5xD(43)(3) <= VNStageIntLLROutputS4xD(202)(0);
  CNStageIntLLRInputS5xD(73)(3) <= VNStageIntLLROutputS4xD(202)(1);
  CNStageIntLLRInputS5xD(160)(3) <= VNStageIntLLROutputS4xD(202)(2);
  CNStageIntLLRInputS5xD(181)(3) <= VNStageIntLLROutputS4xD(202)(3);
  CNStageIntLLRInputS5xD(281)(3) <= VNStageIntLLROutputS4xD(202)(4);
  CNStageIntLLRInputS5xD(365)(3) <= VNStageIntLLROutputS4xD(202)(5);
  CNStageIntLLRInputS5xD(42)(3) <= VNStageIntLLROutputS4xD(203)(0);
  CNStageIntLLRInputS5xD(54)(3) <= VNStageIntLLROutputS4xD(203)(1);
  CNStageIntLLRInputS5xD(119)(3) <= VNStageIntLLROutputS4xD(203)(2);
  CNStageIntLLRInputS5xD(217)(3) <= VNStageIntLLROutputS4xD(203)(3);
  CNStageIntLLRInputS5xD(267)(3) <= VNStageIntLLROutputS4xD(203)(4);
  CNStageIntLLRInputS5xD(326)(3) <= VNStageIntLLROutputS4xD(203)(5);
  CNStageIntLLRInputS5xD(361)(3) <= VNStageIntLLROutputS4xD(203)(6);
  CNStageIntLLRInputS5xD(41)(3) <= VNStageIntLLROutputS4xD(204)(0);
  CNStageIntLLRInputS5xD(68)(3) <= VNStageIntLLROutputS4xD(204)(1);
  CNStageIntLLRInputS5xD(123)(3) <= VNStageIntLLROutputS4xD(204)(2);
  CNStageIntLLRInputS5xD(219)(3) <= VNStageIntLLROutputS4xD(204)(3);
  CNStageIntLLRInputS5xD(251)(3) <= VNStageIntLLROutputS4xD(204)(4);
  CNStageIntLLRInputS5xD(288)(3) <= VNStageIntLLROutputS4xD(204)(5);
  CNStageIntLLRInputS5xD(382)(3) <= VNStageIntLLROutputS4xD(204)(6);
  CNStageIntLLRInputS5xD(170)(3) <= VNStageIntLLROutputS4xD(205)(0);
  CNStageIntLLRInputS5xD(276)(3) <= VNStageIntLLROutputS4xD(205)(1);
  CNStageIntLLRInputS5xD(345)(3) <= VNStageIntLLROutputS4xD(205)(2);
  CNStageIntLLRInputS5xD(40)(3) <= VNStageIntLLROutputS4xD(206)(0);
  CNStageIntLLRInputS5xD(122)(3) <= VNStageIntLLROutputS4xD(206)(1);
  CNStageIntLLRInputS5xD(172)(3) <= VNStageIntLLROutputS4xD(206)(2);
  CNStageIntLLRInputS5xD(332)(3) <= VNStageIntLLROutputS4xD(206)(3);
  CNStageIntLLRInputS5xD(346)(3) <= VNStageIntLLROutputS4xD(206)(4);
  CNStageIntLLRInputS5xD(39)(3) <= VNStageIntLLROutputS4xD(207)(0);
  CNStageIntLLRInputS5xD(95)(3) <= VNStageIntLLROutputS4xD(207)(1);
  CNStageIntLLRInputS5xD(117)(3) <= VNStageIntLLROutputS4xD(207)(2);
  CNStageIntLLRInputS5xD(255)(3) <= VNStageIntLLROutputS4xD(207)(3);
  CNStageIntLLRInputS5xD(292)(3) <= VNStageIntLLROutputS4xD(207)(4);
  CNStageIntLLRInputS5xD(381)(3) <= VNStageIntLLROutputS4xD(207)(5);
  CNStageIntLLRInputS5xD(38)(3) <= VNStageIntLLROutputS4xD(208)(0);
  CNStageIntLLRInputS5xD(82)(3) <= VNStageIntLLROutputS4xD(208)(1);
  CNStageIntLLRInputS5xD(157)(3) <= VNStageIntLLROutputS4xD(208)(2);
  CNStageIntLLRInputS5xD(191)(3) <= VNStageIntLLROutputS4xD(208)(3);
  CNStageIntLLRInputS5xD(286)(3) <= VNStageIntLLROutputS4xD(208)(4);
  CNStageIntLLRInputS5xD(372)(3) <= VNStageIntLLROutputS4xD(208)(5);
  CNStageIntLLRInputS5xD(37)(3) <= VNStageIntLLROutputS4xD(209)(0);
  CNStageIntLLRInputS5xD(97)(3) <= VNStageIntLLROutputS4xD(209)(1);
  CNStageIntLLRInputS5xD(165)(3) <= VNStageIntLLROutputS4xD(209)(2);
  CNStageIntLLRInputS5xD(218)(3) <= VNStageIntLLROutputS4xD(209)(3);
  CNStageIntLLRInputS5xD(323)(3) <= VNStageIntLLROutputS4xD(209)(4);
  CNStageIntLLRInputS5xD(36)(3) <= VNStageIntLLROutputS4xD(210)(0);
  CNStageIntLLRInputS5xD(60)(3) <= VNStageIntLLROutputS4xD(210)(1);
  CNStageIntLLRInputS5xD(129)(3) <= VNStageIntLLROutputS4xD(210)(2);
  CNStageIntLLRInputS5xD(180)(3) <= VNStageIntLLROutputS4xD(210)(3);
  CNStageIntLLRInputS5xD(246)(3) <= VNStageIntLLROutputS4xD(210)(4);
  CNStageIntLLRInputS5xD(330)(3) <= VNStageIntLLROutputS4xD(210)(5);
  CNStageIntLLRInputS5xD(335)(3) <= VNStageIntLLROutputS4xD(210)(6);
  CNStageIntLLRInputS5xD(35)(3) <= VNStageIntLLROutputS4xD(211)(0);
  CNStageIntLLRInputS5xD(70)(3) <= VNStageIntLLROutputS4xD(211)(1);
  CNStageIntLLRInputS5xD(127)(3) <= VNStageIntLLROutputS4xD(211)(2);
  CNStageIntLLRInputS5xD(206)(3) <= VNStageIntLLROutputS4xD(211)(3);
  CNStageIntLLRInputS5xD(260)(3) <= VNStageIntLLROutputS4xD(211)(4);
  CNStageIntLLRInputS5xD(298)(3) <= VNStageIntLLROutputS4xD(211)(5);
  CNStageIntLLRInputS5xD(34)(3) <= VNStageIntLLROutputS4xD(212)(0);
  CNStageIntLLRInputS5xD(65)(3) <= VNStageIntLLROutputS4xD(212)(1);
  CNStageIntLLRInputS5xD(163)(3) <= VNStageIntLLROutputS4xD(212)(2);
  CNStageIntLLRInputS5xD(186)(3) <= VNStageIntLLROutputS4xD(212)(3);
  CNStageIntLLRInputS5xD(296)(3) <= VNStageIntLLROutputS4xD(212)(4);
  CNStageIntLLRInputS5xD(33)(3) <= VNStageIntLLROutputS4xD(213)(0);
  CNStageIntLLRInputS5xD(71)(3) <= VNStageIntLLROutputS4xD(213)(1);
  CNStageIntLLRInputS5xD(142)(3) <= VNStageIntLLROutputS4xD(213)(2);
  CNStageIntLLRInputS5xD(230)(3) <= VNStageIntLLROutputS4xD(213)(3);
  CNStageIntLLRInputS5xD(32)(3) <= VNStageIntLLROutputS4xD(214)(0);
  CNStageIntLLRInputS5xD(59)(3) <= VNStageIntLLROutputS4xD(214)(1);
  CNStageIntLLRInputS5xD(145)(3) <= VNStageIntLLROutputS4xD(214)(2);
  CNStageIntLLRInputS5xD(220)(3) <= VNStageIntLLROutputS4xD(214)(3);
  CNStageIntLLRInputS5xD(240)(3) <= VNStageIntLLROutputS4xD(214)(4);
  CNStageIntLLRInputS5xD(308)(3) <= VNStageIntLLROutputS4xD(214)(5);
  CNStageIntLLRInputS5xD(369)(3) <= VNStageIntLLROutputS4xD(214)(6);
  CNStageIntLLRInputS5xD(31)(3) <= VNStageIntLLROutputS4xD(215)(0);
  CNStageIntLLRInputS5xD(85)(3) <= VNStageIntLLROutputS4xD(215)(1);
  CNStageIntLLRInputS5xD(130)(3) <= VNStageIntLLROutputS4xD(215)(2);
  CNStageIntLLRInputS5xD(216)(3) <= VNStageIntLLROutputS4xD(215)(3);
  CNStageIntLLRInputS5xD(234)(3) <= VNStageIntLLROutputS4xD(215)(4);
  CNStageIntLLRInputS5xD(311)(3) <= VNStageIntLLROutputS4xD(215)(5);
  CNStageIntLLRInputS5xD(377)(3) <= VNStageIntLLROutputS4xD(215)(6);
  CNStageIntLLRInputS5xD(30)(3) <= VNStageIntLLROutputS4xD(216)(0);
  CNStageIntLLRInputS5xD(91)(3) <= VNStageIntLLROutputS4xD(216)(1);
  CNStageIntLLRInputS5xD(164)(3) <= VNStageIntLLROutputS4xD(216)(2);
  CNStageIntLLRInputS5xD(183)(3) <= VNStageIntLLROutputS4xD(216)(3);
  CNStageIntLLRInputS5xD(237)(3) <= VNStageIntLLROutputS4xD(216)(4);
  CNStageIntLLRInputS5xD(299)(3) <= VNStageIntLLROutputS4xD(216)(5);
  CNStageIntLLRInputS5xD(341)(3) <= VNStageIntLLROutputS4xD(216)(6);
  CNStageIntLLRInputS5xD(29)(3) <= VNStageIntLLROutputS4xD(217)(0);
  CNStageIntLLRInputS5xD(75)(3) <= VNStageIntLLROutputS4xD(217)(1);
  CNStageIntLLRInputS5xD(126)(3) <= VNStageIntLLROutputS4xD(217)(2);
  CNStageIntLLRInputS5xD(201)(3) <= VNStageIntLLROutputS4xD(217)(3);
  CNStageIntLLRInputS5xD(227)(3) <= VNStageIntLLROutputS4xD(217)(4);
  CNStageIntLLRInputS5xD(329)(3) <= VNStageIntLLROutputS4xD(217)(5);
  CNStageIntLLRInputS5xD(339)(3) <= VNStageIntLLROutputS4xD(217)(6);
  CNStageIntLLRInputS5xD(28)(3) <= VNStageIntLLROutputS4xD(218)(0);
  CNStageIntLLRInputS5xD(77)(3) <= VNStageIntLLROutputS4xD(218)(1);
  CNStageIntLLRInputS5xD(154)(3) <= VNStageIntLLROutputS4xD(218)(2);
  CNStageIntLLRInputS5xD(202)(3) <= VNStageIntLLROutputS4xD(218)(3);
  CNStageIntLLRInputS5xD(261)(3) <= VNStageIntLLROutputS4xD(218)(4);
  CNStageIntLLRInputS5xD(295)(3) <= VNStageIntLLROutputS4xD(218)(5);
  CNStageIntLLRInputS5xD(375)(3) <= VNStageIntLLROutputS4xD(218)(6);
  CNStageIntLLRInputS5xD(27)(3) <= VNStageIntLLROutputS4xD(219)(0);
  CNStageIntLLRInputS5xD(101)(3) <= VNStageIntLLROutputS4xD(219)(1);
  CNStageIntLLRInputS5xD(138)(3) <= VNStageIntLLROutputS4xD(219)(2);
  CNStageIntLLRInputS5xD(182)(3) <= VNStageIntLLROutputS4xD(219)(3);
  CNStageIntLLRInputS5xD(321)(3) <= VNStageIntLLROutputS4xD(219)(4);
  CNStageIntLLRInputS5xD(354)(3) <= VNStageIntLLROutputS4xD(219)(5);
  CNStageIntLLRInputS5xD(26)(3) <= VNStageIntLLROutputS4xD(220)(0);
  CNStageIntLLRInputS5xD(83)(3) <= VNStageIntLLROutputS4xD(220)(1);
  CNStageIntLLRInputS5xD(166)(3) <= VNStageIntLLROutputS4xD(220)(2);
  CNStageIntLLRInputS5xD(173)(3) <= VNStageIntLLROutputS4xD(220)(3);
  CNStageIntLLRInputS5xD(256)(3) <= VNStageIntLLROutputS4xD(220)(4);
  CNStageIntLLRInputS5xD(305)(3) <= VNStageIntLLROutputS4xD(220)(5);
  CNStageIntLLRInputS5xD(356)(3) <= VNStageIntLLROutputS4xD(220)(6);
  CNStageIntLLRInputS5xD(25)(3) <= VNStageIntLLROutputS4xD(221)(0);
  CNStageIntLLRInputS5xD(94)(3) <= VNStageIntLLROutputS4xD(221)(1);
  CNStageIntLLRInputS5xD(156)(3) <= VNStageIntLLROutputS4xD(221)(2);
  CNStageIntLLRInputS5xD(190)(3) <= VNStageIntLLROutputS4xD(221)(3);
  CNStageIntLLRInputS5xD(268)(3) <= VNStageIntLLROutputS4xD(221)(4);
  CNStageIntLLRInputS5xD(331)(3) <= VNStageIntLLROutputS4xD(221)(5);
  CNStageIntLLRInputS5xD(342)(3) <= VNStageIntLLROutputS4xD(221)(6);
  CNStageIntLLRInputS5xD(24)(3) <= VNStageIntLLROutputS4xD(222)(0);
  CNStageIntLLRInputS5xD(143)(3) <= VNStageIntLLROutputS4xD(222)(1);
  CNStageIntLLRInputS5xD(241)(3) <= VNStageIntLLROutputS4xD(222)(2);
  CNStageIntLLRInputS5xD(376)(3) <= VNStageIntLLROutputS4xD(222)(3);
  CNStageIntLLRInputS5xD(23)(3) <= VNStageIntLLROutputS4xD(223)(0);
  CNStageIntLLRInputS5xD(76)(3) <= VNStageIntLLROutputS4xD(223)(1);
  CNStageIntLLRInputS5xD(162)(3) <= VNStageIntLLROutputS4xD(223)(2);
  CNStageIntLLRInputS5xD(224)(3) <= VNStageIntLLROutputS4xD(223)(3);
  CNStageIntLLRInputS5xD(229)(3) <= VNStageIntLLROutputS4xD(223)(4);
  CNStageIntLLRInputS5xD(309)(3) <= VNStageIntLLROutputS4xD(223)(5);
  CNStageIntLLRInputS5xD(338)(3) <= VNStageIntLLROutputS4xD(223)(6);
  CNStageIntLLRInputS5xD(22)(3) <= VNStageIntLLROutputS4xD(224)(0);
  CNStageIntLLRInputS5xD(90)(3) <= VNStageIntLLROutputS4xD(224)(1);
  CNStageIntLLRInputS5xD(135)(3) <= VNStageIntLLROutputS4xD(224)(2);
  CNStageIntLLRInputS5xD(193)(3) <= VNStageIntLLROutputS4xD(224)(3);
  CNStageIntLLRInputS5xD(270)(3) <= VNStageIntLLROutputS4xD(224)(4);
  CNStageIntLLRInputS5xD(328)(3) <= VNStageIntLLROutputS4xD(224)(5);
  CNStageIntLLRInputS5xD(366)(3) <= VNStageIntLLROutputS4xD(224)(6);
  CNStageIntLLRInputS5xD(21)(3) <= VNStageIntLLROutputS4xD(225)(0);
  CNStageIntLLRInputS5xD(61)(3) <= VNStageIntLLROutputS4xD(225)(1);
  CNStageIntLLRInputS5xD(132)(3) <= VNStageIntLLROutputS4xD(225)(2);
  CNStageIntLLRInputS5xD(188)(3) <= VNStageIntLLROutputS4xD(225)(3);
  CNStageIntLLRInputS5xD(232)(3) <= VNStageIntLLROutputS4xD(225)(4);
  CNStageIntLLRInputS5xD(301)(3) <= VNStageIntLLROutputS4xD(225)(5);
  CNStageIntLLRInputS5xD(20)(3) <= VNStageIntLLROutputS4xD(226)(0);
  CNStageIntLLRInputS5xD(148)(3) <= VNStageIntLLROutputS4xD(226)(1);
  CNStageIntLLRInputS5xD(378)(3) <= VNStageIntLLROutputS4xD(226)(2);
  CNStageIntLLRInputS5xD(19)(3) <= VNStageIntLLROutputS4xD(227)(0);
  CNStageIntLLRInputS5xD(63)(3) <= VNStageIntLLROutputS4xD(227)(1);
  CNStageIntLLRInputS5xD(140)(3) <= VNStageIntLLROutputS4xD(227)(2);
  CNStageIntLLRInputS5xD(178)(3) <= VNStageIntLLROutputS4xD(227)(3);
  CNStageIntLLRInputS5xD(258)(3) <= VNStageIntLLROutputS4xD(227)(4);
  CNStageIntLLRInputS5xD(314)(3) <= VNStageIntLLROutputS4xD(227)(5);
  CNStageIntLLRInputS5xD(368)(3) <= VNStageIntLLROutputS4xD(227)(6);
  CNStageIntLLRInputS5xD(18)(3) <= VNStageIntLLROutputS4xD(228)(0);
  CNStageIntLLRInputS5xD(78)(3) <= VNStageIntLLROutputS4xD(228)(1);
  CNStageIntLLRInputS5xD(114)(3) <= VNStageIntLLROutputS4xD(228)(2);
  CNStageIntLLRInputS5xD(198)(3) <= VNStageIntLLROutputS4xD(228)(3);
  CNStageIntLLRInputS5xD(253)(3) <= VNStageIntLLROutputS4xD(228)(4);
  CNStageIntLLRInputS5xD(307)(3) <= VNStageIntLLROutputS4xD(228)(5);
  CNStageIntLLRInputS5xD(17)(3) <= VNStageIntLLROutputS4xD(229)(0);
  CNStageIntLLRInputS5xD(74)(3) <= VNStageIntLLROutputS4xD(229)(1);
  CNStageIntLLRInputS5xD(124)(3) <= VNStageIntLLROutputS4xD(229)(2);
  CNStageIntLLRInputS5xD(259)(3) <= VNStageIntLLROutputS4xD(229)(3);
  CNStageIntLLRInputS5xD(374)(3) <= VNStageIntLLROutputS4xD(229)(4);
  CNStageIntLLRInputS5xD(16)(3) <= VNStageIntLLROutputS4xD(230)(0);
  CNStageIntLLRInputS5xD(118)(3) <= VNStageIntLLROutputS4xD(230)(1);
  CNStageIntLLRInputS5xD(176)(3) <= VNStageIntLLROutputS4xD(230)(2);
  CNStageIntLLRInputS5xD(249)(3) <= VNStageIntLLROutputS4xD(230)(3);
  CNStageIntLLRInputS5xD(293)(3) <= VNStageIntLLROutputS4xD(230)(4);
  CNStageIntLLRInputS5xD(347)(3) <= VNStageIntLLROutputS4xD(230)(5);
  CNStageIntLLRInputS5xD(15)(3) <= VNStageIntLLROutputS4xD(231)(0);
  CNStageIntLLRInputS5xD(56)(3) <= VNStageIntLLROutputS4xD(231)(1);
  CNStageIntLLRInputS5xD(209)(3) <= VNStageIntLLROutputS4xD(231)(2);
  CNStageIntLLRInputS5xD(272)(3) <= VNStageIntLLROutputS4xD(231)(3);
  CNStageIntLLRInputS5xD(287)(3) <= VNStageIntLLROutputS4xD(231)(4);
  CNStageIntLLRInputS5xD(344)(3) <= VNStageIntLLROutputS4xD(231)(5);
  CNStageIntLLRInputS5xD(14)(3) <= VNStageIntLLROutputS4xD(232)(0);
  CNStageIntLLRInputS5xD(57)(3) <= VNStageIntLLROutputS4xD(232)(1);
  CNStageIntLLRInputS5xD(212)(3) <= VNStageIntLLROutputS4xD(232)(2);
  CNStageIntLLRInputS5xD(278)(3) <= VNStageIntLLROutputS4xD(232)(3);
  CNStageIntLLRInputS5xD(291)(3) <= VNStageIntLLROutputS4xD(232)(4);
  CNStageIntLLRInputS5xD(359)(3) <= VNStageIntLLROutputS4xD(232)(5);
  CNStageIntLLRInputS5xD(13)(3) <= VNStageIntLLROutputS4xD(233)(0);
  CNStageIntLLRInputS5xD(92)(3) <= VNStageIntLLROutputS4xD(233)(1);
  CNStageIntLLRInputS5xD(149)(3) <= VNStageIntLLROutputS4xD(233)(2);
  CNStageIntLLRInputS5xD(263)(3) <= VNStageIntLLROutputS4xD(233)(3);
  CNStageIntLLRInputS5xD(352)(3) <= VNStageIntLLROutputS4xD(233)(4);
  CNStageIntLLRInputS5xD(12)(3) <= VNStageIntLLROutputS4xD(234)(0);
  CNStageIntLLRInputS5xD(84)(3) <= VNStageIntLLROutputS4xD(234)(1);
  CNStageIntLLRInputS5xD(131)(3) <= VNStageIntLLROutputS4xD(234)(2);
  CNStageIntLLRInputS5xD(177)(3) <= VNStageIntLLROutputS4xD(234)(3);
  CNStageIntLLRInputS5xD(265)(3) <= VNStageIntLLROutputS4xD(234)(4);
  CNStageIntLLRInputS5xD(315)(3) <= VNStageIntLLROutputS4xD(234)(5);
  CNStageIntLLRInputS5xD(100)(3) <= VNStageIntLLROutputS4xD(235)(0);
  CNStageIntLLRInputS5xD(144)(3) <= VNStageIntLLROutputS4xD(235)(1);
  CNStageIntLLRInputS5xD(196)(3) <= VNStageIntLLROutputS4xD(235)(2);
  CNStageIntLLRInputS5xD(235)(3) <= VNStageIntLLROutputS4xD(235)(3);
  CNStageIntLLRInputS5xD(336)(3) <= VNStageIntLLROutputS4xD(235)(4);
  CNStageIntLLRInputS5xD(11)(3) <= VNStageIntLLROutputS4xD(236)(0);
  CNStageIntLLRInputS5xD(104)(3) <= VNStageIntLLROutputS4xD(236)(1);
  CNStageIntLLRInputS5xD(155)(3) <= VNStageIntLLROutputS4xD(236)(2);
  CNStageIntLLRInputS5xD(221)(3) <= VNStageIntLLROutputS4xD(236)(3);
  CNStageIntLLRInputS5xD(271)(3) <= VNStageIntLLROutputS4xD(236)(4);
  CNStageIntLLRInputS5xD(310)(3) <= VNStageIntLLROutputS4xD(236)(5);
  CNStageIntLLRInputS5xD(10)(3) <= VNStageIntLLROutputS4xD(237)(0);
  CNStageIntLLRInputS5xD(110)(3) <= VNStageIntLLROutputS4xD(237)(1);
  CNStageIntLLRInputS5xD(125)(3) <= VNStageIntLLROutputS4xD(237)(2);
  CNStageIntLLRInputS5xD(228)(3) <= VNStageIntLLROutputS4xD(237)(3);
  CNStageIntLLRInputS5xD(322)(3) <= VNStageIntLLROutputS4xD(237)(4);
  CNStageIntLLRInputS5xD(334)(3) <= VNStageIntLLROutputS4xD(237)(5);
  CNStageIntLLRInputS5xD(9)(3) <= VNStageIntLLROutputS4xD(238)(0);
  CNStageIntLLRInputS5xD(103)(3) <= VNStageIntLLROutputS4xD(238)(1);
  CNStageIntLLRInputS5xD(113)(3) <= VNStageIntLLROutputS4xD(238)(2);
  CNStageIntLLRInputS5xD(179)(3) <= VNStageIntLLROutputS4xD(238)(3);
  CNStageIntLLRInputS5xD(236)(3) <= VNStageIntLLROutputS4xD(238)(4);
  CNStageIntLLRInputS5xD(294)(3) <= VNStageIntLLROutputS4xD(238)(5);
  CNStageIntLLRInputS5xD(383)(3) <= VNStageIntLLROutputS4xD(238)(6);
  CNStageIntLLRInputS5xD(8)(3) <= VNStageIntLLROutputS4xD(239)(0);
  CNStageIntLLRInputS5xD(98)(3) <= VNStageIntLLROutputS4xD(239)(1);
  CNStageIntLLRInputS5xD(158)(3) <= VNStageIntLLROutputS4xD(239)(2);
  CNStageIntLLRInputS5xD(223)(3) <= VNStageIntLLROutputS4xD(239)(3);
  CNStageIntLLRInputS5xD(264)(3) <= VNStageIntLLROutputS4xD(239)(4);
  CNStageIntLLRInputS5xD(284)(3) <= VNStageIntLLROutputS4xD(239)(5);
  CNStageIntLLRInputS5xD(360)(3) <= VNStageIntLLROutputS4xD(239)(6);
  CNStageIntLLRInputS5xD(7)(3) <= VNStageIntLLROutputS4xD(240)(0);
  CNStageIntLLRInputS5xD(81)(3) <= VNStageIntLLROutputS4xD(240)(1);
  CNStageIntLLRInputS5xD(116)(3) <= VNStageIntLLROutputS4xD(240)(2);
  CNStageIntLLRInputS5xD(210)(3) <= VNStageIntLLROutputS4xD(240)(3);
  CNStageIntLLRInputS5xD(277)(3) <= VNStageIntLLROutputS4xD(240)(4);
  CNStageIntLLRInputS5xD(324)(3) <= VNStageIntLLROutputS4xD(240)(5);
  CNStageIntLLRInputS5xD(343)(3) <= VNStageIntLLROutputS4xD(240)(6);
  CNStageIntLLRInputS5xD(6)(3) <= VNStageIntLLROutputS4xD(241)(0);
  CNStageIntLLRInputS5xD(88)(3) <= VNStageIntLLROutputS4xD(241)(1);
  CNStageIntLLRInputS5xD(175)(3) <= VNStageIntLLROutputS4xD(241)(2);
  CNStageIntLLRInputS5xD(250)(3) <= VNStageIntLLROutputS4xD(241)(3);
  CNStageIntLLRInputS5xD(285)(3) <= VNStageIntLLROutputS4xD(241)(4);
  CNStageIntLLRInputS5xD(355)(3) <= VNStageIntLLROutputS4xD(241)(5);
  CNStageIntLLRInputS5xD(5)(3) <= VNStageIntLLROutputS4xD(242)(0);
  CNStageIntLLRInputS5xD(108)(3) <= VNStageIntLLROutputS4xD(242)(1);
  CNStageIntLLRInputS5xD(146)(3) <= VNStageIntLLROutputS4xD(242)(2);
  CNStageIntLLRInputS5xD(203)(3) <= VNStageIntLLROutputS4xD(242)(3);
  CNStageIntLLRInputS5xD(231)(3) <= VNStageIntLLROutputS4xD(242)(4);
  CNStageIntLLRInputS5xD(303)(3) <= VNStageIntLLROutputS4xD(242)(5);
  CNStageIntLLRInputS5xD(367)(3) <= VNStageIntLLROutputS4xD(242)(6);
  CNStageIntLLRInputS5xD(4)(3) <= VNStageIntLLROutputS4xD(243)(0);
  CNStageIntLLRInputS5xD(106)(3) <= VNStageIntLLROutputS4xD(243)(1);
  CNStageIntLLRInputS5xD(141)(3) <= VNStageIntLLROutputS4xD(243)(2);
  CNStageIntLLRInputS5xD(200)(3) <= VNStageIntLLROutputS4xD(243)(3);
  CNStageIntLLRInputS5xD(252)(3) <= VNStageIntLLROutputS4xD(243)(4);
  CNStageIntLLRInputS5xD(312)(3) <= VNStageIntLLROutputS4xD(243)(5);
  CNStageIntLLRInputS5xD(337)(3) <= VNStageIntLLROutputS4xD(243)(6);
  CNStageIntLLRInputS5xD(147)(3) <= VNStageIntLLROutputS4xD(244)(0);
  CNStageIntLLRInputS5xD(266)(3) <= VNStageIntLLROutputS4xD(244)(1);
  CNStageIntLLRInputS5xD(3)(3) <= VNStageIntLLROutputS4xD(245)(0);
  CNStageIntLLRInputS5xD(66)(3) <= VNStageIntLLROutputS4xD(245)(1);
  CNStageIntLLRInputS5xD(136)(3) <= VNStageIntLLROutputS4xD(245)(2);
  CNStageIntLLRInputS5xD(207)(3) <= VNStageIntLLROutputS4xD(245)(3);
  CNStageIntLLRInputS5xD(262)(3) <= VNStageIntLLROutputS4xD(245)(4);
  CNStageIntLLRInputS5xD(313)(3) <= VNStageIntLLROutputS4xD(245)(5);
  CNStageIntLLRInputS5xD(370)(3) <= VNStageIntLLROutputS4xD(245)(6);
  CNStageIntLLRInputS5xD(2)(3) <= VNStageIntLLROutputS4xD(246)(0);
  CNStageIntLLRInputS5xD(69)(3) <= VNStageIntLLROutputS4xD(246)(1);
  CNStageIntLLRInputS5xD(161)(3) <= VNStageIntLLROutputS4xD(246)(2);
  CNStageIntLLRInputS5xD(185)(3) <= VNStageIntLLROutputS4xD(246)(3);
  CNStageIntLLRInputS5xD(226)(3) <= VNStageIntLLROutputS4xD(246)(4);
  CNStageIntLLRInputS5xD(302)(3) <= VNStageIntLLROutputS4xD(246)(5);
  CNStageIntLLRInputS5xD(1)(3) <= VNStageIntLLROutputS4xD(247)(0);
  CNStageIntLLRInputS5xD(109)(3) <= VNStageIntLLROutputS4xD(247)(1);
  CNStageIntLLRInputS5xD(168)(3) <= VNStageIntLLROutputS4xD(247)(2);
  CNStageIntLLRInputS5xD(194)(3) <= VNStageIntLLROutputS4xD(247)(3);
  CNStageIntLLRInputS5xD(247)(3) <= VNStageIntLLROutputS4xD(247)(4);
  CNStageIntLLRInputS5xD(327)(3) <= VNStageIntLLROutputS4xD(247)(5);
  CNStageIntLLRInputS5xD(349)(3) <= VNStageIntLLROutputS4xD(247)(6);
  CNStageIntLLRInputS5xD(0)(3) <= VNStageIntLLROutputS4xD(248)(0);
  CNStageIntLLRInputS5xD(87)(3) <= VNStageIntLLROutputS4xD(248)(1);
  CNStageIntLLRInputS5xD(151)(3) <= VNStageIntLLROutputS4xD(248)(2);
  CNStageIntLLRInputS5xD(189)(3) <= VNStageIntLLROutputS4xD(248)(3);
  CNStageIntLLRInputS5xD(248)(3) <= VNStageIntLLROutputS4xD(248)(4);
  CNStageIntLLRInputS5xD(280)(3) <= VNStageIntLLROutputS4xD(248)(5);
  CNStageIntLLRInputS5xD(357)(3) <= VNStageIntLLROutputS4xD(248)(6);
  CNStageIntLLRInputS5xD(152)(3) <= VNStageIntLLROutputS4xD(249)(0);
  CNStageIntLLRInputS5xD(192)(3) <= VNStageIntLLROutputS4xD(249)(1);
  CNStageIntLLRInputS5xD(225)(3) <= VNStageIntLLROutputS4xD(249)(2);
  CNStageIntLLRInputS5xD(317)(3) <= VNStageIntLLROutputS4xD(249)(3);
  CNStageIntLLRInputS5xD(353)(3) <= VNStageIntLLROutputS4xD(249)(4);
  CNStageIntLLRInputS5xD(79)(3) <= VNStageIntLLROutputS4xD(250)(0);
  CNStageIntLLRInputS5xD(120)(3) <= VNStageIntLLROutputS4xD(250)(1);
  CNStageIntLLRInputS5xD(184)(3) <= VNStageIntLLROutputS4xD(250)(2);
  CNStageIntLLRInputS5xD(319)(3) <= VNStageIntLLROutputS4xD(250)(3);
  CNStageIntLLRInputS5xD(358)(3) <= VNStageIntLLROutputS4xD(250)(4);
  CNStageIntLLRInputS5xD(62)(3) <= VNStageIntLLROutputS4xD(251)(0);
  CNStageIntLLRInputS5xD(159)(3) <= VNStageIntLLROutputS4xD(251)(1);
  CNStageIntLLRInputS5xD(215)(3) <= VNStageIntLLROutputS4xD(251)(2);
  CNStageIntLLRInputS5xD(289)(3) <= VNStageIntLLROutputS4xD(251)(3);
  CNStageIntLLRInputS5xD(348)(3) <= VNStageIntLLROutputS4xD(251)(4);
  CNStageIntLLRInputS5xD(89)(3) <= VNStageIntLLROutputS4xD(252)(0);
  CNStageIntLLRInputS5xD(112)(3) <= VNStageIntLLROutputS4xD(252)(1);
  CNStageIntLLRInputS5xD(199)(3) <= VNStageIntLLROutputS4xD(252)(2);
  CNStageIntLLRInputS5xD(239)(3) <= VNStageIntLLROutputS4xD(252)(3);
  CNStageIntLLRInputS5xD(325)(3) <= VNStageIntLLROutputS4xD(252)(4);
  CNStageIntLLRInputS5xD(373)(3) <= VNStageIntLLROutputS4xD(252)(5);
  CNStageIntLLRInputS5xD(80)(3) <= VNStageIntLLROutputS4xD(253)(0);
  CNStageIntLLRInputS5xD(121)(3) <= VNStageIntLLROutputS4xD(253)(1);
  CNStageIntLLRInputS5xD(211)(3) <= VNStageIntLLROutputS4xD(253)(2);
  CNStageIntLLRInputS5xD(279)(3) <= VNStageIntLLROutputS4xD(253)(3);
  CNStageIntLLRInputS5xD(283)(3) <= VNStageIntLLROutputS4xD(253)(4);
  CNStageIntLLRInputS5xD(380)(3) <= VNStageIntLLROutputS4xD(253)(5);
  CNStageIntLLRInputS5xD(67)(3) <= VNStageIntLLROutputS4xD(254)(0);
  CNStageIntLLRInputS5xD(222)(3) <= VNStageIntLLROutputS4xD(254)(1);
  CNStageIntLLRInputS5xD(238)(3) <= VNStageIntLLROutputS4xD(254)(2);
  CNStageIntLLRInputS5xD(290)(3) <= VNStageIntLLROutputS4xD(254)(3);
  CNStageIntLLRInputS5xD(362)(3) <= VNStageIntLLROutputS4xD(254)(4);
  CNStageIntLLRInputS5xD(52)(3) <= VNStageIntLLROutputS4xD(255)(0);
  CNStageIntLLRInputS5xD(86)(3) <= VNStageIntLLROutputS4xD(255)(1);
  CNStageIntLLRInputS5xD(167)(3) <= VNStageIntLLROutputS4xD(255)(2);
  CNStageIntLLRInputS5xD(195)(3) <= VNStageIntLLROutputS4xD(255)(3);
  CNStageIntLLRInputS5xD(233)(3) <= VNStageIntLLROutputS4xD(255)(4);
  CNStageIntLLRInputS5xD(318)(3) <= VNStageIntLLROutputS4xD(255)(5);
  CNStageIntLLRInputS5xD(364)(3) <= VNStageIntLLROutputS4xD(255)(6);
  CNStageIntLLRInputS5xD(53)(4) <= VNStageIntLLROutputS4xD(256)(0);
  CNStageIntLLRInputS5xD(106)(4) <= VNStageIntLLROutputS4xD(256)(1);
  CNStageIntLLRInputS5xD(127)(4) <= VNStageIntLLROutputS4xD(256)(2);
  CNStageIntLLRInputS5xD(242)(4) <= VNStageIntLLROutputS4xD(256)(3);
  CNStageIntLLRInputS5xD(296)(4) <= VNStageIntLLROutputS4xD(256)(4);
  CNStageIntLLRInputS5xD(339)(4) <= VNStageIntLLROutputS4xD(256)(5);
  CNStageIntLLRInputS5xD(51)(4) <= VNStageIntLLROutputS4xD(257)(0);
  CNStageIntLLRInputS5xD(85)(4) <= VNStageIntLLROutputS4xD(257)(1);
  CNStageIntLLRInputS5xD(166)(4) <= VNStageIntLLROutputS4xD(257)(2);
  CNStageIntLLRInputS5xD(194)(4) <= VNStageIntLLROutputS4xD(257)(3);
  CNStageIntLLRInputS5xD(232)(4) <= VNStageIntLLROutputS4xD(257)(4);
  CNStageIntLLRInputS5xD(317)(4) <= VNStageIntLLROutputS4xD(257)(5);
  CNStageIntLLRInputS5xD(363)(4) <= VNStageIntLLROutputS4xD(257)(6);
  CNStageIntLLRInputS5xD(50)(4) <= VNStageIntLLROutputS4xD(258)(0);
  CNStageIntLLRInputS5xD(57)(4) <= VNStageIntLLROutputS4xD(258)(1);
  CNStageIntLLRInputS5xD(331)(4) <= VNStageIntLLROutputS4xD(258)(2);
  CNStageIntLLRInputS5xD(54)(4) <= VNStageIntLLROutputS4xD(259)(0);
  CNStageIntLLRInputS5xD(114)(4) <= VNStageIntLLROutputS4xD(259)(1);
  CNStageIntLLRInputS5xD(274)(4) <= VNStageIntLLROutputS4xD(259)(2);
  CNStageIntLLRInputS5xD(303)(4) <= VNStageIntLLROutputS4xD(259)(3);
  CNStageIntLLRInputS5xD(370)(4) <= VNStageIntLLROutputS4xD(259)(4);
  CNStageIntLLRInputS5xD(49)(4) <= VNStageIntLLROutputS4xD(260)(0);
  CNStageIntLLRInputS5xD(71)(4) <= VNStageIntLLROutputS4xD(260)(1);
  CNStageIntLLRInputS5xD(138)(4) <= VNStageIntLLROutputS4xD(260)(2);
  CNStageIntLLRInputS5xD(186)(4) <= VNStageIntLLROutputS4xD(260)(3);
  CNStageIntLLRInputS5xD(243)(4) <= VNStageIntLLROutputS4xD(260)(4);
  CNStageIntLLRInputS5xD(383)(4) <= VNStageIntLLROutputS4xD(260)(5);
  CNStageIntLLRInputS5xD(48)(4) <= VNStageIntLLROutputS4xD(261)(0);
  CNStageIntLLRInputS5xD(63)(4) <= VNStageIntLLROutputS4xD(261)(1);
  CNStageIntLLRInputS5xD(152)(4) <= VNStageIntLLROutputS4xD(261)(2);
  CNStageIntLLRInputS5xD(204)(4) <= VNStageIntLLROutputS4xD(261)(3);
  CNStageIntLLRInputS5xD(305)(4) <= VNStageIntLLROutputS4xD(261)(4);
  CNStageIntLLRInputS5xD(333)(4) <= VNStageIntLLROutputS4xD(261)(5);
  CNStageIntLLRInputS5xD(47)(4) <= VNStageIntLLROutputS4xD(262)(0);
  CNStageIntLLRInputS5xD(95)(4) <= VNStageIntLLROutputS4xD(262)(1);
  CNStageIntLLRInputS5xD(149)(4) <= VNStageIntLLROutputS4xD(262)(2);
  CNStageIntLLRInputS5xD(212)(4) <= VNStageIntLLROutputS4xD(262)(3);
  CNStageIntLLRInputS5xD(319)(4) <= VNStageIntLLROutputS4xD(262)(4);
  CNStageIntLLRInputS5xD(362)(4) <= VNStageIntLLROutputS4xD(262)(5);
  CNStageIntLLRInputS5xD(46)(4) <= VNStageIntLLROutputS4xD(263)(0);
  CNStageIntLLRInputS5xD(104)(4) <= VNStageIntLLROutputS4xD(263)(1);
  CNStageIntLLRInputS5xD(169)(4) <= VNStageIntLLROutputS4xD(263)(2);
  CNStageIntLLRInputS5xD(207)(4) <= VNStageIntLLROutputS4xD(263)(3);
  CNStageIntLLRInputS5xD(253)(4) <= VNStageIntLLROutputS4xD(263)(4);
  CNStageIntLLRInputS5xD(315)(4) <= VNStageIntLLROutputS4xD(263)(5);
  CNStageIntLLRInputS5xD(378)(4) <= VNStageIntLLROutputS4xD(263)(6);
  CNStageIntLLRInputS5xD(45)(4) <= VNStageIntLLROutputS4xD(264)(0);
  CNStageIntLLRInputS5xD(98)(4) <= VNStageIntLLROutputS4xD(264)(1);
  CNStageIntLLRInputS5xD(132)(4) <= VNStageIntLLROutputS4xD(264)(2);
  CNStageIntLLRInputS5xD(213)(4) <= VNStageIntLLROutputS4xD(264)(3);
  CNStageIntLLRInputS5xD(256)(4) <= VNStageIntLLROutputS4xD(264)(4);
  CNStageIntLLRInputS5xD(281)(4) <= VNStageIntLLROutputS4xD(264)(5);
  CNStageIntLLRInputS5xD(349)(4) <= VNStageIntLLROutputS4xD(264)(6);
  CNStageIntLLRInputS5xD(44)(4) <= VNStageIntLLROutputS4xD(265)(0);
  CNStageIntLLRInputS5xD(133)(4) <= VNStageIntLLROutputS4xD(265)(1);
  CNStageIntLLRInputS5xD(203)(4) <= VNStageIntLLROutputS4xD(265)(2);
  CNStageIntLLRInputS5xD(244)(4) <= VNStageIntLLROutputS4xD(265)(3);
  CNStageIntLLRInputS5xD(43)(4) <= VNStageIntLLROutputS4xD(266)(0);
  CNStageIntLLRInputS5xD(168)(4) <= VNStageIntLLROutputS4xD(266)(1);
  CNStageIntLLRInputS5xD(173)(4) <= VNStageIntLLROutputS4xD(266)(2);
  CNStageIntLLRInputS5xD(273)(4) <= VNStageIntLLROutputS4xD(266)(3);
  CNStageIntLLRInputS5xD(300)(4) <= VNStageIntLLROutputS4xD(266)(4);
  CNStageIntLLRInputS5xD(42)(4) <= VNStageIntLLROutputS4xD(267)(0);
  CNStageIntLLRInputS5xD(72)(4) <= VNStageIntLLROutputS4xD(267)(1);
  CNStageIntLLRInputS5xD(159)(4) <= VNStageIntLLROutputS4xD(267)(2);
  CNStageIntLLRInputS5xD(180)(4) <= VNStageIntLLROutputS4xD(267)(3);
  CNStageIntLLRInputS5xD(241)(4) <= VNStageIntLLROutputS4xD(267)(4);
  CNStageIntLLRInputS5xD(280)(4) <= VNStageIntLLROutputS4xD(267)(5);
  CNStageIntLLRInputS5xD(364)(4) <= VNStageIntLLROutputS4xD(267)(6);
  CNStageIntLLRInputS5xD(41)(4) <= VNStageIntLLROutputS4xD(268)(0);
  CNStageIntLLRInputS5xD(109)(4) <= VNStageIntLLROutputS4xD(268)(1);
  CNStageIntLLRInputS5xD(118)(4) <= VNStageIntLLROutputS4xD(268)(2);
  CNStageIntLLRInputS5xD(216)(4) <= VNStageIntLLROutputS4xD(268)(3);
  CNStageIntLLRInputS5xD(266)(4) <= VNStageIntLLROutputS4xD(268)(4);
  CNStageIntLLRInputS5xD(325)(4) <= VNStageIntLLROutputS4xD(268)(5);
  CNStageIntLLRInputS5xD(360)(4) <= VNStageIntLLROutputS4xD(268)(6);
  CNStageIntLLRInputS5xD(67)(4) <= VNStageIntLLROutputS4xD(269)(0);
  CNStageIntLLRInputS5xD(122)(4) <= VNStageIntLLROutputS4xD(269)(1);
  CNStageIntLLRInputS5xD(218)(4) <= VNStageIntLLROutputS4xD(269)(2);
  CNStageIntLLRInputS5xD(250)(4) <= VNStageIntLLROutputS4xD(269)(3);
  CNStageIntLLRInputS5xD(287)(4) <= VNStageIntLLROutputS4xD(269)(4);
  CNStageIntLLRInputS5xD(381)(4) <= VNStageIntLLROutputS4xD(269)(5);
  CNStageIntLLRInputS5xD(40)(4) <= VNStageIntLLROutputS4xD(270)(0);
  CNStageIntLLRInputS5xD(79)(4) <= VNStageIntLLROutputS4xD(270)(1);
  CNStageIntLLRInputS5xD(170)(4) <= VNStageIntLLROutputS4xD(270)(2);
  CNStageIntLLRInputS5xD(190)(4) <= VNStageIntLLROutputS4xD(270)(3);
  CNStageIntLLRInputS5xD(275)(4) <= VNStageIntLLROutputS4xD(270)(4);
  CNStageIntLLRInputS5xD(292)(4) <= VNStageIntLLROutputS4xD(270)(5);
  CNStageIntLLRInputS5xD(344)(4) <= VNStageIntLLROutputS4xD(270)(6);
  CNStageIntLLRInputS5xD(39)(4) <= VNStageIntLLROutputS4xD(271)(0);
  CNStageIntLLRInputS5xD(105)(4) <= VNStageIntLLROutputS4xD(271)(1);
  CNStageIntLLRInputS5xD(171)(4) <= VNStageIntLLROutputS4xD(271)(2);
  CNStageIntLLRInputS5xD(268)(4) <= VNStageIntLLROutputS4xD(271)(3);
  CNStageIntLLRInputS5xD(332)(4) <= VNStageIntLLROutputS4xD(271)(4);
  CNStageIntLLRInputS5xD(345)(4) <= VNStageIntLLROutputS4xD(271)(5);
  CNStageIntLLRInputS5xD(38)(4) <= VNStageIntLLROutputS4xD(272)(0);
  CNStageIntLLRInputS5xD(94)(4) <= VNStageIntLLROutputS4xD(272)(1);
  CNStageIntLLRInputS5xD(116)(4) <= VNStageIntLLROutputS4xD(272)(2);
  CNStageIntLLRInputS5xD(184)(4) <= VNStageIntLLROutputS4xD(272)(3);
  CNStageIntLLRInputS5xD(254)(4) <= VNStageIntLLROutputS4xD(272)(4);
  CNStageIntLLRInputS5xD(291)(4) <= VNStageIntLLROutputS4xD(272)(5);
  CNStageIntLLRInputS5xD(380)(4) <= VNStageIntLLROutputS4xD(272)(6);
  CNStageIntLLRInputS5xD(37)(4) <= VNStageIntLLROutputS4xD(273)(0);
  CNStageIntLLRInputS5xD(81)(4) <= VNStageIntLLROutputS4xD(273)(1);
  CNStageIntLLRInputS5xD(156)(4) <= VNStageIntLLROutputS4xD(273)(2);
  CNStageIntLLRInputS5xD(272)(4) <= VNStageIntLLROutputS4xD(273)(3);
  CNStageIntLLRInputS5xD(285)(4) <= VNStageIntLLROutputS4xD(273)(4);
  CNStageIntLLRInputS5xD(371)(4) <= VNStageIntLLROutputS4xD(273)(5);
  CNStageIntLLRInputS5xD(36)(4) <= VNStageIntLLROutputS4xD(274)(0);
  CNStageIntLLRInputS5xD(164)(4) <= VNStageIntLLROutputS4xD(274)(1);
  CNStageIntLLRInputS5xD(217)(4) <= VNStageIntLLROutputS4xD(274)(2);
  CNStageIntLLRInputS5xD(248)(4) <= VNStageIntLLROutputS4xD(274)(3);
  CNStageIntLLRInputS5xD(35)(4) <= VNStageIntLLROutputS4xD(275)(0);
  CNStageIntLLRInputS5xD(59)(4) <= VNStageIntLLROutputS4xD(275)(1);
  CNStageIntLLRInputS5xD(128)(4) <= VNStageIntLLROutputS4xD(275)(2);
  CNStageIntLLRInputS5xD(179)(4) <= VNStageIntLLROutputS4xD(275)(3);
  CNStageIntLLRInputS5xD(329)(4) <= VNStageIntLLROutputS4xD(275)(4);
  CNStageIntLLRInputS5xD(34)(4) <= VNStageIntLLROutputS4xD(276)(0);
  CNStageIntLLRInputS5xD(69)(4) <= VNStageIntLLROutputS4xD(276)(1);
  CNStageIntLLRInputS5xD(126)(4) <= VNStageIntLLROutputS4xD(276)(2);
  CNStageIntLLRInputS5xD(205)(4) <= VNStageIntLLROutputS4xD(276)(3);
  CNStageIntLLRInputS5xD(259)(4) <= VNStageIntLLROutputS4xD(276)(4);
  CNStageIntLLRInputS5xD(297)(4) <= VNStageIntLLROutputS4xD(276)(5);
  CNStageIntLLRInputS5xD(33)(4) <= VNStageIntLLROutputS4xD(277)(0);
  CNStageIntLLRInputS5xD(64)(4) <= VNStageIntLLROutputS4xD(277)(1);
  CNStageIntLLRInputS5xD(162)(4) <= VNStageIntLLROutputS4xD(277)(2);
  CNStageIntLLRInputS5xD(185)(4) <= VNStageIntLLROutputS4xD(277)(3);
  CNStageIntLLRInputS5xD(252)(4) <= VNStageIntLLROutputS4xD(277)(4);
  CNStageIntLLRInputS5xD(295)(4) <= VNStageIntLLROutputS4xD(277)(5);
  CNStageIntLLRInputS5xD(334)(4) <= VNStageIntLLROutputS4xD(277)(6);
  CNStageIntLLRInputS5xD(32)(4) <= VNStageIntLLROutputS4xD(278)(0);
  CNStageIntLLRInputS5xD(70)(4) <= VNStageIntLLROutputS4xD(278)(1);
  CNStageIntLLRInputS5xD(141)(4) <= VNStageIntLLROutputS4xD(278)(2);
  CNStageIntLLRInputS5xD(229)(4) <= VNStageIntLLROutputS4xD(278)(3);
  CNStageIntLLRInputS5xD(328)(4) <= VNStageIntLLROutputS4xD(278)(4);
  CNStageIntLLRInputS5xD(31)(4) <= VNStageIntLLROutputS4xD(279)(0);
  CNStageIntLLRInputS5xD(58)(4) <= VNStageIntLLROutputS4xD(279)(1);
  CNStageIntLLRInputS5xD(144)(4) <= VNStageIntLLROutputS4xD(279)(2);
  CNStageIntLLRInputS5xD(219)(4) <= VNStageIntLLROutputS4xD(279)(3);
  CNStageIntLLRInputS5xD(239)(4) <= VNStageIntLLROutputS4xD(279)(4);
  CNStageIntLLRInputS5xD(368)(4) <= VNStageIntLLROutputS4xD(279)(5);
  CNStageIntLLRInputS5xD(30)(4) <= VNStageIntLLROutputS4xD(280)(0);
  CNStageIntLLRInputS5xD(84)(4) <= VNStageIntLLROutputS4xD(280)(1);
  CNStageIntLLRInputS5xD(129)(4) <= VNStageIntLLROutputS4xD(280)(2);
  CNStageIntLLRInputS5xD(215)(4) <= VNStageIntLLROutputS4xD(280)(3);
  CNStageIntLLRInputS5xD(233)(4) <= VNStageIntLLROutputS4xD(280)(4);
  CNStageIntLLRInputS5xD(310)(4) <= VNStageIntLLROutputS4xD(280)(5);
  CNStageIntLLRInputS5xD(376)(4) <= VNStageIntLLROutputS4xD(280)(6);
  CNStageIntLLRInputS5xD(29)(4) <= VNStageIntLLROutputS4xD(281)(0);
  CNStageIntLLRInputS5xD(90)(4) <= VNStageIntLLROutputS4xD(281)(1);
  CNStageIntLLRInputS5xD(163)(4) <= VNStageIntLLROutputS4xD(281)(2);
  CNStageIntLLRInputS5xD(182)(4) <= VNStageIntLLROutputS4xD(281)(3);
  CNStageIntLLRInputS5xD(236)(4) <= VNStageIntLLROutputS4xD(281)(4);
  CNStageIntLLRInputS5xD(298)(4) <= VNStageIntLLROutputS4xD(281)(5);
  CNStageIntLLRInputS5xD(340)(4) <= VNStageIntLLROutputS4xD(281)(6);
  CNStageIntLLRInputS5xD(28)(4) <= VNStageIntLLROutputS4xD(282)(0);
  CNStageIntLLRInputS5xD(74)(4) <= VNStageIntLLROutputS4xD(282)(1);
  CNStageIntLLRInputS5xD(125)(4) <= VNStageIntLLROutputS4xD(282)(2);
  CNStageIntLLRInputS5xD(200)(4) <= VNStageIntLLROutputS4xD(282)(3);
  CNStageIntLLRInputS5xD(226)(4) <= VNStageIntLLROutputS4xD(282)(4);
  CNStageIntLLRInputS5xD(338)(4) <= VNStageIntLLROutputS4xD(282)(5);
  CNStageIntLLRInputS5xD(27)(4) <= VNStageIntLLROutputS4xD(283)(0);
  CNStageIntLLRInputS5xD(76)(4) <= VNStageIntLLROutputS4xD(283)(1);
  CNStageIntLLRInputS5xD(153)(4) <= VNStageIntLLROutputS4xD(283)(2);
  CNStageIntLLRInputS5xD(201)(4) <= VNStageIntLLROutputS4xD(283)(3);
  CNStageIntLLRInputS5xD(260)(4) <= VNStageIntLLROutputS4xD(283)(4);
  CNStageIntLLRInputS5xD(294)(4) <= VNStageIntLLROutputS4xD(283)(5);
  CNStageIntLLRInputS5xD(374)(4) <= VNStageIntLLROutputS4xD(283)(6);
  CNStageIntLLRInputS5xD(26)(4) <= VNStageIntLLROutputS4xD(284)(0);
  CNStageIntLLRInputS5xD(100)(4) <= VNStageIntLLROutputS4xD(284)(1);
  CNStageIntLLRInputS5xD(137)(4) <= VNStageIntLLROutputS4xD(284)(2);
  CNStageIntLLRInputS5xD(181)(4) <= VNStageIntLLROutputS4xD(284)(3);
  CNStageIntLLRInputS5xD(245)(4) <= VNStageIntLLROutputS4xD(284)(4);
  CNStageIntLLRInputS5xD(320)(4) <= VNStageIntLLROutputS4xD(284)(5);
  CNStageIntLLRInputS5xD(353)(4) <= VNStageIntLLROutputS4xD(284)(6);
  CNStageIntLLRInputS5xD(25)(4) <= VNStageIntLLROutputS4xD(285)(0);
  CNStageIntLLRInputS5xD(82)(4) <= VNStageIntLLROutputS4xD(285)(1);
  CNStageIntLLRInputS5xD(165)(4) <= VNStageIntLLROutputS4xD(285)(2);
  CNStageIntLLRInputS5xD(172)(4) <= VNStageIntLLROutputS4xD(285)(3);
  CNStageIntLLRInputS5xD(255)(4) <= VNStageIntLLROutputS4xD(285)(4);
  CNStageIntLLRInputS5xD(304)(4) <= VNStageIntLLROutputS4xD(285)(5);
  CNStageIntLLRInputS5xD(355)(4) <= VNStageIntLLROutputS4xD(285)(6);
  CNStageIntLLRInputS5xD(24)(4) <= VNStageIntLLROutputS4xD(286)(0);
  CNStageIntLLRInputS5xD(93)(4) <= VNStageIntLLROutputS4xD(286)(1);
  CNStageIntLLRInputS5xD(155)(4) <= VNStageIntLLROutputS4xD(286)(2);
  CNStageIntLLRInputS5xD(189)(4) <= VNStageIntLLROutputS4xD(286)(3);
  CNStageIntLLRInputS5xD(267)(4) <= VNStageIntLLROutputS4xD(286)(4);
  CNStageIntLLRInputS5xD(330)(4) <= VNStageIntLLROutputS4xD(286)(5);
  CNStageIntLLRInputS5xD(341)(4) <= VNStageIntLLROutputS4xD(286)(6);
  CNStageIntLLRInputS5xD(23)(4) <= VNStageIntLLROutputS4xD(287)(0);
  CNStageIntLLRInputS5xD(101)(4) <= VNStageIntLLROutputS4xD(287)(1);
  CNStageIntLLRInputS5xD(142)(4) <= VNStageIntLLROutputS4xD(287)(2);
  CNStageIntLLRInputS5xD(193)(4) <= VNStageIntLLROutputS4xD(287)(3);
  CNStageIntLLRInputS5xD(240)(4) <= VNStageIntLLROutputS4xD(287)(4);
  CNStageIntLLRInputS5xD(322)(4) <= VNStageIntLLROutputS4xD(287)(5);
  CNStageIntLLRInputS5xD(375)(4) <= VNStageIntLLROutputS4xD(287)(6);
  CNStageIntLLRInputS5xD(22)(4) <= VNStageIntLLROutputS4xD(288)(0);
  CNStageIntLLRInputS5xD(75)(4) <= VNStageIntLLROutputS4xD(288)(1);
  CNStageIntLLRInputS5xD(161)(4) <= VNStageIntLLROutputS4xD(288)(2);
  CNStageIntLLRInputS5xD(224)(4) <= VNStageIntLLROutputS4xD(288)(3);
  CNStageIntLLRInputS5xD(228)(4) <= VNStageIntLLROutputS4xD(288)(4);
  CNStageIntLLRInputS5xD(308)(4) <= VNStageIntLLROutputS4xD(288)(5);
  CNStageIntLLRInputS5xD(337)(4) <= VNStageIntLLROutputS4xD(288)(6);
  CNStageIntLLRInputS5xD(21)(4) <= VNStageIntLLROutputS4xD(289)(0);
  CNStageIntLLRInputS5xD(89)(4) <= VNStageIntLLROutputS4xD(289)(1);
  CNStageIntLLRInputS5xD(134)(4) <= VNStageIntLLROutputS4xD(289)(2);
  CNStageIntLLRInputS5xD(192)(4) <= VNStageIntLLROutputS4xD(289)(3);
  CNStageIntLLRInputS5xD(269)(4) <= VNStageIntLLROutputS4xD(289)(4);
  CNStageIntLLRInputS5xD(327)(4) <= VNStageIntLLROutputS4xD(289)(5);
  CNStageIntLLRInputS5xD(365)(4) <= VNStageIntLLROutputS4xD(289)(6);
  CNStageIntLLRInputS5xD(20)(4) <= VNStageIntLLROutputS4xD(290)(0);
  CNStageIntLLRInputS5xD(60)(4) <= VNStageIntLLROutputS4xD(290)(1);
  CNStageIntLLRInputS5xD(131)(4) <= VNStageIntLLROutputS4xD(290)(2);
  CNStageIntLLRInputS5xD(187)(4) <= VNStageIntLLROutputS4xD(290)(3);
  CNStageIntLLRInputS5xD(231)(4) <= VNStageIntLLROutputS4xD(290)(4);
  CNStageIntLLRInputS5xD(350)(4) <= VNStageIntLLROutputS4xD(290)(5);
  CNStageIntLLRInputS5xD(19)(4) <= VNStageIntLLROutputS4xD(291)(0);
  CNStageIntLLRInputS5xD(96)(4) <= VNStageIntLLROutputS4xD(291)(1);
  CNStageIntLLRInputS5xD(147)(4) <= VNStageIntLLROutputS4xD(291)(2);
  CNStageIntLLRInputS5xD(223)(4) <= VNStageIntLLROutputS4xD(291)(3);
  CNStageIntLLRInputS5xD(249)(4) <= VNStageIntLLROutputS4xD(291)(4);
  CNStageIntLLRInputS5xD(377)(4) <= VNStageIntLLROutputS4xD(291)(5);
  CNStageIntLLRInputS5xD(18)(4) <= VNStageIntLLROutputS4xD(292)(0);
  CNStageIntLLRInputS5xD(62)(4) <= VNStageIntLLROutputS4xD(292)(1);
  CNStageIntLLRInputS5xD(139)(4) <= VNStageIntLLROutputS4xD(292)(2);
  CNStageIntLLRInputS5xD(177)(4) <= VNStageIntLLROutputS4xD(292)(3);
  CNStageIntLLRInputS5xD(257)(4) <= VNStageIntLLROutputS4xD(292)(4);
  CNStageIntLLRInputS5xD(313)(4) <= VNStageIntLLROutputS4xD(292)(5);
  CNStageIntLLRInputS5xD(367)(4) <= VNStageIntLLROutputS4xD(292)(6);
  CNStageIntLLRInputS5xD(17)(4) <= VNStageIntLLROutputS4xD(293)(0);
  CNStageIntLLRInputS5xD(77)(4) <= VNStageIntLLROutputS4xD(293)(1);
  CNStageIntLLRInputS5xD(113)(4) <= VNStageIntLLROutputS4xD(293)(2);
  CNStageIntLLRInputS5xD(197)(4) <= VNStageIntLLROutputS4xD(293)(3);
  CNStageIntLLRInputS5xD(306)(4) <= VNStageIntLLROutputS4xD(293)(4);
  CNStageIntLLRInputS5xD(354)(4) <= VNStageIntLLROutputS4xD(293)(5);
  CNStageIntLLRInputS5xD(16)(4) <= VNStageIntLLROutputS4xD(294)(0);
  CNStageIntLLRInputS5xD(73)(4) <= VNStageIntLLROutputS4xD(294)(1);
  CNStageIntLLRInputS5xD(123)(4) <= VNStageIntLLROutputS4xD(294)(2);
  CNStageIntLLRInputS5xD(196)(4) <= VNStageIntLLROutputS4xD(294)(3);
  CNStageIntLLRInputS5xD(258)(4) <= VNStageIntLLROutputS4xD(294)(4);
  CNStageIntLLRInputS5xD(284)(4) <= VNStageIntLLROutputS4xD(294)(5);
  CNStageIntLLRInputS5xD(373)(4) <= VNStageIntLLROutputS4xD(294)(6);
  CNStageIntLLRInputS5xD(15)(4) <= VNStageIntLLROutputS4xD(295)(0);
  CNStageIntLLRInputS5xD(92)(4) <= VNStageIntLLROutputS4xD(295)(1);
  CNStageIntLLRInputS5xD(117)(4) <= VNStageIntLLROutputS4xD(295)(2);
  CNStageIntLLRInputS5xD(175)(4) <= VNStageIntLLROutputS4xD(295)(3);
  CNStageIntLLRInputS5xD(346)(4) <= VNStageIntLLROutputS4xD(295)(4);
  CNStageIntLLRInputS5xD(14)(4) <= VNStageIntLLROutputS4xD(296)(0);
  CNStageIntLLRInputS5xD(55)(4) <= VNStageIntLLROutputS4xD(296)(1);
  CNStageIntLLRInputS5xD(121)(4) <= VNStageIntLLROutputS4xD(296)(2);
  CNStageIntLLRInputS5xD(208)(4) <= VNStageIntLLROutputS4xD(296)(3);
  CNStageIntLLRInputS5xD(286)(4) <= VNStageIntLLROutputS4xD(296)(4);
  CNStageIntLLRInputS5xD(343)(4) <= VNStageIntLLROutputS4xD(296)(5);
  CNStageIntLLRInputS5xD(13)(4) <= VNStageIntLLROutputS4xD(297)(0);
  CNStageIntLLRInputS5xD(56)(4) <= VNStageIntLLROutputS4xD(297)(1);
  CNStageIntLLRInputS5xD(111)(4) <= VNStageIntLLROutputS4xD(297)(2);
  CNStageIntLLRInputS5xD(211)(4) <= VNStageIntLLROutputS4xD(297)(3);
  CNStageIntLLRInputS5xD(277)(4) <= VNStageIntLLROutputS4xD(297)(4);
  CNStageIntLLRInputS5xD(290)(4) <= VNStageIntLLROutputS4xD(297)(5);
  CNStageIntLLRInputS5xD(358)(4) <= VNStageIntLLROutputS4xD(297)(6);
  CNStageIntLLRInputS5xD(12)(4) <= VNStageIntLLROutputS4xD(298)(0);
  CNStageIntLLRInputS5xD(91)(4) <= VNStageIntLLROutputS4xD(298)(1);
  CNStageIntLLRInputS5xD(148)(4) <= VNStageIntLLROutputS4xD(298)(2);
  CNStageIntLLRInputS5xD(198)(4) <= VNStageIntLLROutputS4xD(298)(3);
  CNStageIntLLRInputS5xD(262)(4) <= VNStageIntLLROutputS4xD(298)(4);
  CNStageIntLLRInputS5xD(282)(4) <= VNStageIntLLROutputS4xD(298)(5);
  CNStageIntLLRInputS5xD(351)(4) <= VNStageIntLLROutputS4xD(298)(6);
  CNStageIntLLRInputS5xD(83)(4) <= VNStageIntLLROutputS4xD(299)(0);
  CNStageIntLLRInputS5xD(130)(4) <= VNStageIntLLROutputS4xD(299)(1);
  CNStageIntLLRInputS5xD(176)(4) <= VNStageIntLLROutputS4xD(299)(2);
  CNStageIntLLRInputS5xD(264)(4) <= VNStageIntLLROutputS4xD(299)(3);
  CNStageIntLLRInputS5xD(314)(4) <= VNStageIntLLROutputS4xD(299)(4);
  CNStageIntLLRInputS5xD(11)(4) <= VNStageIntLLROutputS4xD(300)(0);
  CNStageIntLLRInputS5xD(99)(4) <= VNStageIntLLROutputS4xD(300)(1);
  CNStageIntLLRInputS5xD(143)(4) <= VNStageIntLLROutputS4xD(300)(2);
  CNStageIntLLRInputS5xD(195)(4) <= VNStageIntLLROutputS4xD(300)(3);
  CNStageIntLLRInputS5xD(299)(4) <= VNStageIntLLROutputS4xD(300)(4);
  CNStageIntLLRInputS5xD(335)(4) <= VNStageIntLLROutputS4xD(300)(5);
  CNStageIntLLRInputS5xD(10)(4) <= VNStageIntLLROutputS4xD(301)(0);
  CNStageIntLLRInputS5xD(103)(4) <= VNStageIntLLROutputS4xD(301)(1);
  CNStageIntLLRInputS5xD(154)(4) <= VNStageIntLLROutputS4xD(301)(2);
  CNStageIntLLRInputS5xD(220)(4) <= VNStageIntLLROutputS4xD(301)(3);
  CNStageIntLLRInputS5xD(270)(4) <= VNStageIntLLROutputS4xD(301)(4);
  CNStageIntLLRInputS5xD(309)(4) <= VNStageIntLLROutputS4xD(301)(5);
  CNStageIntLLRInputS5xD(9)(4) <= VNStageIntLLROutputS4xD(302)(0);
  CNStageIntLLRInputS5xD(110)(4) <= VNStageIntLLROutputS4xD(302)(1);
  CNStageIntLLRInputS5xD(124)(4) <= VNStageIntLLROutputS4xD(302)(2);
  CNStageIntLLRInputS5xD(206)(4) <= VNStageIntLLROutputS4xD(302)(3);
  CNStageIntLLRInputS5xD(227)(4) <= VNStageIntLLROutputS4xD(302)(4);
  CNStageIntLLRInputS5xD(321)(4) <= VNStageIntLLROutputS4xD(302)(5);
  CNStageIntLLRInputS5xD(8)(4) <= VNStageIntLLROutputS4xD(303)(0);
  CNStageIntLLRInputS5xD(102)(4) <= VNStageIntLLROutputS4xD(303)(1);
  CNStageIntLLRInputS5xD(112)(4) <= VNStageIntLLROutputS4xD(303)(2);
  CNStageIntLLRInputS5xD(178)(4) <= VNStageIntLLROutputS4xD(303)(3);
  CNStageIntLLRInputS5xD(235)(4) <= VNStageIntLLROutputS4xD(303)(4);
  CNStageIntLLRInputS5xD(293)(4) <= VNStageIntLLROutputS4xD(303)(5);
  CNStageIntLLRInputS5xD(382)(4) <= VNStageIntLLROutputS4xD(303)(6);
  CNStageIntLLRInputS5xD(7)(4) <= VNStageIntLLROutputS4xD(304)(0);
  CNStageIntLLRInputS5xD(97)(4) <= VNStageIntLLROutputS4xD(304)(1);
  CNStageIntLLRInputS5xD(157)(4) <= VNStageIntLLROutputS4xD(304)(2);
  CNStageIntLLRInputS5xD(222)(4) <= VNStageIntLLROutputS4xD(304)(3);
  CNStageIntLLRInputS5xD(263)(4) <= VNStageIntLLROutputS4xD(304)(4);
  CNStageIntLLRInputS5xD(283)(4) <= VNStageIntLLROutputS4xD(304)(5);
  CNStageIntLLRInputS5xD(359)(4) <= VNStageIntLLROutputS4xD(304)(6);
  CNStageIntLLRInputS5xD(6)(4) <= VNStageIntLLROutputS4xD(305)(0);
  CNStageIntLLRInputS5xD(80)(4) <= VNStageIntLLROutputS4xD(305)(1);
  CNStageIntLLRInputS5xD(115)(4) <= VNStageIntLLROutputS4xD(305)(2);
  CNStageIntLLRInputS5xD(209)(4) <= VNStageIntLLROutputS4xD(305)(3);
  CNStageIntLLRInputS5xD(276)(4) <= VNStageIntLLROutputS4xD(305)(4);
  CNStageIntLLRInputS5xD(323)(4) <= VNStageIntLLROutputS4xD(305)(5);
  CNStageIntLLRInputS5xD(342)(4) <= VNStageIntLLROutputS4xD(305)(6);
  CNStageIntLLRInputS5xD(5)(4) <= VNStageIntLLROutputS4xD(306)(0);
  CNStageIntLLRInputS5xD(87)(4) <= VNStageIntLLROutputS4xD(306)(1);
  CNStageIntLLRInputS5xD(136)(4) <= VNStageIntLLROutputS4xD(306)(2);
  CNStageIntLLRInputS5xD(174)(4) <= VNStageIntLLROutputS4xD(306)(3);
  CNStageIntLLRInputS5xD(4)(4) <= VNStageIntLLROutputS4xD(307)(0);
  CNStageIntLLRInputS5xD(107)(4) <= VNStageIntLLROutputS4xD(307)(1);
  CNStageIntLLRInputS5xD(145)(4) <= VNStageIntLLROutputS4xD(307)(2);
  CNStageIntLLRInputS5xD(202)(4) <= VNStageIntLLROutputS4xD(307)(3);
  CNStageIntLLRInputS5xD(230)(4) <= VNStageIntLLROutputS4xD(307)(4);
  CNStageIntLLRInputS5xD(302)(4) <= VNStageIntLLROutputS4xD(307)(5);
  CNStageIntLLRInputS5xD(366)(4) <= VNStageIntLLROutputS4xD(307)(6);
  CNStageIntLLRInputS5xD(140)(4) <= VNStageIntLLROutputS4xD(308)(0);
  CNStageIntLLRInputS5xD(199)(4) <= VNStageIntLLROutputS4xD(308)(1);
  CNStageIntLLRInputS5xD(251)(4) <= VNStageIntLLROutputS4xD(308)(2);
  CNStageIntLLRInputS5xD(311)(4) <= VNStageIntLLROutputS4xD(308)(3);
  CNStageIntLLRInputS5xD(336)(4) <= VNStageIntLLROutputS4xD(308)(4);
  CNStageIntLLRInputS5xD(3)(4) <= VNStageIntLLROutputS4xD(309)(0);
  CNStageIntLLRInputS5xD(86)(4) <= VNStageIntLLROutputS4xD(309)(1);
  CNStageIntLLRInputS5xD(146)(4) <= VNStageIntLLROutputS4xD(309)(2);
  CNStageIntLLRInputS5xD(214)(4) <= VNStageIntLLROutputS4xD(309)(3);
  CNStageIntLLRInputS5xD(265)(4) <= VNStageIntLLROutputS4xD(309)(4);
  CNStageIntLLRInputS5xD(307)(4) <= VNStageIntLLROutputS4xD(309)(5);
  CNStageIntLLRInputS5xD(2)(4) <= VNStageIntLLROutputS4xD(310)(0);
  CNStageIntLLRInputS5xD(65)(4) <= VNStageIntLLROutputS4xD(310)(1);
  CNStageIntLLRInputS5xD(135)(4) <= VNStageIntLLROutputS4xD(310)(2);
  CNStageIntLLRInputS5xD(261)(4) <= VNStageIntLLROutputS4xD(310)(3);
  CNStageIntLLRInputS5xD(312)(4) <= VNStageIntLLROutputS4xD(310)(4);
  CNStageIntLLRInputS5xD(369)(4) <= VNStageIntLLROutputS4xD(310)(5);
  CNStageIntLLRInputS5xD(1)(4) <= VNStageIntLLROutputS4xD(311)(0);
  CNStageIntLLRInputS5xD(68)(4) <= VNStageIntLLROutputS4xD(311)(1);
  CNStageIntLLRInputS5xD(160)(4) <= VNStageIntLLROutputS4xD(311)(2);
  CNStageIntLLRInputS5xD(225)(4) <= VNStageIntLLROutputS4xD(311)(3);
  CNStageIntLLRInputS5xD(301)(4) <= VNStageIntLLROutputS4xD(311)(4);
  CNStageIntLLRInputS5xD(0)(4) <= VNStageIntLLROutputS4xD(312)(0);
  CNStageIntLLRInputS5xD(108)(4) <= VNStageIntLLROutputS4xD(312)(1);
  CNStageIntLLRInputS5xD(167)(4) <= VNStageIntLLROutputS4xD(312)(2);
  CNStageIntLLRInputS5xD(246)(4) <= VNStageIntLLROutputS4xD(312)(3);
  CNStageIntLLRInputS5xD(326)(4) <= VNStageIntLLROutputS4xD(312)(4);
  CNStageIntLLRInputS5xD(348)(4) <= VNStageIntLLROutputS4xD(312)(5);
  CNStageIntLLRInputS5xD(150)(4) <= VNStageIntLLROutputS4xD(313)(0);
  CNStageIntLLRInputS5xD(188)(4) <= VNStageIntLLROutputS4xD(313)(1);
  CNStageIntLLRInputS5xD(247)(4) <= VNStageIntLLROutputS4xD(313)(2);
  CNStageIntLLRInputS5xD(356)(4) <= VNStageIntLLROutputS4xD(313)(3);
  CNStageIntLLRInputS5xD(191)(4) <= VNStageIntLLROutputS4xD(314)(0);
  CNStageIntLLRInputS5xD(278)(4) <= VNStageIntLLROutputS4xD(314)(1);
  CNStageIntLLRInputS5xD(316)(4) <= VNStageIntLLROutputS4xD(314)(2);
  CNStageIntLLRInputS5xD(352)(4) <= VNStageIntLLROutputS4xD(314)(3);
  CNStageIntLLRInputS5xD(78)(4) <= VNStageIntLLROutputS4xD(315)(0);
  CNStageIntLLRInputS5xD(119)(4) <= VNStageIntLLROutputS4xD(315)(1);
  CNStageIntLLRInputS5xD(183)(4) <= VNStageIntLLROutputS4xD(315)(2);
  CNStageIntLLRInputS5xD(271)(4) <= VNStageIntLLROutputS4xD(315)(3);
  CNStageIntLLRInputS5xD(318)(4) <= VNStageIntLLROutputS4xD(315)(4);
  CNStageIntLLRInputS5xD(357)(4) <= VNStageIntLLROutputS4xD(315)(5);
  CNStageIntLLRInputS5xD(61)(4) <= VNStageIntLLROutputS4xD(316)(0);
  CNStageIntLLRInputS5xD(158)(4) <= VNStageIntLLROutputS4xD(316)(1);
  CNStageIntLLRInputS5xD(234)(4) <= VNStageIntLLROutputS4xD(316)(2);
  CNStageIntLLRInputS5xD(288)(4) <= VNStageIntLLROutputS4xD(316)(3);
  CNStageIntLLRInputS5xD(347)(4) <= VNStageIntLLROutputS4xD(316)(4);
  CNStageIntLLRInputS5xD(88)(4) <= VNStageIntLLROutputS4xD(317)(0);
  CNStageIntLLRInputS5xD(238)(4) <= VNStageIntLLROutputS4xD(317)(1);
  CNStageIntLLRInputS5xD(324)(4) <= VNStageIntLLROutputS4xD(317)(2);
  CNStageIntLLRInputS5xD(372)(4) <= VNStageIntLLROutputS4xD(317)(3);
  CNStageIntLLRInputS5xD(120)(4) <= VNStageIntLLROutputS4xD(318)(0);
  CNStageIntLLRInputS5xD(210)(4) <= VNStageIntLLROutputS4xD(318)(1);
  CNStageIntLLRInputS5xD(279)(4) <= VNStageIntLLROutputS4xD(318)(2);
  CNStageIntLLRInputS5xD(379)(4) <= VNStageIntLLROutputS4xD(318)(3);
  CNStageIntLLRInputS5xD(52)(4) <= VNStageIntLLROutputS4xD(319)(0);
  CNStageIntLLRInputS5xD(66)(4) <= VNStageIntLLROutputS4xD(319)(1);
  CNStageIntLLRInputS5xD(151)(4) <= VNStageIntLLROutputS4xD(319)(2);
  CNStageIntLLRInputS5xD(221)(4) <= VNStageIntLLROutputS4xD(319)(3);
  CNStageIntLLRInputS5xD(237)(4) <= VNStageIntLLROutputS4xD(319)(4);
  CNStageIntLLRInputS5xD(289)(4) <= VNStageIntLLROutputS4xD(319)(5);
  CNStageIntLLRInputS5xD(361)(4) <= VNStageIntLLROutputS4xD(319)(6);
  CNStageIntLLRInputS5xD(53)(5) <= VNStageIntLLROutputS4xD(320)(0);
  CNStageIntLLRInputS5xD(126)(5) <= VNStageIntLLROutputS4xD(320)(1);
  CNStageIntLLRInputS5xD(196)(5) <= VNStageIntLLROutputS4xD(320)(2);
  CNStageIntLLRInputS5xD(295)(5) <= VNStageIntLLROutputS4xD(320)(3);
  CNStageIntLLRInputS5xD(338)(5) <= VNStageIntLLROutputS4xD(320)(4);
  CNStageIntLLRInputS5xD(51)(5) <= VNStageIntLLROutputS4xD(321)(0);
  CNStageIntLLRInputS5xD(65)(5) <= VNStageIntLLROutputS4xD(321)(1);
  CNStageIntLLRInputS5xD(150)(5) <= VNStageIntLLROutputS4xD(321)(2);
  CNStageIntLLRInputS5xD(220)(5) <= VNStageIntLLROutputS4xD(321)(3);
  CNStageIntLLRInputS5xD(236)(5) <= VNStageIntLLROutputS4xD(321)(4);
  CNStageIntLLRInputS5xD(288)(5) <= VNStageIntLLROutputS4xD(321)(5);
  CNStageIntLLRInputS5xD(360)(5) <= VNStageIntLLROutputS4xD(321)(6);
  CNStageIntLLRInputS5xD(50)(5) <= VNStageIntLLROutputS4xD(322)(0);
  CNStageIntLLRInputS5xD(84)(5) <= VNStageIntLLROutputS4xD(322)(1);
  CNStageIntLLRInputS5xD(165)(5) <= VNStageIntLLROutputS4xD(322)(2);
  CNStageIntLLRInputS5xD(231)(5) <= VNStageIntLLROutputS4xD(322)(3);
  CNStageIntLLRInputS5xD(316)(5) <= VNStageIntLLROutputS4xD(322)(4);
  CNStageIntLLRInputS5xD(362)(5) <= VNStageIntLLROutputS4xD(322)(5);
  CNStageIntLLRInputS5xD(56)(5) <= VNStageIntLLROutputS4xD(323)(0);
  CNStageIntLLRInputS5xD(136)(5) <= VNStageIntLLROutputS4xD(323)(1);
  CNStageIntLLRInputS5xD(184)(5) <= VNStageIntLLROutputS4xD(323)(2);
  CNStageIntLLRInputS5xD(268)(5) <= VNStageIntLLROutputS4xD(323)(3);
  CNStageIntLLRInputS5xD(330)(5) <= VNStageIntLLROutputS4xD(323)(4);
  CNStageIntLLRInputS5xD(49)(5) <= VNStageIntLLROutputS4xD(324)(0);
  CNStageIntLLRInputS5xD(109)(5) <= VNStageIntLLROutputS4xD(324)(1);
  CNStageIntLLRInputS5xD(113)(5) <= VNStageIntLLROutputS4xD(324)(2);
  CNStageIntLLRInputS5xD(223)(5) <= VNStageIntLLROutputS4xD(324)(3);
  CNStageIntLLRInputS5xD(273)(5) <= VNStageIntLLROutputS4xD(324)(4);
  CNStageIntLLRInputS5xD(302)(5) <= VNStageIntLLROutputS4xD(324)(5);
  CNStageIntLLRInputS5xD(369)(5) <= VNStageIntLLROutputS4xD(324)(6);
  CNStageIntLLRInputS5xD(48)(5) <= VNStageIntLLROutputS4xD(325)(0);
  CNStageIntLLRInputS5xD(70)(5) <= VNStageIntLLROutputS4xD(325)(1);
  CNStageIntLLRInputS5xD(137)(5) <= VNStageIntLLROutputS4xD(325)(2);
  CNStageIntLLRInputS5xD(185)(5) <= VNStageIntLLROutputS4xD(325)(3);
  CNStageIntLLRInputS5xD(242)(5) <= VNStageIntLLROutputS4xD(325)(4);
  CNStageIntLLRInputS5xD(284)(5) <= VNStageIntLLROutputS4xD(325)(5);
  CNStageIntLLRInputS5xD(382)(5) <= VNStageIntLLROutputS4xD(325)(6);
  CNStageIntLLRInputS5xD(47)(5) <= VNStageIntLLROutputS4xD(326)(0);
  CNStageIntLLRInputS5xD(62)(5) <= VNStageIntLLROutputS4xD(326)(1);
  CNStageIntLLRInputS5xD(203)(5) <= VNStageIntLLROutputS4xD(326)(2);
  CNStageIntLLRInputS5xD(241)(5) <= VNStageIntLLROutputS4xD(326)(3);
  CNStageIntLLRInputS5xD(304)(5) <= VNStageIntLLROutputS4xD(326)(4);
  CNStageIntLLRInputS5xD(46)(5) <= VNStageIntLLROutputS4xD(327)(0);
  CNStageIntLLRInputS5xD(94)(5) <= VNStageIntLLROutputS4xD(327)(1);
  CNStageIntLLRInputS5xD(148)(5) <= VNStageIntLLROutputS4xD(327)(2);
  CNStageIntLLRInputS5xD(211)(5) <= VNStageIntLLROutputS4xD(327)(3);
  CNStageIntLLRInputS5xD(272)(5) <= VNStageIntLLROutputS4xD(327)(4);
  CNStageIntLLRInputS5xD(318)(5) <= VNStageIntLLROutputS4xD(327)(5);
  CNStageIntLLRInputS5xD(361)(5) <= VNStageIntLLROutputS4xD(327)(6);
  CNStageIntLLRInputS5xD(45)(5) <= VNStageIntLLROutputS4xD(328)(0);
  CNStageIntLLRInputS5xD(103)(5) <= VNStageIntLLROutputS4xD(328)(1);
  CNStageIntLLRInputS5xD(168)(5) <= VNStageIntLLROutputS4xD(328)(2);
  CNStageIntLLRInputS5xD(314)(5) <= VNStageIntLLROutputS4xD(328)(3);
  CNStageIntLLRInputS5xD(377)(5) <= VNStageIntLLROutputS4xD(328)(4);
  CNStageIntLLRInputS5xD(44)(5) <= VNStageIntLLROutputS4xD(329)(0);
  CNStageIntLLRInputS5xD(97)(5) <= VNStageIntLLROutputS4xD(329)(1);
  CNStageIntLLRInputS5xD(131)(5) <= VNStageIntLLROutputS4xD(329)(2);
  CNStageIntLLRInputS5xD(212)(5) <= VNStageIntLLROutputS4xD(329)(3);
  CNStageIntLLRInputS5xD(255)(5) <= VNStageIntLLROutputS4xD(329)(4);
  CNStageIntLLRInputS5xD(280)(5) <= VNStageIntLLROutputS4xD(329)(5);
  CNStageIntLLRInputS5xD(348)(5) <= VNStageIntLLROutputS4xD(329)(6);
  CNStageIntLLRInputS5xD(43)(5) <= VNStageIntLLROutputS4xD(330)(0);
  CNStageIntLLRInputS5xD(101)(5) <= VNStageIntLLROutputS4xD(330)(1);
  CNStageIntLLRInputS5xD(132)(5) <= VNStageIntLLROutputS4xD(330)(2);
  CNStageIntLLRInputS5xD(202)(5) <= VNStageIntLLROutputS4xD(330)(3);
  CNStageIntLLRInputS5xD(243)(5) <= VNStageIntLLROutputS4xD(330)(4);
  CNStageIntLLRInputS5xD(42)(5) <= VNStageIntLLROutputS4xD(331)(0);
  CNStageIntLLRInputS5xD(92)(5) <= VNStageIntLLROutputS4xD(331)(1);
  CNStageIntLLRInputS5xD(167)(5) <= VNStageIntLLROutputS4xD(331)(2);
  CNStageIntLLRInputS5xD(172)(5) <= VNStageIntLLROutputS4xD(331)(3);
  CNStageIntLLRInputS5xD(350)(5) <= VNStageIntLLROutputS4xD(331)(4);
  CNStageIntLLRInputS5xD(41)(5) <= VNStageIntLLROutputS4xD(332)(0);
  CNStageIntLLRInputS5xD(71)(5) <= VNStageIntLLROutputS4xD(332)(1);
  CNStageIntLLRInputS5xD(158)(5) <= VNStageIntLLROutputS4xD(332)(2);
  CNStageIntLLRInputS5xD(179)(5) <= VNStageIntLLROutputS4xD(332)(3);
  CNStageIntLLRInputS5xD(240)(5) <= VNStageIntLLROutputS4xD(332)(4);
  CNStageIntLLRInputS5xD(363)(5) <= VNStageIntLLROutputS4xD(332)(5);
  CNStageIntLLRInputS5xD(108)(5) <= VNStageIntLLROutputS4xD(333)(0);
  CNStageIntLLRInputS5xD(117)(5) <= VNStageIntLLROutputS4xD(333)(1);
  CNStageIntLLRInputS5xD(215)(5) <= VNStageIntLLROutputS4xD(333)(2);
  CNStageIntLLRInputS5xD(265)(5) <= VNStageIntLLROutputS4xD(333)(3);
  CNStageIntLLRInputS5xD(324)(5) <= VNStageIntLLROutputS4xD(333)(4);
  CNStageIntLLRInputS5xD(359)(5) <= VNStageIntLLROutputS4xD(333)(5);
  CNStageIntLLRInputS5xD(40)(5) <= VNStageIntLLROutputS4xD(334)(0);
  CNStageIntLLRInputS5xD(66)(5) <= VNStageIntLLROutputS4xD(334)(1);
  CNStageIntLLRInputS5xD(217)(5) <= VNStageIntLLROutputS4xD(334)(2);
  CNStageIntLLRInputS5xD(286)(5) <= VNStageIntLLROutputS4xD(334)(3);
  CNStageIntLLRInputS5xD(380)(5) <= VNStageIntLLROutputS4xD(334)(4);
  CNStageIntLLRInputS5xD(39)(5) <= VNStageIntLLROutputS4xD(335)(0);
  CNStageIntLLRInputS5xD(78)(5) <= VNStageIntLLROutputS4xD(335)(1);
  CNStageIntLLRInputS5xD(170)(5) <= VNStageIntLLROutputS4xD(335)(2);
  CNStageIntLLRInputS5xD(189)(5) <= VNStageIntLLROutputS4xD(335)(3);
  CNStageIntLLRInputS5xD(274)(5) <= VNStageIntLLROutputS4xD(335)(4);
  CNStageIntLLRInputS5xD(291)(5) <= VNStageIntLLROutputS4xD(335)(5);
  CNStageIntLLRInputS5xD(343)(5) <= VNStageIntLLROutputS4xD(335)(6);
  CNStageIntLLRInputS5xD(38)(5) <= VNStageIntLLROutputS4xD(336)(0);
  CNStageIntLLRInputS5xD(104)(5) <= VNStageIntLLROutputS4xD(336)(1);
  CNStageIntLLRInputS5xD(121)(5) <= VNStageIntLLROutputS4xD(336)(2);
  CNStageIntLLRInputS5xD(267)(5) <= VNStageIntLLROutputS4xD(336)(3);
  CNStageIntLLRInputS5xD(332)(5) <= VNStageIntLLROutputS4xD(336)(4);
  CNStageIntLLRInputS5xD(344)(5) <= VNStageIntLLROutputS4xD(336)(5);
  CNStageIntLLRInputS5xD(37)(5) <= VNStageIntLLROutputS4xD(337)(0);
  CNStageIntLLRInputS5xD(93)(5) <= VNStageIntLLROutputS4xD(337)(1);
  CNStageIntLLRInputS5xD(115)(5) <= VNStageIntLLROutputS4xD(337)(2);
  CNStageIntLLRInputS5xD(183)(5) <= VNStageIntLLROutputS4xD(337)(3);
  CNStageIntLLRInputS5xD(253)(5) <= VNStageIntLLROutputS4xD(337)(4);
  CNStageIntLLRInputS5xD(290)(5) <= VNStageIntLLROutputS4xD(337)(5);
  CNStageIntLLRInputS5xD(379)(5) <= VNStageIntLLROutputS4xD(337)(6);
  CNStageIntLLRInputS5xD(36)(5) <= VNStageIntLLROutputS4xD(338)(0);
  CNStageIntLLRInputS5xD(80)(5) <= VNStageIntLLROutputS4xD(338)(1);
  CNStageIntLLRInputS5xD(155)(5) <= VNStageIntLLROutputS4xD(338)(2);
  CNStageIntLLRInputS5xD(190)(5) <= VNStageIntLLROutputS4xD(338)(3);
  CNStageIntLLRInputS5xD(370)(5) <= VNStageIntLLROutputS4xD(338)(4);
  CNStageIntLLRInputS5xD(35)(5) <= VNStageIntLLROutputS4xD(339)(0);
  CNStageIntLLRInputS5xD(96)(5) <= VNStageIntLLROutputS4xD(339)(1);
  CNStageIntLLRInputS5xD(163)(5) <= VNStageIntLLROutputS4xD(339)(2);
  CNStageIntLLRInputS5xD(216)(5) <= VNStageIntLLROutputS4xD(339)(3);
  CNStageIntLLRInputS5xD(247)(5) <= VNStageIntLLROutputS4xD(339)(4);
  CNStageIntLLRInputS5xD(322)(5) <= VNStageIntLLROutputS4xD(339)(5);
  CNStageIntLLRInputS5xD(34)(5) <= VNStageIntLLROutputS4xD(340)(0);
  CNStageIntLLRInputS5xD(58)(5) <= VNStageIntLLROutputS4xD(340)(1);
  CNStageIntLLRInputS5xD(127)(5) <= VNStageIntLLROutputS4xD(340)(2);
  CNStageIntLLRInputS5xD(178)(5) <= VNStageIntLLROutputS4xD(340)(3);
  CNStageIntLLRInputS5xD(245)(5) <= VNStageIntLLROutputS4xD(340)(4);
  CNStageIntLLRInputS5xD(334)(5) <= VNStageIntLLROutputS4xD(340)(5);
  CNStageIntLLRInputS5xD(33)(5) <= VNStageIntLLROutputS4xD(341)(0);
  CNStageIntLLRInputS5xD(68)(5) <= VNStageIntLLROutputS4xD(341)(1);
  CNStageIntLLRInputS5xD(125)(5) <= VNStageIntLLROutputS4xD(341)(2);
  CNStageIntLLRInputS5xD(204)(5) <= VNStageIntLLROutputS4xD(341)(3);
  CNStageIntLLRInputS5xD(258)(5) <= VNStageIntLLROutputS4xD(341)(4);
  CNStageIntLLRInputS5xD(296)(5) <= VNStageIntLLROutputS4xD(341)(5);
  CNStageIntLLRInputS5xD(32)(5) <= VNStageIntLLROutputS4xD(342)(0);
  CNStageIntLLRInputS5xD(63)(5) <= VNStageIntLLROutputS4xD(342)(1);
  CNStageIntLLRInputS5xD(161)(5) <= VNStageIntLLROutputS4xD(342)(2);
  CNStageIntLLRInputS5xD(251)(5) <= VNStageIntLLROutputS4xD(342)(3);
  CNStageIntLLRInputS5xD(294)(5) <= VNStageIntLLROutputS4xD(342)(4);
  CNStageIntLLRInputS5xD(31)(5) <= VNStageIntLLROutputS4xD(343)(0);
  CNStageIntLLRInputS5xD(69)(5) <= VNStageIntLLROutputS4xD(343)(1);
  CNStageIntLLRInputS5xD(140)(5) <= VNStageIntLLROutputS4xD(343)(2);
  CNStageIntLLRInputS5xD(206)(5) <= VNStageIntLLROutputS4xD(343)(3);
  CNStageIntLLRInputS5xD(228)(5) <= VNStageIntLLROutputS4xD(343)(4);
  CNStageIntLLRInputS5xD(327)(5) <= VNStageIntLLROutputS4xD(343)(5);
  CNStageIntLLRInputS5xD(30)(5) <= VNStageIntLLROutputS4xD(344)(0);
  CNStageIntLLRInputS5xD(57)(5) <= VNStageIntLLROutputS4xD(344)(1);
  CNStageIntLLRInputS5xD(143)(5) <= VNStageIntLLROutputS4xD(344)(2);
  CNStageIntLLRInputS5xD(218)(5) <= VNStageIntLLROutputS4xD(344)(3);
  CNStageIntLLRInputS5xD(238)(5) <= VNStageIntLLROutputS4xD(344)(4);
  CNStageIntLLRInputS5xD(307)(5) <= VNStageIntLLROutputS4xD(344)(5);
  CNStageIntLLRInputS5xD(367)(5) <= VNStageIntLLROutputS4xD(344)(6);
  CNStageIntLLRInputS5xD(29)(5) <= VNStageIntLLROutputS4xD(345)(0);
  CNStageIntLLRInputS5xD(83)(5) <= VNStageIntLLROutputS4xD(345)(1);
  CNStageIntLLRInputS5xD(128)(5) <= VNStageIntLLROutputS4xD(345)(2);
  CNStageIntLLRInputS5xD(232)(5) <= VNStageIntLLROutputS4xD(345)(3);
  CNStageIntLLRInputS5xD(309)(5) <= VNStageIntLLROutputS4xD(345)(4);
  CNStageIntLLRInputS5xD(375)(5) <= VNStageIntLLROutputS4xD(345)(5);
  CNStageIntLLRInputS5xD(28)(5) <= VNStageIntLLROutputS4xD(346)(0);
  CNStageIntLLRInputS5xD(89)(5) <= VNStageIntLLROutputS4xD(346)(1);
  CNStageIntLLRInputS5xD(162)(5) <= VNStageIntLLROutputS4xD(346)(2);
  CNStageIntLLRInputS5xD(181)(5) <= VNStageIntLLROutputS4xD(346)(3);
  CNStageIntLLRInputS5xD(235)(5) <= VNStageIntLLROutputS4xD(346)(4);
  CNStageIntLLRInputS5xD(297)(5) <= VNStageIntLLROutputS4xD(346)(5);
  CNStageIntLLRInputS5xD(339)(5) <= VNStageIntLLROutputS4xD(346)(6);
  CNStageIntLLRInputS5xD(27)(5) <= VNStageIntLLROutputS4xD(347)(0);
  CNStageIntLLRInputS5xD(73)(5) <= VNStageIntLLROutputS4xD(347)(1);
  CNStageIntLLRInputS5xD(124)(5) <= VNStageIntLLROutputS4xD(347)(2);
  CNStageIntLLRInputS5xD(199)(5) <= VNStageIntLLROutputS4xD(347)(3);
  CNStageIntLLRInputS5xD(225)(5) <= VNStageIntLLROutputS4xD(347)(4);
  CNStageIntLLRInputS5xD(328)(5) <= VNStageIntLLROutputS4xD(347)(5);
  CNStageIntLLRInputS5xD(337)(5) <= VNStageIntLLROutputS4xD(347)(6);
  CNStageIntLLRInputS5xD(26)(5) <= VNStageIntLLROutputS4xD(348)(0);
  CNStageIntLLRInputS5xD(75)(5) <= VNStageIntLLROutputS4xD(348)(1);
  CNStageIntLLRInputS5xD(152)(5) <= VNStageIntLLROutputS4xD(348)(2);
  CNStageIntLLRInputS5xD(200)(5) <= VNStageIntLLROutputS4xD(348)(3);
  CNStageIntLLRInputS5xD(259)(5) <= VNStageIntLLROutputS4xD(348)(4);
  CNStageIntLLRInputS5xD(293)(5) <= VNStageIntLLROutputS4xD(348)(5);
  CNStageIntLLRInputS5xD(373)(5) <= VNStageIntLLROutputS4xD(348)(6);
  CNStageIntLLRInputS5xD(25)(5) <= VNStageIntLLROutputS4xD(349)(0);
  CNStageIntLLRInputS5xD(99)(5) <= VNStageIntLLROutputS4xD(349)(1);
  CNStageIntLLRInputS5xD(180)(5) <= VNStageIntLLROutputS4xD(349)(2);
  CNStageIntLLRInputS5xD(244)(5) <= VNStageIntLLROutputS4xD(349)(3);
  CNStageIntLLRInputS5xD(319)(5) <= VNStageIntLLROutputS4xD(349)(4);
  CNStageIntLLRInputS5xD(352)(5) <= VNStageIntLLROutputS4xD(349)(5);
  CNStageIntLLRInputS5xD(24)(5) <= VNStageIntLLROutputS4xD(350)(0);
  CNStageIntLLRInputS5xD(81)(5) <= VNStageIntLLROutputS4xD(350)(1);
  CNStageIntLLRInputS5xD(164)(5) <= VNStageIntLLROutputS4xD(350)(2);
  CNStageIntLLRInputS5xD(171)(5) <= VNStageIntLLROutputS4xD(350)(3);
  CNStageIntLLRInputS5xD(254)(5) <= VNStageIntLLROutputS4xD(350)(4);
  CNStageIntLLRInputS5xD(303)(5) <= VNStageIntLLROutputS4xD(350)(5);
  CNStageIntLLRInputS5xD(23)(5) <= VNStageIntLLROutputS4xD(351)(0);
  CNStageIntLLRInputS5xD(154)(5) <= VNStageIntLLROutputS4xD(351)(1);
  CNStageIntLLRInputS5xD(188)(5) <= VNStageIntLLROutputS4xD(351)(2);
  CNStageIntLLRInputS5xD(266)(5) <= VNStageIntLLROutputS4xD(351)(3);
  CNStageIntLLRInputS5xD(329)(5) <= VNStageIntLLROutputS4xD(351)(4);
  CNStageIntLLRInputS5xD(340)(5) <= VNStageIntLLROutputS4xD(351)(5);
  CNStageIntLLRInputS5xD(22)(5) <= VNStageIntLLROutputS4xD(352)(0);
  CNStageIntLLRInputS5xD(100)(5) <= VNStageIntLLROutputS4xD(352)(1);
  CNStageIntLLRInputS5xD(141)(5) <= VNStageIntLLROutputS4xD(352)(2);
  CNStageIntLLRInputS5xD(192)(5) <= VNStageIntLLROutputS4xD(352)(3);
  CNStageIntLLRInputS5xD(239)(5) <= VNStageIntLLROutputS4xD(352)(4);
  CNStageIntLLRInputS5xD(321)(5) <= VNStageIntLLROutputS4xD(352)(5);
  CNStageIntLLRInputS5xD(374)(5) <= VNStageIntLLROutputS4xD(352)(6);
  CNStageIntLLRInputS5xD(21)(5) <= VNStageIntLLROutputS4xD(353)(0);
  CNStageIntLLRInputS5xD(74)(5) <= VNStageIntLLROutputS4xD(353)(1);
  CNStageIntLLRInputS5xD(160)(5) <= VNStageIntLLROutputS4xD(353)(2);
  CNStageIntLLRInputS5xD(224)(5) <= VNStageIntLLROutputS4xD(353)(3);
  CNStageIntLLRInputS5xD(227)(5) <= VNStageIntLLROutputS4xD(353)(4);
  CNStageIntLLRInputS5xD(336)(5) <= VNStageIntLLROutputS4xD(353)(5);
  CNStageIntLLRInputS5xD(20)(5) <= VNStageIntLLROutputS4xD(354)(0);
  CNStageIntLLRInputS5xD(88)(5) <= VNStageIntLLROutputS4xD(354)(1);
  CNStageIntLLRInputS5xD(133)(5) <= VNStageIntLLROutputS4xD(354)(2);
  CNStageIntLLRInputS5xD(191)(5) <= VNStageIntLLROutputS4xD(354)(3);
  CNStageIntLLRInputS5xD(326)(5) <= VNStageIntLLROutputS4xD(354)(4);
  CNStageIntLLRInputS5xD(364)(5) <= VNStageIntLLROutputS4xD(354)(5);
  CNStageIntLLRInputS5xD(19)(5) <= VNStageIntLLROutputS4xD(355)(0);
  CNStageIntLLRInputS5xD(59)(5) <= VNStageIntLLROutputS4xD(355)(1);
  CNStageIntLLRInputS5xD(130)(5) <= VNStageIntLLROutputS4xD(355)(2);
  CNStageIntLLRInputS5xD(186)(5) <= VNStageIntLLROutputS4xD(355)(3);
  CNStageIntLLRInputS5xD(230)(5) <= VNStageIntLLROutputS4xD(355)(4);
  CNStageIntLLRInputS5xD(300)(5) <= VNStageIntLLROutputS4xD(355)(5);
  CNStageIntLLRInputS5xD(349)(5) <= VNStageIntLLROutputS4xD(355)(6);
  CNStageIntLLRInputS5xD(18)(5) <= VNStageIntLLROutputS4xD(356)(0);
  CNStageIntLLRInputS5xD(95)(5) <= VNStageIntLLROutputS4xD(356)(1);
  CNStageIntLLRInputS5xD(146)(5) <= VNStageIntLLROutputS4xD(356)(2);
  CNStageIntLLRInputS5xD(222)(5) <= VNStageIntLLROutputS4xD(356)(3);
  CNStageIntLLRInputS5xD(299)(5) <= VNStageIntLLROutputS4xD(356)(4);
  CNStageIntLLRInputS5xD(376)(5) <= VNStageIntLLROutputS4xD(356)(5);
  CNStageIntLLRInputS5xD(17)(5) <= VNStageIntLLROutputS4xD(357)(0);
  CNStageIntLLRInputS5xD(61)(5) <= VNStageIntLLROutputS4xD(357)(1);
  CNStageIntLLRInputS5xD(138)(5) <= VNStageIntLLROutputS4xD(357)(2);
  CNStageIntLLRInputS5xD(176)(5) <= VNStageIntLLROutputS4xD(357)(3);
  CNStageIntLLRInputS5xD(256)(5) <= VNStageIntLLROutputS4xD(357)(4);
  CNStageIntLLRInputS5xD(312)(5) <= VNStageIntLLROutputS4xD(357)(5);
  CNStageIntLLRInputS5xD(366)(5) <= VNStageIntLLROutputS4xD(357)(6);
  CNStageIntLLRInputS5xD(16)(5) <= VNStageIntLLROutputS4xD(358)(0);
  CNStageIntLLRInputS5xD(76)(5) <= VNStageIntLLROutputS4xD(358)(1);
  CNStageIntLLRInputS5xD(112)(5) <= VNStageIntLLROutputS4xD(358)(2);
  CNStageIntLLRInputS5xD(252)(5) <= VNStageIntLLROutputS4xD(358)(3);
  CNStageIntLLRInputS5xD(305)(5) <= VNStageIntLLROutputS4xD(358)(4);
  CNStageIntLLRInputS5xD(353)(5) <= VNStageIntLLROutputS4xD(358)(5);
  CNStageIntLLRInputS5xD(15)(5) <= VNStageIntLLROutputS4xD(359)(0);
  CNStageIntLLRInputS5xD(72)(5) <= VNStageIntLLROutputS4xD(359)(1);
  CNStageIntLLRInputS5xD(122)(5) <= VNStageIntLLROutputS4xD(359)(2);
  CNStageIntLLRInputS5xD(195)(5) <= VNStageIntLLROutputS4xD(359)(3);
  CNStageIntLLRInputS5xD(257)(5) <= VNStageIntLLROutputS4xD(359)(4);
  CNStageIntLLRInputS5xD(283)(5) <= VNStageIntLLROutputS4xD(359)(5);
  CNStageIntLLRInputS5xD(372)(5) <= VNStageIntLLROutputS4xD(359)(6);
  CNStageIntLLRInputS5xD(14)(5) <= VNStageIntLLROutputS4xD(360)(0);
  CNStageIntLLRInputS5xD(91)(5) <= VNStageIntLLROutputS4xD(360)(1);
  CNStageIntLLRInputS5xD(116)(5) <= VNStageIntLLROutputS4xD(360)(2);
  CNStageIntLLRInputS5xD(174)(5) <= VNStageIntLLROutputS4xD(360)(3);
  CNStageIntLLRInputS5xD(248)(5) <= VNStageIntLLROutputS4xD(360)(4);
  CNStageIntLLRInputS5xD(292)(5) <= VNStageIntLLROutputS4xD(360)(5);
  CNStageIntLLRInputS5xD(345)(5) <= VNStageIntLLROutputS4xD(360)(6);
  CNStageIntLLRInputS5xD(13)(5) <= VNStageIntLLROutputS4xD(361)(0);
  CNStageIntLLRInputS5xD(54)(5) <= VNStageIntLLROutputS4xD(361)(1);
  CNStageIntLLRInputS5xD(120)(5) <= VNStageIntLLROutputS4xD(361)(2);
  CNStageIntLLRInputS5xD(207)(5) <= VNStageIntLLROutputS4xD(361)(3);
  CNStageIntLLRInputS5xD(271)(5) <= VNStageIntLLROutputS4xD(361)(4);
  CNStageIntLLRInputS5xD(285)(5) <= VNStageIntLLROutputS4xD(361)(5);
  CNStageIntLLRInputS5xD(342)(5) <= VNStageIntLLROutputS4xD(361)(6);
  CNStageIntLLRInputS5xD(12)(5) <= VNStageIntLLROutputS4xD(362)(0);
  CNStageIntLLRInputS5xD(55)(5) <= VNStageIntLLROutputS4xD(362)(1);
  CNStageIntLLRInputS5xD(169)(5) <= VNStageIntLLROutputS4xD(362)(2);
  CNStageIntLLRInputS5xD(210)(5) <= VNStageIntLLROutputS4xD(362)(3);
  CNStageIntLLRInputS5xD(276)(5) <= VNStageIntLLROutputS4xD(362)(4);
  CNStageIntLLRInputS5xD(289)(5) <= VNStageIntLLROutputS4xD(362)(5);
  CNStageIntLLRInputS5xD(357)(5) <= VNStageIntLLROutputS4xD(362)(6);
  CNStageIntLLRInputS5xD(90)(5) <= VNStageIntLLROutputS4xD(363)(0);
  CNStageIntLLRInputS5xD(147)(5) <= VNStageIntLLROutputS4xD(363)(1);
  CNStageIntLLRInputS5xD(197)(5) <= VNStageIntLLROutputS4xD(363)(2);
  CNStageIntLLRInputS5xD(261)(5) <= VNStageIntLLROutputS4xD(363)(3);
  CNStageIntLLRInputS5xD(281)(5) <= VNStageIntLLROutputS4xD(363)(4);
  CNStageIntLLRInputS5xD(11)(5) <= VNStageIntLLROutputS4xD(364)(0);
  CNStageIntLLRInputS5xD(82)(5) <= VNStageIntLLROutputS4xD(364)(1);
  CNStageIntLLRInputS5xD(129)(5) <= VNStageIntLLROutputS4xD(364)(2);
  CNStageIntLLRInputS5xD(175)(5) <= VNStageIntLLROutputS4xD(364)(3);
  CNStageIntLLRInputS5xD(263)(5) <= VNStageIntLLROutputS4xD(364)(4);
  CNStageIntLLRInputS5xD(313)(5) <= VNStageIntLLROutputS4xD(364)(5);
  CNStageIntLLRInputS5xD(10)(5) <= VNStageIntLLROutputS4xD(365)(0);
  CNStageIntLLRInputS5xD(98)(5) <= VNStageIntLLROutputS4xD(365)(1);
  CNStageIntLLRInputS5xD(142)(5) <= VNStageIntLLROutputS4xD(365)(2);
  CNStageIntLLRInputS5xD(194)(5) <= VNStageIntLLROutputS4xD(365)(3);
  CNStageIntLLRInputS5xD(234)(5) <= VNStageIntLLROutputS4xD(365)(4);
  CNStageIntLLRInputS5xD(298)(5) <= VNStageIntLLROutputS4xD(365)(5);
  CNStageIntLLRInputS5xD(9)(5) <= VNStageIntLLROutputS4xD(366)(0);
  CNStageIntLLRInputS5xD(102)(5) <= VNStageIntLLROutputS4xD(366)(1);
  CNStageIntLLRInputS5xD(153)(5) <= VNStageIntLLROutputS4xD(366)(2);
  CNStageIntLLRInputS5xD(219)(5) <= VNStageIntLLROutputS4xD(366)(3);
  CNStageIntLLRInputS5xD(269)(5) <= VNStageIntLLROutputS4xD(366)(4);
  CNStageIntLLRInputS5xD(308)(5) <= VNStageIntLLROutputS4xD(366)(5);
  CNStageIntLLRInputS5xD(8)(5) <= VNStageIntLLROutputS4xD(367)(0);
  CNStageIntLLRInputS5xD(110)(5) <= VNStageIntLLROutputS4xD(367)(1);
  CNStageIntLLRInputS5xD(123)(5) <= VNStageIntLLROutputS4xD(367)(2);
  CNStageIntLLRInputS5xD(205)(5) <= VNStageIntLLROutputS4xD(367)(3);
  CNStageIntLLRInputS5xD(226)(5) <= VNStageIntLLROutputS4xD(367)(4);
  CNStageIntLLRInputS5xD(320)(5) <= VNStageIntLLROutputS4xD(367)(5);
  CNStageIntLLRInputS5xD(333)(5) <= VNStageIntLLROutputS4xD(367)(6);
  CNStageIntLLRInputS5xD(7)(5) <= VNStageIntLLROutputS4xD(368)(0);
  CNStageIntLLRInputS5xD(177)(5) <= VNStageIntLLROutputS4xD(368)(1);
  CNStageIntLLRInputS5xD(381)(5) <= VNStageIntLLROutputS4xD(368)(2);
  CNStageIntLLRInputS5xD(6)(5) <= VNStageIntLLROutputS4xD(369)(0);
  CNStageIntLLRInputS5xD(156)(5) <= VNStageIntLLROutputS4xD(369)(1);
  CNStageIntLLRInputS5xD(221)(5) <= VNStageIntLLROutputS4xD(369)(2);
  CNStageIntLLRInputS5xD(262)(5) <= VNStageIntLLROutputS4xD(369)(3);
  CNStageIntLLRInputS5xD(358)(5) <= VNStageIntLLROutputS4xD(369)(4);
  CNStageIntLLRInputS5xD(5)(5) <= VNStageIntLLROutputS4xD(370)(0);
  CNStageIntLLRInputS5xD(114)(5) <= VNStageIntLLROutputS4xD(370)(1);
  CNStageIntLLRInputS5xD(208)(5) <= VNStageIntLLROutputS4xD(370)(2);
  CNStageIntLLRInputS5xD(275)(5) <= VNStageIntLLROutputS4xD(370)(3);
  CNStageIntLLRInputS5xD(341)(5) <= VNStageIntLLROutputS4xD(370)(4);
  CNStageIntLLRInputS5xD(4)(5) <= VNStageIntLLROutputS4xD(371)(0);
  CNStageIntLLRInputS5xD(135)(5) <= VNStageIntLLROutputS4xD(371)(1);
  CNStageIntLLRInputS5xD(173)(5) <= VNStageIntLLROutputS4xD(371)(2);
  CNStageIntLLRInputS5xD(249)(5) <= VNStageIntLLROutputS4xD(371)(3);
  CNStageIntLLRInputS5xD(354)(5) <= VNStageIntLLROutputS4xD(371)(4);
  CNStageIntLLRInputS5xD(106)(5) <= VNStageIntLLROutputS4xD(372)(0);
  CNStageIntLLRInputS5xD(144)(5) <= VNStageIntLLROutputS4xD(372)(1);
  CNStageIntLLRInputS5xD(201)(5) <= VNStageIntLLROutputS4xD(372)(2);
  CNStageIntLLRInputS5xD(229)(5) <= VNStageIntLLROutputS4xD(372)(3);
  CNStageIntLLRInputS5xD(301)(5) <= VNStageIntLLROutputS4xD(372)(4);
  CNStageIntLLRInputS5xD(365)(5) <= VNStageIntLLROutputS4xD(372)(5);
  CNStageIntLLRInputS5xD(3)(5) <= VNStageIntLLROutputS4xD(373)(0);
  CNStageIntLLRInputS5xD(139)(5) <= VNStageIntLLROutputS4xD(373)(1);
  CNStageIntLLRInputS5xD(250)(5) <= VNStageIntLLROutputS4xD(373)(2);
  CNStageIntLLRInputS5xD(310)(5) <= VNStageIntLLROutputS4xD(373)(3);
  CNStageIntLLRInputS5xD(335)(5) <= VNStageIntLLROutputS4xD(373)(4);
  CNStageIntLLRInputS5xD(2)(5) <= VNStageIntLLROutputS4xD(374)(0);
  CNStageIntLLRInputS5xD(85)(5) <= VNStageIntLLROutputS4xD(374)(1);
  CNStageIntLLRInputS5xD(145)(5) <= VNStageIntLLROutputS4xD(374)(2);
  CNStageIntLLRInputS5xD(213)(5) <= VNStageIntLLROutputS4xD(374)(3);
  CNStageIntLLRInputS5xD(264)(5) <= VNStageIntLLROutputS4xD(374)(4);
  CNStageIntLLRInputS5xD(306)(5) <= VNStageIntLLROutputS4xD(374)(5);
  CNStageIntLLRInputS5xD(383)(5) <= VNStageIntLLROutputS4xD(374)(6);
  CNStageIntLLRInputS5xD(1)(5) <= VNStageIntLLROutputS4xD(375)(0);
  CNStageIntLLRInputS5xD(64)(5) <= VNStageIntLLROutputS4xD(375)(1);
  CNStageIntLLRInputS5xD(134)(5) <= VNStageIntLLROutputS4xD(375)(2);
  CNStageIntLLRInputS5xD(260)(5) <= VNStageIntLLROutputS4xD(375)(3);
  CNStageIntLLRInputS5xD(311)(5) <= VNStageIntLLROutputS4xD(375)(4);
  CNStageIntLLRInputS5xD(368)(5) <= VNStageIntLLROutputS4xD(375)(5);
  CNStageIntLLRInputS5xD(0)(5) <= VNStageIntLLROutputS4xD(376)(0);
  CNStageIntLLRInputS5xD(67)(5) <= VNStageIntLLROutputS4xD(376)(1);
  CNStageIntLLRInputS5xD(159)(5) <= VNStageIntLLROutputS4xD(376)(2);
  CNStageIntLLRInputS5xD(278)(5) <= VNStageIntLLROutputS4xD(376)(3);
  CNStageIntLLRInputS5xD(107)(5) <= VNStageIntLLROutputS4xD(377)(0);
  CNStageIntLLRInputS5xD(166)(5) <= VNStageIntLLROutputS4xD(377)(1);
  CNStageIntLLRInputS5xD(193)(5) <= VNStageIntLLROutputS4xD(377)(2);
  CNStageIntLLRInputS5xD(325)(5) <= VNStageIntLLROutputS4xD(377)(3);
  CNStageIntLLRInputS5xD(347)(5) <= VNStageIntLLROutputS4xD(377)(4);
  CNStageIntLLRInputS5xD(86)(5) <= VNStageIntLLROutputS4xD(378)(0);
  CNStageIntLLRInputS5xD(149)(5) <= VNStageIntLLROutputS4xD(378)(1);
  CNStageIntLLRInputS5xD(187)(5) <= VNStageIntLLROutputS4xD(378)(2);
  CNStageIntLLRInputS5xD(246)(5) <= VNStageIntLLROutputS4xD(378)(3);
  CNStageIntLLRInputS5xD(331)(5) <= VNStageIntLLROutputS4xD(378)(4);
  CNStageIntLLRInputS5xD(355)(5) <= VNStageIntLLROutputS4xD(378)(5);
  CNStageIntLLRInputS5xD(105)(5) <= VNStageIntLLROutputS4xD(379)(0);
  CNStageIntLLRInputS5xD(151)(5) <= VNStageIntLLROutputS4xD(379)(1);
  CNStageIntLLRInputS5xD(277)(5) <= VNStageIntLLROutputS4xD(379)(2);
  CNStageIntLLRInputS5xD(315)(5) <= VNStageIntLLROutputS4xD(379)(3);
  CNStageIntLLRInputS5xD(351)(5) <= VNStageIntLLROutputS4xD(379)(4);
  CNStageIntLLRInputS5xD(77)(5) <= VNStageIntLLROutputS4xD(380)(0);
  CNStageIntLLRInputS5xD(118)(5) <= VNStageIntLLROutputS4xD(380)(1);
  CNStageIntLLRInputS5xD(182)(5) <= VNStageIntLLROutputS4xD(380)(2);
  CNStageIntLLRInputS5xD(270)(5) <= VNStageIntLLROutputS4xD(380)(3);
  CNStageIntLLRInputS5xD(317)(5) <= VNStageIntLLROutputS4xD(380)(4);
  CNStageIntLLRInputS5xD(356)(5) <= VNStageIntLLROutputS4xD(380)(5);
  CNStageIntLLRInputS5xD(60)(5) <= VNStageIntLLROutputS4xD(381)(0);
  CNStageIntLLRInputS5xD(157)(5) <= VNStageIntLLROutputS4xD(381)(1);
  CNStageIntLLRInputS5xD(214)(5) <= VNStageIntLLROutputS4xD(381)(2);
  CNStageIntLLRInputS5xD(233)(5) <= VNStageIntLLROutputS4xD(381)(3);
  CNStageIntLLRInputS5xD(287)(5) <= VNStageIntLLROutputS4xD(381)(4);
  CNStageIntLLRInputS5xD(346)(5) <= VNStageIntLLROutputS4xD(381)(5);
  CNStageIntLLRInputS5xD(87)(5) <= VNStageIntLLROutputS4xD(382)(0);
  CNStageIntLLRInputS5xD(111)(5) <= VNStageIntLLROutputS4xD(382)(1);
  CNStageIntLLRInputS5xD(198)(5) <= VNStageIntLLROutputS4xD(382)(2);
  CNStageIntLLRInputS5xD(237)(5) <= VNStageIntLLROutputS4xD(382)(3);
  CNStageIntLLRInputS5xD(323)(5) <= VNStageIntLLROutputS4xD(382)(4);
  CNStageIntLLRInputS5xD(371)(5) <= VNStageIntLLROutputS4xD(382)(5);
  CNStageIntLLRInputS5xD(52)(5) <= VNStageIntLLROutputS4xD(383)(0);
  CNStageIntLLRInputS5xD(79)(5) <= VNStageIntLLROutputS4xD(383)(1);
  CNStageIntLLRInputS5xD(119)(5) <= VNStageIntLLROutputS4xD(383)(2);
  CNStageIntLLRInputS5xD(209)(5) <= VNStageIntLLROutputS4xD(383)(3);
  CNStageIntLLRInputS5xD(279)(5) <= VNStageIntLLROutputS4xD(383)(4);
  CNStageIntLLRInputS5xD(282)(5) <= VNStageIntLLROutputS4xD(383)(5);
  CNStageIntLLRInputS5xD(378)(5) <= VNStageIntLLROutputS4xD(383)(6);

  -- Variable Nodes (Iteration 5)
  VNStageIntLLRInputS5xD(56)(0) <= CNStageIntLLROutputS5xD(0)(0);
  VNStageIntLLRInputS5xD(120)(0) <= CNStageIntLLROutputS5xD(0)(1);
  VNStageIntLLRInputS5xD(184)(0) <= CNStageIntLLROutputS5xD(0)(2);
  VNStageIntLLRInputS5xD(248)(0) <= CNStageIntLLROutputS5xD(0)(3);
  VNStageIntLLRInputS5xD(312)(0) <= CNStageIntLLROutputS5xD(0)(4);
  VNStageIntLLRInputS5xD(376)(0) <= CNStageIntLLROutputS5xD(0)(5);
  VNStageIntLLRInputS5xD(55)(0) <= CNStageIntLLROutputS5xD(1)(0);
  VNStageIntLLRInputS5xD(119)(0) <= CNStageIntLLROutputS5xD(1)(1);
  VNStageIntLLRInputS5xD(183)(0) <= CNStageIntLLROutputS5xD(1)(2);
  VNStageIntLLRInputS5xD(247)(0) <= CNStageIntLLROutputS5xD(1)(3);
  VNStageIntLLRInputS5xD(311)(0) <= CNStageIntLLROutputS5xD(1)(4);
  VNStageIntLLRInputS5xD(375)(0) <= CNStageIntLLROutputS5xD(1)(5);
  VNStageIntLLRInputS5xD(54)(0) <= CNStageIntLLROutputS5xD(2)(0);
  VNStageIntLLRInputS5xD(118)(0) <= CNStageIntLLROutputS5xD(2)(1);
  VNStageIntLLRInputS5xD(182)(0) <= CNStageIntLLROutputS5xD(2)(2);
  VNStageIntLLRInputS5xD(246)(0) <= CNStageIntLLROutputS5xD(2)(3);
  VNStageIntLLRInputS5xD(310)(0) <= CNStageIntLLROutputS5xD(2)(4);
  VNStageIntLLRInputS5xD(374)(0) <= CNStageIntLLROutputS5xD(2)(5);
  VNStageIntLLRInputS5xD(53)(0) <= CNStageIntLLROutputS5xD(3)(0);
  VNStageIntLLRInputS5xD(117)(0) <= CNStageIntLLROutputS5xD(3)(1);
  VNStageIntLLRInputS5xD(181)(0) <= CNStageIntLLROutputS5xD(3)(2);
  VNStageIntLLRInputS5xD(245)(0) <= CNStageIntLLROutputS5xD(3)(3);
  VNStageIntLLRInputS5xD(309)(0) <= CNStageIntLLROutputS5xD(3)(4);
  VNStageIntLLRInputS5xD(373)(0) <= CNStageIntLLROutputS5xD(3)(5);
  VNStageIntLLRInputS5xD(51)(0) <= CNStageIntLLROutputS5xD(4)(0);
  VNStageIntLLRInputS5xD(115)(0) <= CNStageIntLLROutputS5xD(4)(1);
  VNStageIntLLRInputS5xD(179)(0) <= CNStageIntLLROutputS5xD(4)(2);
  VNStageIntLLRInputS5xD(243)(0) <= CNStageIntLLROutputS5xD(4)(3);
  VNStageIntLLRInputS5xD(307)(0) <= CNStageIntLLROutputS5xD(4)(4);
  VNStageIntLLRInputS5xD(371)(0) <= CNStageIntLLROutputS5xD(4)(5);
  VNStageIntLLRInputS5xD(50)(0) <= CNStageIntLLROutputS5xD(5)(0);
  VNStageIntLLRInputS5xD(114)(0) <= CNStageIntLLROutputS5xD(5)(1);
  VNStageIntLLRInputS5xD(178)(0) <= CNStageIntLLROutputS5xD(5)(2);
  VNStageIntLLRInputS5xD(242)(0) <= CNStageIntLLROutputS5xD(5)(3);
  VNStageIntLLRInputS5xD(306)(0) <= CNStageIntLLROutputS5xD(5)(4);
  VNStageIntLLRInputS5xD(370)(0) <= CNStageIntLLROutputS5xD(5)(5);
  VNStageIntLLRInputS5xD(49)(0) <= CNStageIntLLROutputS5xD(6)(0);
  VNStageIntLLRInputS5xD(113)(0) <= CNStageIntLLROutputS5xD(6)(1);
  VNStageIntLLRInputS5xD(177)(0) <= CNStageIntLLROutputS5xD(6)(2);
  VNStageIntLLRInputS5xD(241)(0) <= CNStageIntLLROutputS5xD(6)(3);
  VNStageIntLLRInputS5xD(305)(0) <= CNStageIntLLROutputS5xD(6)(4);
  VNStageIntLLRInputS5xD(369)(0) <= CNStageIntLLROutputS5xD(6)(5);
  VNStageIntLLRInputS5xD(48)(0) <= CNStageIntLLROutputS5xD(7)(0);
  VNStageIntLLRInputS5xD(112)(0) <= CNStageIntLLROutputS5xD(7)(1);
  VNStageIntLLRInputS5xD(176)(0) <= CNStageIntLLROutputS5xD(7)(2);
  VNStageIntLLRInputS5xD(240)(0) <= CNStageIntLLROutputS5xD(7)(3);
  VNStageIntLLRInputS5xD(304)(0) <= CNStageIntLLROutputS5xD(7)(4);
  VNStageIntLLRInputS5xD(368)(0) <= CNStageIntLLROutputS5xD(7)(5);
  VNStageIntLLRInputS5xD(47)(0) <= CNStageIntLLROutputS5xD(8)(0);
  VNStageIntLLRInputS5xD(111)(0) <= CNStageIntLLROutputS5xD(8)(1);
  VNStageIntLLRInputS5xD(175)(0) <= CNStageIntLLROutputS5xD(8)(2);
  VNStageIntLLRInputS5xD(239)(0) <= CNStageIntLLROutputS5xD(8)(3);
  VNStageIntLLRInputS5xD(303)(0) <= CNStageIntLLROutputS5xD(8)(4);
  VNStageIntLLRInputS5xD(367)(0) <= CNStageIntLLROutputS5xD(8)(5);
  VNStageIntLLRInputS5xD(46)(0) <= CNStageIntLLROutputS5xD(9)(0);
  VNStageIntLLRInputS5xD(110)(0) <= CNStageIntLLROutputS5xD(9)(1);
  VNStageIntLLRInputS5xD(174)(0) <= CNStageIntLLROutputS5xD(9)(2);
  VNStageIntLLRInputS5xD(238)(0) <= CNStageIntLLROutputS5xD(9)(3);
  VNStageIntLLRInputS5xD(302)(0) <= CNStageIntLLROutputS5xD(9)(4);
  VNStageIntLLRInputS5xD(366)(0) <= CNStageIntLLROutputS5xD(9)(5);
  VNStageIntLLRInputS5xD(45)(0) <= CNStageIntLLROutputS5xD(10)(0);
  VNStageIntLLRInputS5xD(109)(0) <= CNStageIntLLROutputS5xD(10)(1);
  VNStageIntLLRInputS5xD(173)(0) <= CNStageIntLLROutputS5xD(10)(2);
  VNStageIntLLRInputS5xD(237)(0) <= CNStageIntLLROutputS5xD(10)(3);
  VNStageIntLLRInputS5xD(301)(0) <= CNStageIntLLROutputS5xD(10)(4);
  VNStageIntLLRInputS5xD(365)(0) <= CNStageIntLLROutputS5xD(10)(5);
  VNStageIntLLRInputS5xD(44)(0) <= CNStageIntLLROutputS5xD(11)(0);
  VNStageIntLLRInputS5xD(108)(0) <= CNStageIntLLROutputS5xD(11)(1);
  VNStageIntLLRInputS5xD(172)(0) <= CNStageIntLLROutputS5xD(11)(2);
  VNStageIntLLRInputS5xD(236)(0) <= CNStageIntLLROutputS5xD(11)(3);
  VNStageIntLLRInputS5xD(300)(0) <= CNStageIntLLROutputS5xD(11)(4);
  VNStageIntLLRInputS5xD(364)(0) <= CNStageIntLLROutputS5xD(11)(5);
  VNStageIntLLRInputS5xD(42)(0) <= CNStageIntLLROutputS5xD(12)(0);
  VNStageIntLLRInputS5xD(106)(0) <= CNStageIntLLROutputS5xD(12)(1);
  VNStageIntLLRInputS5xD(170)(0) <= CNStageIntLLROutputS5xD(12)(2);
  VNStageIntLLRInputS5xD(234)(0) <= CNStageIntLLROutputS5xD(12)(3);
  VNStageIntLLRInputS5xD(298)(0) <= CNStageIntLLROutputS5xD(12)(4);
  VNStageIntLLRInputS5xD(362)(0) <= CNStageIntLLROutputS5xD(12)(5);
  VNStageIntLLRInputS5xD(41)(0) <= CNStageIntLLROutputS5xD(13)(0);
  VNStageIntLLRInputS5xD(105)(0) <= CNStageIntLLROutputS5xD(13)(1);
  VNStageIntLLRInputS5xD(169)(0) <= CNStageIntLLROutputS5xD(13)(2);
  VNStageIntLLRInputS5xD(233)(0) <= CNStageIntLLROutputS5xD(13)(3);
  VNStageIntLLRInputS5xD(297)(0) <= CNStageIntLLROutputS5xD(13)(4);
  VNStageIntLLRInputS5xD(361)(0) <= CNStageIntLLROutputS5xD(13)(5);
  VNStageIntLLRInputS5xD(40)(0) <= CNStageIntLLROutputS5xD(14)(0);
  VNStageIntLLRInputS5xD(104)(0) <= CNStageIntLLROutputS5xD(14)(1);
  VNStageIntLLRInputS5xD(168)(0) <= CNStageIntLLROutputS5xD(14)(2);
  VNStageIntLLRInputS5xD(232)(0) <= CNStageIntLLROutputS5xD(14)(3);
  VNStageIntLLRInputS5xD(296)(0) <= CNStageIntLLROutputS5xD(14)(4);
  VNStageIntLLRInputS5xD(360)(0) <= CNStageIntLLROutputS5xD(14)(5);
  VNStageIntLLRInputS5xD(39)(0) <= CNStageIntLLROutputS5xD(15)(0);
  VNStageIntLLRInputS5xD(103)(0) <= CNStageIntLLROutputS5xD(15)(1);
  VNStageIntLLRInputS5xD(167)(0) <= CNStageIntLLROutputS5xD(15)(2);
  VNStageIntLLRInputS5xD(231)(0) <= CNStageIntLLROutputS5xD(15)(3);
  VNStageIntLLRInputS5xD(295)(0) <= CNStageIntLLROutputS5xD(15)(4);
  VNStageIntLLRInputS5xD(359)(0) <= CNStageIntLLROutputS5xD(15)(5);
  VNStageIntLLRInputS5xD(38)(0) <= CNStageIntLLROutputS5xD(16)(0);
  VNStageIntLLRInputS5xD(102)(0) <= CNStageIntLLROutputS5xD(16)(1);
  VNStageIntLLRInputS5xD(166)(0) <= CNStageIntLLROutputS5xD(16)(2);
  VNStageIntLLRInputS5xD(230)(0) <= CNStageIntLLROutputS5xD(16)(3);
  VNStageIntLLRInputS5xD(294)(0) <= CNStageIntLLROutputS5xD(16)(4);
  VNStageIntLLRInputS5xD(358)(0) <= CNStageIntLLROutputS5xD(16)(5);
  VNStageIntLLRInputS5xD(37)(0) <= CNStageIntLLROutputS5xD(17)(0);
  VNStageIntLLRInputS5xD(101)(0) <= CNStageIntLLROutputS5xD(17)(1);
  VNStageIntLLRInputS5xD(165)(0) <= CNStageIntLLROutputS5xD(17)(2);
  VNStageIntLLRInputS5xD(229)(0) <= CNStageIntLLROutputS5xD(17)(3);
  VNStageIntLLRInputS5xD(293)(0) <= CNStageIntLLROutputS5xD(17)(4);
  VNStageIntLLRInputS5xD(357)(0) <= CNStageIntLLROutputS5xD(17)(5);
  VNStageIntLLRInputS5xD(36)(0) <= CNStageIntLLROutputS5xD(18)(0);
  VNStageIntLLRInputS5xD(100)(0) <= CNStageIntLLROutputS5xD(18)(1);
  VNStageIntLLRInputS5xD(164)(0) <= CNStageIntLLROutputS5xD(18)(2);
  VNStageIntLLRInputS5xD(228)(0) <= CNStageIntLLROutputS5xD(18)(3);
  VNStageIntLLRInputS5xD(292)(0) <= CNStageIntLLROutputS5xD(18)(4);
  VNStageIntLLRInputS5xD(356)(0) <= CNStageIntLLROutputS5xD(18)(5);
  VNStageIntLLRInputS5xD(35)(0) <= CNStageIntLLROutputS5xD(19)(0);
  VNStageIntLLRInputS5xD(99)(0) <= CNStageIntLLROutputS5xD(19)(1);
  VNStageIntLLRInputS5xD(163)(0) <= CNStageIntLLROutputS5xD(19)(2);
  VNStageIntLLRInputS5xD(227)(0) <= CNStageIntLLROutputS5xD(19)(3);
  VNStageIntLLRInputS5xD(291)(0) <= CNStageIntLLROutputS5xD(19)(4);
  VNStageIntLLRInputS5xD(355)(0) <= CNStageIntLLROutputS5xD(19)(5);
  VNStageIntLLRInputS5xD(34)(0) <= CNStageIntLLROutputS5xD(20)(0);
  VNStageIntLLRInputS5xD(98)(0) <= CNStageIntLLROutputS5xD(20)(1);
  VNStageIntLLRInputS5xD(162)(0) <= CNStageIntLLROutputS5xD(20)(2);
  VNStageIntLLRInputS5xD(226)(0) <= CNStageIntLLROutputS5xD(20)(3);
  VNStageIntLLRInputS5xD(290)(0) <= CNStageIntLLROutputS5xD(20)(4);
  VNStageIntLLRInputS5xD(354)(0) <= CNStageIntLLROutputS5xD(20)(5);
  VNStageIntLLRInputS5xD(33)(0) <= CNStageIntLLROutputS5xD(21)(0);
  VNStageIntLLRInputS5xD(97)(0) <= CNStageIntLLROutputS5xD(21)(1);
  VNStageIntLLRInputS5xD(161)(0) <= CNStageIntLLROutputS5xD(21)(2);
  VNStageIntLLRInputS5xD(225)(0) <= CNStageIntLLROutputS5xD(21)(3);
  VNStageIntLLRInputS5xD(289)(0) <= CNStageIntLLROutputS5xD(21)(4);
  VNStageIntLLRInputS5xD(353)(0) <= CNStageIntLLROutputS5xD(21)(5);
  VNStageIntLLRInputS5xD(32)(0) <= CNStageIntLLROutputS5xD(22)(0);
  VNStageIntLLRInputS5xD(96)(0) <= CNStageIntLLROutputS5xD(22)(1);
  VNStageIntLLRInputS5xD(160)(0) <= CNStageIntLLROutputS5xD(22)(2);
  VNStageIntLLRInputS5xD(224)(0) <= CNStageIntLLROutputS5xD(22)(3);
  VNStageIntLLRInputS5xD(288)(0) <= CNStageIntLLROutputS5xD(22)(4);
  VNStageIntLLRInputS5xD(352)(0) <= CNStageIntLLROutputS5xD(22)(5);
  VNStageIntLLRInputS5xD(31)(0) <= CNStageIntLLROutputS5xD(23)(0);
  VNStageIntLLRInputS5xD(95)(0) <= CNStageIntLLROutputS5xD(23)(1);
  VNStageIntLLRInputS5xD(159)(0) <= CNStageIntLLROutputS5xD(23)(2);
  VNStageIntLLRInputS5xD(223)(0) <= CNStageIntLLROutputS5xD(23)(3);
  VNStageIntLLRInputS5xD(287)(0) <= CNStageIntLLROutputS5xD(23)(4);
  VNStageIntLLRInputS5xD(351)(0) <= CNStageIntLLROutputS5xD(23)(5);
  VNStageIntLLRInputS5xD(30)(0) <= CNStageIntLLROutputS5xD(24)(0);
  VNStageIntLLRInputS5xD(94)(0) <= CNStageIntLLROutputS5xD(24)(1);
  VNStageIntLLRInputS5xD(158)(0) <= CNStageIntLLROutputS5xD(24)(2);
  VNStageIntLLRInputS5xD(222)(0) <= CNStageIntLLROutputS5xD(24)(3);
  VNStageIntLLRInputS5xD(286)(0) <= CNStageIntLLROutputS5xD(24)(4);
  VNStageIntLLRInputS5xD(350)(0) <= CNStageIntLLROutputS5xD(24)(5);
  VNStageIntLLRInputS5xD(29)(0) <= CNStageIntLLROutputS5xD(25)(0);
  VNStageIntLLRInputS5xD(93)(0) <= CNStageIntLLROutputS5xD(25)(1);
  VNStageIntLLRInputS5xD(157)(0) <= CNStageIntLLROutputS5xD(25)(2);
  VNStageIntLLRInputS5xD(221)(0) <= CNStageIntLLROutputS5xD(25)(3);
  VNStageIntLLRInputS5xD(285)(0) <= CNStageIntLLROutputS5xD(25)(4);
  VNStageIntLLRInputS5xD(349)(0) <= CNStageIntLLROutputS5xD(25)(5);
  VNStageIntLLRInputS5xD(28)(0) <= CNStageIntLLROutputS5xD(26)(0);
  VNStageIntLLRInputS5xD(92)(0) <= CNStageIntLLROutputS5xD(26)(1);
  VNStageIntLLRInputS5xD(156)(0) <= CNStageIntLLROutputS5xD(26)(2);
  VNStageIntLLRInputS5xD(220)(0) <= CNStageIntLLROutputS5xD(26)(3);
  VNStageIntLLRInputS5xD(284)(0) <= CNStageIntLLROutputS5xD(26)(4);
  VNStageIntLLRInputS5xD(348)(0) <= CNStageIntLLROutputS5xD(26)(5);
  VNStageIntLLRInputS5xD(27)(0) <= CNStageIntLLROutputS5xD(27)(0);
  VNStageIntLLRInputS5xD(91)(0) <= CNStageIntLLROutputS5xD(27)(1);
  VNStageIntLLRInputS5xD(155)(0) <= CNStageIntLLROutputS5xD(27)(2);
  VNStageIntLLRInputS5xD(219)(0) <= CNStageIntLLROutputS5xD(27)(3);
  VNStageIntLLRInputS5xD(283)(0) <= CNStageIntLLROutputS5xD(27)(4);
  VNStageIntLLRInputS5xD(347)(0) <= CNStageIntLLROutputS5xD(27)(5);
  VNStageIntLLRInputS5xD(26)(0) <= CNStageIntLLROutputS5xD(28)(0);
  VNStageIntLLRInputS5xD(90)(0) <= CNStageIntLLROutputS5xD(28)(1);
  VNStageIntLLRInputS5xD(154)(0) <= CNStageIntLLROutputS5xD(28)(2);
  VNStageIntLLRInputS5xD(218)(0) <= CNStageIntLLROutputS5xD(28)(3);
  VNStageIntLLRInputS5xD(282)(0) <= CNStageIntLLROutputS5xD(28)(4);
  VNStageIntLLRInputS5xD(346)(0) <= CNStageIntLLROutputS5xD(28)(5);
  VNStageIntLLRInputS5xD(25)(0) <= CNStageIntLLROutputS5xD(29)(0);
  VNStageIntLLRInputS5xD(89)(0) <= CNStageIntLLROutputS5xD(29)(1);
  VNStageIntLLRInputS5xD(153)(0) <= CNStageIntLLROutputS5xD(29)(2);
  VNStageIntLLRInputS5xD(217)(0) <= CNStageIntLLROutputS5xD(29)(3);
  VNStageIntLLRInputS5xD(281)(0) <= CNStageIntLLROutputS5xD(29)(4);
  VNStageIntLLRInputS5xD(345)(0) <= CNStageIntLLROutputS5xD(29)(5);
  VNStageIntLLRInputS5xD(24)(0) <= CNStageIntLLROutputS5xD(30)(0);
  VNStageIntLLRInputS5xD(88)(0) <= CNStageIntLLROutputS5xD(30)(1);
  VNStageIntLLRInputS5xD(152)(0) <= CNStageIntLLROutputS5xD(30)(2);
  VNStageIntLLRInputS5xD(216)(0) <= CNStageIntLLROutputS5xD(30)(3);
  VNStageIntLLRInputS5xD(280)(0) <= CNStageIntLLROutputS5xD(30)(4);
  VNStageIntLLRInputS5xD(344)(0) <= CNStageIntLLROutputS5xD(30)(5);
  VNStageIntLLRInputS5xD(23)(0) <= CNStageIntLLROutputS5xD(31)(0);
  VNStageIntLLRInputS5xD(87)(0) <= CNStageIntLLROutputS5xD(31)(1);
  VNStageIntLLRInputS5xD(151)(0) <= CNStageIntLLROutputS5xD(31)(2);
  VNStageIntLLRInputS5xD(215)(0) <= CNStageIntLLROutputS5xD(31)(3);
  VNStageIntLLRInputS5xD(279)(0) <= CNStageIntLLROutputS5xD(31)(4);
  VNStageIntLLRInputS5xD(343)(0) <= CNStageIntLLROutputS5xD(31)(5);
  VNStageIntLLRInputS5xD(22)(0) <= CNStageIntLLROutputS5xD(32)(0);
  VNStageIntLLRInputS5xD(86)(0) <= CNStageIntLLROutputS5xD(32)(1);
  VNStageIntLLRInputS5xD(150)(0) <= CNStageIntLLROutputS5xD(32)(2);
  VNStageIntLLRInputS5xD(214)(0) <= CNStageIntLLROutputS5xD(32)(3);
  VNStageIntLLRInputS5xD(278)(0) <= CNStageIntLLROutputS5xD(32)(4);
  VNStageIntLLRInputS5xD(342)(0) <= CNStageIntLLROutputS5xD(32)(5);
  VNStageIntLLRInputS5xD(21)(0) <= CNStageIntLLROutputS5xD(33)(0);
  VNStageIntLLRInputS5xD(85)(0) <= CNStageIntLLROutputS5xD(33)(1);
  VNStageIntLLRInputS5xD(149)(0) <= CNStageIntLLROutputS5xD(33)(2);
  VNStageIntLLRInputS5xD(213)(0) <= CNStageIntLLROutputS5xD(33)(3);
  VNStageIntLLRInputS5xD(277)(0) <= CNStageIntLLROutputS5xD(33)(4);
  VNStageIntLLRInputS5xD(341)(0) <= CNStageIntLLROutputS5xD(33)(5);
  VNStageIntLLRInputS5xD(20)(0) <= CNStageIntLLROutputS5xD(34)(0);
  VNStageIntLLRInputS5xD(84)(0) <= CNStageIntLLROutputS5xD(34)(1);
  VNStageIntLLRInputS5xD(148)(0) <= CNStageIntLLROutputS5xD(34)(2);
  VNStageIntLLRInputS5xD(212)(0) <= CNStageIntLLROutputS5xD(34)(3);
  VNStageIntLLRInputS5xD(276)(0) <= CNStageIntLLROutputS5xD(34)(4);
  VNStageIntLLRInputS5xD(340)(0) <= CNStageIntLLROutputS5xD(34)(5);
  VNStageIntLLRInputS5xD(19)(0) <= CNStageIntLLROutputS5xD(35)(0);
  VNStageIntLLRInputS5xD(83)(0) <= CNStageIntLLROutputS5xD(35)(1);
  VNStageIntLLRInputS5xD(147)(0) <= CNStageIntLLROutputS5xD(35)(2);
  VNStageIntLLRInputS5xD(211)(0) <= CNStageIntLLROutputS5xD(35)(3);
  VNStageIntLLRInputS5xD(275)(0) <= CNStageIntLLROutputS5xD(35)(4);
  VNStageIntLLRInputS5xD(339)(0) <= CNStageIntLLROutputS5xD(35)(5);
  VNStageIntLLRInputS5xD(18)(0) <= CNStageIntLLROutputS5xD(36)(0);
  VNStageIntLLRInputS5xD(82)(0) <= CNStageIntLLROutputS5xD(36)(1);
  VNStageIntLLRInputS5xD(146)(0) <= CNStageIntLLROutputS5xD(36)(2);
  VNStageIntLLRInputS5xD(210)(0) <= CNStageIntLLROutputS5xD(36)(3);
  VNStageIntLLRInputS5xD(274)(0) <= CNStageIntLLROutputS5xD(36)(4);
  VNStageIntLLRInputS5xD(338)(0) <= CNStageIntLLROutputS5xD(36)(5);
  VNStageIntLLRInputS5xD(17)(0) <= CNStageIntLLROutputS5xD(37)(0);
  VNStageIntLLRInputS5xD(81)(0) <= CNStageIntLLROutputS5xD(37)(1);
  VNStageIntLLRInputS5xD(145)(0) <= CNStageIntLLROutputS5xD(37)(2);
  VNStageIntLLRInputS5xD(209)(0) <= CNStageIntLLROutputS5xD(37)(3);
  VNStageIntLLRInputS5xD(273)(0) <= CNStageIntLLROutputS5xD(37)(4);
  VNStageIntLLRInputS5xD(337)(0) <= CNStageIntLLROutputS5xD(37)(5);
  VNStageIntLLRInputS5xD(16)(0) <= CNStageIntLLROutputS5xD(38)(0);
  VNStageIntLLRInputS5xD(80)(0) <= CNStageIntLLROutputS5xD(38)(1);
  VNStageIntLLRInputS5xD(144)(0) <= CNStageIntLLROutputS5xD(38)(2);
  VNStageIntLLRInputS5xD(208)(0) <= CNStageIntLLROutputS5xD(38)(3);
  VNStageIntLLRInputS5xD(272)(0) <= CNStageIntLLROutputS5xD(38)(4);
  VNStageIntLLRInputS5xD(336)(0) <= CNStageIntLLROutputS5xD(38)(5);
  VNStageIntLLRInputS5xD(15)(0) <= CNStageIntLLROutputS5xD(39)(0);
  VNStageIntLLRInputS5xD(79)(0) <= CNStageIntLLROutputS5xD(39)(1);
  VNStageIntLLRInputS5xD(143)(0) <= CNStageIntLLROutputS5xD(39)(2);
  VNStageIntLLRInputS5xD(207)(0) <= CNStageIntLLROutputS5xD(39)(3);
  VNStageIntLLRInputS5xD(271)(0) <= CNStageIntLLROutputS5xD(39)(4);
  VNStageIntLLRInputS5xD(335)(0) <= CNStageIntLLROutputS5xD(39)(5);
  VNStageIntLLRInputS5xD(14)(0) <= CNStageIntLLROutputS5xD(40)(0);
  VNStageIntLLRInputS5xD(78)(0) <= CNStageIntLLROutputS5xD(40)(1);
  VNStageIntLLRInputS5xD(142)(0) <= CNStageIntLLROutputS5xD(40)(2);
  VNStageIntLLRInputS5xD(206)(0) <= CNStageIntLLROutputS5xD(40)(3);
  VNStageIntLLRInputS5xD(270)(0) <= CNStageIntLLROutputS5xD(40)(4);
  VNStageIntLLRInputS5xD(334)(0) <= CNStageIntLLROutputS5xD(40)(5);
  VNStageIntLLRInputS5xD(12)(0) <= CNStageIntLLROutputS5xD(41)(0);
  VNStageIntLLRInputS5xD(76)(0) <= CNStageIntLLROutputS5xD(41)(1);
  VNStageIntLLRInputS5xD(140)(0) <= CNStageIntLLROutputS5xD(41)(2);
  VNStageIntLLRInputS5xD(204)(0) <= CNStageIntLLROutputS5xD(41)(3);
  VNStageIntLLRInputS5xD(268)(0) <= CNStageIntLLROutputS5xD(41)(4);
  VNStageIntLLRInputS5xD(332)(0) <= CNStageIntLLROutputS5xD(41)(5);
  VNStageIntLLRInputS5xD(11)(0) <= CNStageIntLLROutputS5xD(42)(0);
  VNStageIntLLRInputS5xD(75)(0) <= CNStageIntLLROutputS5xD(42)(1);
  VNStageIntLLRInputS5xD(139)(0) <= CNStageIntLLROutputS5xD(42)(2);
  VNStageIntLLRInputS5xD(203)(0) <= CNStageIntLLROutputS5xD(42)(3);
  VNStageIntLLRInputS5xD(267)(0) <= CNStageIntLLROutputS5xD(42)(4);
  VNStageIntLLRInputS5xD(331)(0) <= CNStageIntLLROutputS5xD(42)(5);
  VNStageIntLLRInputS5xD(10)(0) <= CNStageIntLLROutputS5xD(43)(0);
  VNStageIntLLRInputS5xD(74)(0) <= CNStageIntLLROutputS5xD(43)(1);
  VNStageIntLLRInputS5xD(138)(0) <= CNStageIntLLROutputS5xD(43)(2);
  VNStageIntLLRInputS5xD(202)(0) <= CNStageIntLLROutputS5xD(43)(3);
  VNStageIntLLRInputS5xD(266)(0) <= CNStageIntLLROutputS5xD(43)(4);
  VNStageIntLLRInputS5xD(330)(0) <= CNStageIntLLROutputS5xD(43)(5);
  VNStageIntLLRInputS5xD(9)(0) <= CNStageIntLLROutputS5xD(44)(0);
  VNStageIntLLRInputS5xD(73)(0) <= CNStageIntLLROutputS5xD(44)(1);
  VNStageIntLLRInputS5xD(137)(0) <= CNStageIntLLROutputS5xD(44)(2);
  VNStageIntLLRInputS5xD(201)(0) <= CNStageIntLLROutputS5xD(44)(3);
  VNStageIntLLRInputS5xD(265)(0) <= CNStageIntLLROutputS5xD(44)(4);
  VNStageIntLLRInputS5xD(329)(0) <= CNStageIntLLROutputS5xD(44)(5);
  VNStageIntLLRInputS5xD(8)(0) <= CNStageIntLLROutputS5xD(45)(0);
  VNStageIntLLRInputS5xD(72)(0) <= CNStageIntLLROutputS5xD(45)(1);
  VNStageIntLLRInputS5xD(136)(0) <= CNStageIntLLROutputS5xD(45)(2);
  VNStageIntLLRInputS5xD(200)(0) <= CNStageIntLLROutputS5xD(45)(3);
  VNStageIntLLRInputS5xD(264)(0) <= CNStageIntLLROutputS5xD(45)(4);
  VNStageIntLLRInputS5xD(328)(0) <= CNStageIntLLROutputS5xD(45)(5);
  VNStageIntLLRInputS5xD(7)(0) <= CNStageIntLLROutputS5xD(46)(0);
  VNStageIntLLRInputS5xD(71)(0) <= CNStageIntLLROutputS5xD(46)(1);
  VNStageIntLLRInputS5xD(135)(0) <= CNStageIntLLROutputS5xD(46)(2);
  VNStageIntLLRInputS5xD(199)(0) <= CNStageIntLLROutputS5xD(46)(3);
  VNStageIntLLRInputS5xD(263)(0) <= CNStageIntLLROutputS5xD(46)(4);
  VNStageIntLLRInputS5xD(327)(0) <= CNStageIntLLROutputS5xD(46)(5);
  VNStageIntLLRInputS5xD(6)(0) <= CNStageIntLLROutputS5xD(47)(0);
  VNStageIntLLRInputS5xD(70)(0) <= CNStageIntLLROutputS5xD(47)(1);
  VNStageIntLLRInputS5xD(134)(0) <= CNStageIntLLROutputS5xD(47)(2);
  VNStageIntLLRInputS5xD(198)(0) <= CNStageIntLLROutputS5xD(47)(3);
  VNStageIntLLRInputS5xD(262)(0) <= CNStageIntLLROutputS5xD(47)(4);
  VNStageIntLLRInputS5xD(326)(0) <= CNStageIntLLROutputS5xD(47)(5);
  VNStageIntLLRInputS5xD(5)(0) <= CNStageIntLLROutputS5xD(48)(0);
  VNStageIntLLRInputS5xD(69)(0) <= CNStageIntLLROutputS5xD(48)(1);
  VNStageIntLLRInputS5xD(133)(0) <= CNStageIntLLROutputS5xD(48)(2);
  VNStageIntLLRInputS5xD(197)(0) <= CNStageIntLLROutputS5xD(48)(3);
  VNStageIntLLRInputS5xD(261)(0) <= CNStageIntLLROutputS5xD(48)(4);
  VNStageIntLLRInputS5xD(325)(0) <= CNStageIntLLROutputS5xD(48)(5);
  VNStageIntLLRInputS5xD(4)(0) <= CNStageIntLLROutputS5xD(49)(0);
  VNStageIntLLRInputS5xD(68)(0) <= CNStageIntLLROutputS5xD(49)(1);
  VNStageIntLLRInputS5xD(132)(0) <= CNStageIntLLROutputS5xD(49)(2);
  VNStageIntLLRInputS5xD(196)(0) <= CNStageIntLLROutputS5xD(49)(3);
  VNStageIntLLRInputS5xD(260)(0) <= CNStageIntLLROutputS5xD(49)(4);
  VNStageIntLLRInputS5xD(324)(0) <= CNStageIntLLROutputS5xD(49)(5);
  VNStageIntLLRInputS5xD(2)(0) <= CNStageIntLLROutputS5xD(50)(0);
  VNStageIntLLRInputS5xD(66)(0) <= CNStageIntLLROutputS5xD(50)(1);
  VNStageIntLLRInputS5xD(130)(0) <= CNStageIntLLROutputS5xD(50)(2);
  VNStageIntLLRInputS5xD(194)(0) <= CNStageIntLLROutputS5xD(50)(3);
  VNStageIntLLRInputS5xD(258)(0) <= CNStageIntLLROutputS5xD(50)(4);
  VNStageIntLLRInputS5xD(322)(0) <= CNStageIntLLROutputS5xD(50)(5);
  VNStageIntLLRInputS5xD(1)(0) <= CNStageIntLLROutputS5xD(51)(0);
  VNStageIntLLRInputS5xD(65)(0) <= CNStageIntLLROutputS5xD(51)(1);
  VNStageIntLLRInputS5xD(129)(0) <= CNStageIntLLROutputS5xD(51)(2);
  VNStageIntLLRInputS5xD(193)(0) <= CNStageIntLLROutputS5xD(51)(3);
  VNStageIntLLRInputS5xD(257)(0) <= CNStageIntLLROutputS5xD(51)(4);
  VNStageIntLLRInputS5xD(321)(0) <= CNStageIntLLROutputS5xD(51)(5);
  VNStageIntLLRInputS5xD(63)(0) <= CNStageIntLLROutputS5xD(52)(0);
  VNStageIntLLRInputS5xD(127)(0) <= CNStageIntLLROutputS5xD(52)(1);
  VNStageIntLLRInputS5xD(191)(0) <= CNStageIntLLROutputS5xD(52)(2);
  VNStageIntLLRInputS5xD(255)(0) <= CNStageIntLLROutputS5xD(52)(3);
  VNStageIntLLRInputS5xD(319)(0) <= CNStageIntLLROutputS5xD(52)(4);
  VNStageIntLLRInputS5xD(383)(0) <= CNStageIntLLROutputS5xD(52)(5);
  VNStageIntLLRInputS5xD(0)(0) <= CNStageIntLLROutputS5xD(53)(0);
  VNStageIntLLRInputS5xD(64)(0) <= CNStageIntLLROutputS5xD(53)(1);
  VNStageIntLLRInputS5xD(128)(0) <= CNStageIntLLROutputS5xD(53)(2);
  VNStageIntLLRInputS5xD(192)(0) <= CNStageIntLLROutputS5xD(53)(3);
  VNStageIntLLRInputS5xD(256)(0) <= CNStageIntLLROutputS5xD(53)(4);
  VNStageIntLLRInputS5xD(320)(0) <= CNStageIntLLROutputS5xD(53)(5);
  VNStageIntLLRInputS5xD(42)(1) <= CNStageIntLLROutputS5xD(54)(0);
  VNStageIntLLRInputS5xD(112)(1) <= CNStageIntLLROutputS5xD(54)(1);
  VNStageIntLLRInputS5xD(182)(1) <= CNStageIntLLROutputS5xD(54)(2);
  VNStageIntLLRInputS5xD(203)(1) <= CNStageIntLLROutputS5xD(54)(3);
  VNStageIntLLRInputS5xD(259)(0) <= CNStageIntLLROutputS5xD(54)(4);
  VNStageIntLLRInputS5xD(361)(1) <= CNStageIntLLROutputS5xD(54)(5);
  VNStageIntLLRInputS5xD(41)(1) <= CNStageIntLLROutputS5xD(55)(0);
  VNStageIntLLRInputS5xD(117)(1) <= CNStageIntLLROutputS5xD(55)(1);
  VNStageIntLLRInputS5xD(138)(1) <= CNStageIntLLROutputS5xD(55)(2);
  VNStageIntLLRInputS5xD(194)(1) <= CNStageIntLLROutputS5xD(55)(3);
  VNStageIntLLRInputS5xD(296)(1) <= CNStageIntLLROutputS5xD(55)(4);
  VNStageIntLLRInputS5xD(362)(1) <= CNStageIntLLROutputS5xD(55)(5);
  VNStageIntLLRInputS5xD(40)(1) <= CNStageIntLLROutputS5xD(56)(0);
  VNStageIntLLRInputS5xD(73)(1) <= CNStageIntLLROutputS5xD(56)(1);
  VNStageIntLLRInputS5xD(129)(1) <= CNStageIntLLROutputS5xD(56)(2);
  VNStageIntLLRInputS5xD(231)(1) <= CNStageIntLLROutputS5xD(56)(3);
  VNStageIntLLRInputS5xD(297)(1) <= CNStageIntLLROutputS5xD(56)(4);
  VNStageIntLLRInputS5xD(323)(0) <= CNStageIntLLROutputS5xD(56)(5);
  VNStageIntLLRInputS5xD(39)(1) <= CNStageIntLLROutputS5xD(57)(0);
  VNStageIntLLRInputS5xD(127)(1) <= CNStageIntLLROutputS5xD(57)(1);
  VNStageIntLLRInputS5xD(166)(1) <= CNStageIntLLROutputS5xD(57)(2);
  VNStageIntLLRInputS5xD(232)(1) <= CNStageIntLLROutputS5xD(57)(3);
  VNStageIntLLRInputS5xD(258)(1) <= CNStageIntLLROutputS5xD(57)(4);
  VNStageIntLLRInputS5xD(344)(1) <= CNStageIntLLROutputS5xD(57)(5);
  VNStageIntLLRInputS5xD(38)(1) <= CNStageIntLLROutputS5xD(58)(0);
  VNStageIntLLRInputS5xD(101)(1) <= CNStageIntLLROutputS5xD(58)(1);
  VNStageIntLLRInputS5xD(167)(1) <= CNStageIntLLROutputS5xD(58)(2);
  VNStageIntLLRInputS5xD(193)(1) <= CNStageIntLLROutputS5xD(58)(3);
  VNStageIntLLRInputS5xD(279)(1) <= CNStageIntLLROutputS5xD(58)(4);
  VNStageIntLLRInputS5xD(340)(1) <= CNStageIntLLROutputS5xD(58)(5);
  VNStageIntLLRInputS5xD(37)(1) <= CNStageIntLLROutputS5xD(59)(0);
  VNStageIntLLRInputS5xD(102)(1) <= CNStageIntLLROutputS5xD(59)(1);
  VNStageIntLLRInputS5xD(191)(1) <= CNStageIntLLROutputS5xD(59)(2);
  VNStageIntLLRInputS5xD(214)(1) <= CNStageIntLLROutputS5xD(59)(3);
  VNStageIntLLRInputS5xD(275)(1) <= CNStageIntLLROutputS5xD(59)(4);
  VNStageIntLLRInputS5xD(355)(1) <= CNStageIntLLROutputS5xD(59)(5);
  VNStageIntLLRInputS5xD(36)(1) <= CNStageIntLLROutputS5xD(60)(0);
  VNStageIntLLRInputS5xD(126)(0) <= CNStageIntLLROutputS5xD(60)(1);
  VNStageIntLLRInputS5xD(149)(1) <= CNStageIntLLROutputS5xD(60)(2);
  VNStageIntLLRInputS5xD(210)(1) <= CNStageIntLLROutputS5xD(60)(3);
  VNStageIntLLRInputS5xD(290)(1) <= CNStageIntLLROutputS5xD(60)(4);
  VNStageIntLLRInputS5xD(381)(0) <= CNStageIntLLROutputS5xD(60)(5);
  VNStageIntLLRInputS5xD(35)(1) <= CNStageIntLLROutputS5xD(61)(0);
  VNStageIntLLRInputS5xD(84)(1) <= CNStageIntLLROutputS5xD(61)(1);
  VNStageIntLLRInputS5xD(145)(1) <= CNStageIntLLROutputS5xD(61)(2);
  VNStageIntLLRInputS5xD(225)(1) <= CNStageIntLLROutputS5xD(61)(3);
  VNStageIntLLRInputS5xD(316)(0) <= CNStageIntLLROutputS5xD(61)(4);
  VNStageIntLLRInputS5xD(357)(1) <= CNStageIntLLROutputS5xD(61)(5);
  VNStageIntLLRInputS5xD(34)(1) <= CNStageIntLLROutputS5xD(62)(0);
  VNStageIntLLRInputS5xD(80)(1) <= CNStageIntLLROutputS5xD(62)(1);
  VNStageIntLLRInputS5xD(160)(1) <= CNStageIntLLROutputS5xD(62)(2);
  VNStageIntLLRInputS5xD(251)(0) <= CNStageIntLLROutputS5xD(62)(3);
  VNStageIntLLRInputS5xD(292)(1) <= CNStageIntLLROutputS5xD(62)(4);
  VNStageIntLLRInputS5xD(326)(1) <= CNStageIntLLROutputS5xD(62)(5);
  VNStageIntLLRInputS5xD(33)(1) <= CNStageIntLLROutputS5xD(63)(0);
  VNStageIntLLRInputS5xD(95)(1) <= CNStageIntLLROutputS5xD(63)(1);
  VNStageIntLLRInputS5xD(186)(0) <= CNStageIntLLROutputS5xD(63)(2);
  VNStageIntLLRInputS5xD(227)(1) <= CNStageIntLLROutputS5xD(63)(3);
  VNStageIntLLRInputS5xD(261)(1) <= CNStageIntLLROutputS5xD(63)(4);
  VNStageIntLLRInputS5xD(342)(1) <= CNStageIntLLROutputS5xD(63)(5);
  VNStageIntLLRInputS5xD(32)(1) <= CNStageIntLLROutputS5xD(64)(0);
  VNStageIntLLRInputS5xD(121)(0) <= CNStageIntLLROutputS5xD(64)(1);
  VNStageIntLLRInputS5xD(162)(1) <= CNStageIntLLROutputS5xD(64)(2);
  VNStageIntLLRInputS5xD(196)(1) <= CNStageIntLLROutputS5xD(64)(3);
  VNStageIntLLRInputS5xD(277)(1) <= CNStageIntLLROutputS5xD(64)(4);
  VNStageIntLLRInputS5xD(375)(1) <= CNStageIntLLROutputS5xD(64)(5);
  VNStageIntLLRInputS5xD(31)(1) <= CNStageIntLLROutputS5xD(65)(0);
  VNStageIntLLRInputS5xD(97)(1) <= CNStageIntLLROutputS5xD(65)(1);
  VNStageIntLLRInputS5xD(131)(0) <= CNStageIntLLROutputS5xD(65)(2);
  VNStageIntLLRInputS5xD(212)(1) <= CNStageIntLLROutputS5xD(65)(3);
  VNStageIntLLRInputS5xD(310)(1) <= CNStageIntLLROutputS5xD(65)(4);
  VNStageIntLLRInputS5xD(321)(1) <= CNStageIntLLROutputS5xD(65)(5);
  VNStageIntLLRInputS5xD(30)(1) <= CNStageIntLLROutputS5xD(66)(0);
  VNStageIntLLRInputS5xD(66)(1) <= CNStageIntLLROutputS5xD(66)(1);
  VNStageIntLLRInputS5xD(147)(1) <= CNStageIntLLROutputS5xD(66)(2);
  VNStageIntLLRInputS5xD(245)(1) <= CNStageIntLLROutputS5xD(66)(3);
  VNStageIntLLRInputS5xD(319)(1) <= CNStageIntLLROutputS5xD(66)(4);
  VNStageIntLLRInputS5xD(334)(1) <= CNStageIntLLROutputS5xD(66)(5);
  VNStageIntLLRInputS5xD(29)(1) <= CNStageIntLLROutputS5xD(67)(0);
  VNStageIntLLRInputS5xD(82)(1) <= CNStageIntLLROutputS5xD(67)(1);
  VNStageIntLLRInputS5xD(180)(0) <= CNStageIntLLROutputS5xD(67)(2);
  VNStageIntLLRInputS5xD(254)(0) <= CNStageIntLLROutputS5xD(67)(3);
  VNStageIntLLRInputS5xD(269)(0) <= CNStageIntLLROutputS5xD(67)(4);
  VNStageIntLLRInputS5xD(376)(1) <= CNStageIntLLROutputS5xD(67)(5);
  VNStageIntLLRInputS5xD(28)(1) <= CNStageIntLLROutputS5xD(68)(0);
  VNStageIntLLRInputS5xD(115)(1) <= CNStageIntLLROutputS5xD(68)(1);
  VNStageIntLLRInputS5xD(189)(0) <= CNStageIntLLROutputS5xD(68)(2);
  VNStageIntLLRInputS5xD(204)(1) <= CNStageIntLLROutputS5xD(68)(3);
  VNStageIntLLRInputS5xD(311)(1) <= CNStageIntLLROutputS5xD(68)(4);
  VNStageIntLLRInputS5xD(341)(1) <= CNStageIntLLROutputS5xD(68)(5);
  VNStageIntLLRInputS5xD(27)(1) <= CNStageIntLLROutputS5xD(69)(0);
  VNStageIntLLRInputS5xD(124)(0) <= CNStageIntLLROutputS5xD(69)(1);
  VNStageIntLLRInputS5xD(139)(1) <= CNStageIntLLROutputS5xD(69)(2);
  VNStageIntLLRInputS5xD(246)(1) <= CNStageIntLLROutputS5xD(69)(3);
  VNStageIntLLRInputS5xD(276)(1) <= CNStageIntLLROutputS5xD(69)(4);
  VNStageIntLLRInputS5xD(343)(1) <= CNStageIntLLROutputS5xD(69)(5);
  VNStageIntLLRInputS5xD(26)(1) <= CNStageIntLLROutputS5xD(70)(0);
  VNStageIntLLRInputS5xD(74)(1) <= CNStageIntLLROutputS5xD(70)(1);
  VNStageIntLLRInputS5xD(181)(1) <= CNStageIntLLROutputS5xD(70)(2);
  VNStageIntLLRInputS5xD(211)(1) <= CNStageIntLLROutputS5xD(70)(3);
  VNStageIntLLRInputS5xD(278)(1) <= CNStageIntLLROutputS5xD(70)(4);
  VNStageIntLLRInputS5xD(325)(1) <= CNStageIntLLROutputS5xD(70)(5);
  VNStageIntLLRInputS5xD(25)(1) <= CNStageIntLLROutputS5xD(71)(0);
  VNStageIntLLRInputS5xD(116)(0) <= CNStageIntLLROutputS5xD(71)(1);
  VNStageIntLLRInputS5xD(146)(1) <= CNStageIntLLROutputS5xD(71)(2);
  VNStageIntLLRInputS5xD(213)(1) <= CNStageIntLLROutputS5xD(71)(3);
  VNStageIntLLRInputS5xD(260)(1) <= CNStageIntLLROutputS5xD(71)(4);
  VNStageIntLLRInputS5xD(332)(1) <= CNStageIntLLROutputS5xD(71)(5);
  VNStageIntLLRInputS5xD(24)(1) <= CNStageIntLLROutputS5xD(72)(0);
  VNStageIntLLRInputS5xD(81)(1) <= CNStageIntLLROutputS5xD(72)(1);
  VNStageIntLLRInputS5xD(148)(1) <= CNStageIntLLROutputS5xD(72)(2);
  VNStageIntLLRInputS5xD(195)(0) <= CNStageIntLLROutputS5xD(72)(3);
  VNStageIntLLRInputS5xD(267)(1) <= CNStageIntLLROutputS5xD(72)(4);
  VNStageIntLLRInputS5xD(359)(1) <= CNStageIntLLROutputS5xD(72)(5);
  VNStageIntLLRInputS5xD(23)(1) <= CNStageIntLLROutputS5xD(73)(0);
  VNStageIntLLRInputS5xD(83)(1) <= CNStageIntLLROutputS5xD(73)(1);
  VNStageIntLLRInputS5xD(130)(1) <= CNStageIntLLROutputS5xD(73)(2);
  VNStageIntLLRInputS5xD(202)(1) <= CNStageIntLLROutputS5xD(73)(3);
  VNStageIntLLRInputS5xD(294)(1) <= CNStageIntLLROutputS5xD(73)(4);
  VNStageIntLLRInputS5xD(347)(1) <= CNStageIntLLROutputS5xD(73)(5);
  VNStageIntLLRInputS5xD(22)(1) <= CNStageIntLLROutputS5xD(74)(0);
  VNStageIntLLRInputS5xD(65)(1) <= CNStageIntLLROutputS5xD(74)(1);
  VNStageIntLLRInputS5xD(137)(1) <= CNStageIntLLROutputS5xD(74)(2);
  VNStageIntLLRInputS5xD(229)(1) <= CNStageIntLLROutputS5xD(74)(3);
  VNStageIntLLRInputS5xD(282)(1) <= CNStageIntLLROutputS5xD(74)(4);
  VNStageIntLLRInputS5xD(353)(1) <= CNStageIntLLROutputS5xD(74)(5);
  VNStageIntLLRInputS5xD(21)(1) <= CNStageIntLLROutputS5xD(75)(0);
  VNStageIntLLRInputS5xD(72)(1) <= CNStageIntLLROutputS5xD(75)(1);
  VNStageIntLLRInputS5xD(164)(1) <= CNStageIntLLROutputS5xD(75)(2);
  VNStageIntLLRInputS5xD(217)(1) <= CNStageIntLLROutputS5xD(75)(3);
  VNStageIntLLRInputS5xD(288)(1) <= CNStageIntLLROutputS5xD(75)(4);
  VNStageIntLLRInputS5xD(348)(1) <= CNStageIntLLROutputS5xD(75)(5);
  VNStageIntLLRInputS5xD(20)(1) <= CNStageIntLLROutputS5xD(76)(0);
  VNStageIntLLRInputS5xD(99)(1) <= CNStageIntLLROutputS5xD(76)(1);
  VNStageIntLLRInputS5xD(152)(1) <= CNStageIntLLROutputS5xD(76)(2);
  VNStageIntLLRInputS5xD(223)(1) <= CNStageIntLLROutputS5xD(76)(3);
  VNStageIntLLRInputS5xD(283)(1) <= CNStageIntLLROutputS5xD(76)(4);
  VNStageIntLLRInputS5xD(358)(1) <= CNStageIntLLROutputS5xD(76)(5);
  VNStageIntLLRInputS5xD(19)(1) <= CNStageIntLLROutputS5xD(77)(0);
  VNStageIntLLRInputS5xD(87)(1) <= CNStageIntLLROutputS5xD(77)(1);
  VNStageIntLLRInputS5xD(158)(1) <= CNStageIntLLROutputS5xD(77)(2);
  VNStageIntLLRInputS5xD(218)(1) <= CNStageIntLLROutputS5xD(77)(3);
  VNStageIntLLRInputS5xD(293)(1) <= CNStageIntLLROutputS5xD(77)(4);
  VNStageIntLLRInputS5xD(380)(0) <= CNStageIntLLROutputS5xD(77)(5);
  VNStageIntLLRInputS5xD(18)(1) <= CNStageIntLLROutputS5xD(78)(0);
  VNStageIntLLRInputS5xD(93)(1) <= CNStageIntLLROutputS5xD(78)(1);
  VNStageIntLLRInputS5xD(153)(1) <= CNStageIntLLROutputS5xD(78)(2);
  VNStageIntLLRInputS5xD(228)(1) <= CNStageIntLLROutputS5xD(78)(3);
  VNStageIntLLRInputS5xD(315)(0) <= CNStageIntLLROutputS5xD(78)(4);
  VNStageIntLLRInputS5xD(335)(1) <= CNStageIntLLROutputS5xD(78)(5);
  VNStageIntLLRInputS5xD(17)(1) <= CNStageIntLLROutputS5xD(79)(0);
  VNStageIntLLRInputS5xD(88)(1) <= CNStageIntLLROutputS5xD(79)(1);
  VNStageIntLLRInputS5xD(163)(1) <= CNStageIntLLROutputS5xD(79)(2);
  VNStageIntLLRInputS5xD(250)(0) <= CNStageIntLLROutputS5xD(79)(3);
  VNStageIntLLRInputS5xD(270)(1) <= CNStageIntLLROutputS5xD(79)(4);
  VNStageIntLLRInputS5xD(383)(1) <= CNStageIntLLROutputS5xD(79)(5);
  VNStageIntLLRInputS5xD(15)(1) <= CNStageIntLLROutputS5xD(80)(0);
  VNStageIntLLRInputS5xD(120)(1) <= CNStageIntLLROutputS5xD(80)(1);
  VNStageIntLLRInputS5xD(140)(1) <= CNStageIntLLROutputS5xD(80)(2);
  VNStageIntLLRInputS5xD(253)(0) <= CNStageIntLLROutputS5xD(80)(3);
  VNStageIntLLRInputS5xD(305)(1) <= CNStageIntLLROutputS5xD(80)(4);
  VNStageIntLLRInputS5xD(338)(1) <= CNStageIntLLROutputS5xD(80)(5);
  VNStageIntLLRInputS5xD(14)(1) <= CNStageIntLLROutputS5xD(81)(0);
  VNStageIntLLRInputS5xD(75)(1) <= CNStageIntLLROutputS5xD(81)(1);
  VNStageIntLLRInputS5xD(188)(0) <= CNStageIntLLROutputS5xD(81)(2);
  VNStageIntLLRInputS5xD(240)(1) <= CNStageIntLLROutputS5xD(81)(3);
  VNStageIntLLRInputS5xD(273)(1) <= CNStageIntLLROutputS5xD(81)(4);
  VNStageIntLLRInputS5xD(350)(1) <= CNStageIntLLROutputS5xD(81)(5);
  VNStageIntLLRInputS5xD(13)(0) <= CNStageIntLLROutputS5xD(82)(0);
  VNStageIntLLRInputS5xD(123)(0) <= CNStageIntLLROutputS5xD(82)(1);
  VNStageIntLLRInputS5xD(175)(1) <= CNStageIntLLROutputS5xD(82)(2);
  VNStageIntLLRInputS5xD(208)(1) <= CNStageIntLLROutputS5xD(82)(3);
  VNStageIntLLRInputS5xD(285)(1) <= CNStageIntLLROutputS5xD(82)(4);
  VNStageIntLLRInputS5xD(364)(1) <= CNStageIntLLROutputS5xD(82)(5);
  VNStageIntLLRInputS5xD(12)(1) <= CNStageIntLLROutputS5xD(83)(0);
  VNStageIntLLRInputS5xD(110)(1) <= CNStageIntLLROutputS5xD(83)(1);
  VNStageIntLLRInputS5xD(143)(1) <= CNStageIntLLROutputS5xD(83)(2);
  VNStageIntLLRInputS5xD(220)(1) <= CNStageIntLLROutputS5xD(83)(3);
  VNStageIntLLRInputS5xD(299)(0) <= CNStageIntLLROutputS5xD(83)(4);
  VNStageIntLLRInputS5xD(345)(1) <= CNStageIntLLROutputS5xD(83)(5);
  VNStageIntLLRInputS5xD(11)(1) <= CNStageIntLLROutputS5xD(84)(0);
  VNStageIntLLRInputS5xD(78)(1) <= CNStageIntLLROutputS5xD(84)(1);
  VNStageIntLLRInputS5xD(155)(1) <= CNStageIntLLROutputS5xD(84)(2);
  VNStageIntLLRInputS5xD(234)(1) <= CNStageIntLLROutputS5xD(84)(3);
  VNStageIntLLRInputS5xD(280)(1) <= CNStageIntLLROutputS5xD(84)(4);
  VNStageIntLLRInputS5xD(322)(1) <= CNStageIntLLROutputS5xD(84)(5);
  VNStageIntLLRInputS5xD(10)(1) <= CNStageIntLLROutputS5xD(85)(0);
  VNStageIntLLRInputS5xD(90)(1) <= CNStageIntLLROutputS5xD(85)(1);
  VNStageIntLLRInputS5xD(169)(1) <= CNStageIntLLROutputS5xD(85)(2);
  VNStageIntLLRInputS5xD(215)(1) <= CNStageIntLLROutputS5xD(85)(3);
  VNStageIntLLRInputS5xD(257)(1) <= CNStageIntLLROutputS5xD(85)(4);
  VNStageIntLLRInputS5xD(374)(1) <= CNStageIntLLROutputS5xD(85)(5);
  VNStageIntLLRInputS5xD(9)(1) <= CNStageIntLLROutputS5xD(86)(0);
  VNStageIntLLRInputS5xD(104)(1) <= CNStageIntLLROutputS5xD(86)(1);
  VNStageIntLLRInputS5xD(150)(1) <= CNStageIntLLROutputS5xD(86)(2);
  VNStageIntLLRInputS5xD(255)(1) <= CNStageIntLLROutputS5xD(86)(3);
  VNStageIntLLRInputS5xD(309)(1) <= CNStageIntLLROutputS5xD(86)(4);
  VNStageIntLLRInputS5xD(378)(0) <= CNStageIntLLROutputS5xD(86)(5);
  VNStageIntLLRInputS5xD(7)(1) <= CNStageIntLLROutputS5xD(87)(0);
  VNStageIntLLRInputS5xD(125)(0) <= CNStageIntLLROutputS5xD(87)(1);
  VNStageIntLLRInputS5xD(179)(1) <= CNStageIntLLROutputS5xD(87)(2);
  VNStageIntLLRInputS5xD(248)(1) <= CNStageIntLLROutputS5xD(87)(3);
  VNStageIntLLRInputS5xD(306)(1) <= CNStageIntLLROutputS5xD(87)(4);
  VNStageIntLLRInputS5xD(382)(0) <= CNStageIntLLROutputS5xD(87)(5);
  VNStageIntLLRInputS5xD(6)(1) <= CNStageIntLLROutputS5xD(88)(0);
  VNStageIntLLRInputS5xD(114)(1) <= CNStageIntLLROutputS5xD(88)(1);
  VNStageIntLLRInputS5xD(183)(1) <= CNStageIntLLROutputS5xD(88)(2);
  VNStageIntLLRInputS5xD(241)(1) <= CNStageIntLLROutputS5xD(88)(3);
  VNStageIntLLRInputS5xD(317)(0) <= CNStageIntLLROutputS5xD(88)(4);
  VNStageIntLLRInputS5xD(354)(1) <= CNStageIntLLROutputS5xD(88)(5);
  VNStageIntLLRInputS5xD(5)(1) <= CNStageIntLLROutputS5xD(89)(0);
  VNStageIntLLRInputS5xD(118)(1) <= CNStageIntLLROutputS5xD(89)(1);
  VNStageIntLLRInputS5xD(176)(1) <= CNStageIntLLROutputS5xD(89)(2);
  VNStageIntLLRInputS5xD(252)(0) <= CNStageIntLLROutputS5xD(89)(3);
  VNStageIntLLRInputS5xD(289)(1) <= CNStageIntLLROutputS5xD(89)(4);
  VNStageIntLLRInputS5xD(346)(1) <= CNStageIntLLROutputS5xD(89)(5);
  VNStageIntLLRInputS5xD(4)(1) <= CNStageIntLLROutputS5xD(90)(0);
  VNStageIntLLRInputS5xD(111)(1) <= CNStageIntLLROutputS5xD(90)(1);
  VNStageIntLLRInputS5xD(187)(0) <= CNStageIntLLROutputS5xD(90)(2);
  VNStageIntLLRInputS5xD(224)(1) <= CNStageIntLLROutputS5xD(90)(3);
  VNStageIntLLRInputS5xD(281)(1) <= CNStageIntLLROutputS5xD(90)(4);
  VNStageIntLLRInputS5xD(363)(0) <= CNStageIntLLROutputS5xD(90)(5);
  VNStageIntLLRInputS5xD(3)(0) <= CNStageIntLLROutputS5xD(91)(0);
  VNStageIntLLRInputS5xD(122)(0) <= CNStageIntLLROutputS5xD(91)(1);
  VNStageIntLLRInputS5xD(159)(1) <= CNStageIntLLROutputS5xD(91)(2);
  VNStageIntLLRInputS5xD(216)(1) <= CNStageIntLLROutputS5xD(91)(3);
  VNStageIntLLRInputS5xD(298)(1) <= CNStageIntLLROutputS5xD(91)(4);
  VNStageIntLLRInputS5xD(360)(1) <= CNStageIntLLROutputS5xD(91)(5);
  VNStageIntLLRInputS5xD(2)(1) <= CNStageIntLLROutputS5xD(92)(0);
  VNStageIntLLRInputS5xD(94)(1) <= CNStageIntLLROutputS5xD(92)(1);
  VNStageIntLLRInputS5xD(151)(1) <= CNStageIntLLROutputS5xD(92)(2);
  VNStageIntLLRInputS5xD(233)(1) <= CNStageIntLLROutputS5xD(92)(3);
  VNStageIntLLRInputS5xD(295)(1) <= CNStageIntLLROutputS5xD(92)(4);
  VNStageIntLLRInputS5xD(331)(1) <= CNStageIntLLROutputS5xD(92)(5);
  VNStageIntLLRInputS5xD(63)(1) <= CNStageIntLLROutputS5xD(93)(0);
  VNStageIntLLRInputS5xD(103)(1) <= CNStageIntLLROutputS5xD(93)(1);
  VNStageIntLLRInputS5xD(165)(1) <= CNStageIntLLROutputS5xD(93)(2);
  VNStageIntLLRInputS5xD(201)(1) <= CNStageIntLLROutputS5xD(93)(3);
  VNStageIntLLRInputS5xD(286)(1) <= CNStageIntLLROutputS5xD(93)(4);
  VNStageIntLLRInputS5xD(337)(1) <= CNStageIntLLROutputS5xD(93)(5);
  VNStageIntLLRInputS5xD(62)(0) <= CNStageIntLLROutputS5xD(94)(0);
  VNStageIntLLRInputS5xD(100)(1) <= CNStageIntLLROutputS5xD(94)(1);
  VNStageIntLLRInputS5xD(136)(1) <= CNStageIntLLROutputS5xD(94)(2);
  VNStageIntLLRInputS5xD(221)(1) <= CNStageIntLLROutputS5xD(94)(3);
  VNStageIntLLRInputS5xD(272)(1) <= CNStageIntLLROutputS5xD(94)(4);
  VNStageIntLLRInputS5xD(327)(1) <= CNStageIntLLROutputS5xD(94)(5);
  VNStageIntLLRInputS5xD(61)(0) <= CNStageIntLLROutputS5xD(95)(0);
  VNStageIntLLRInputS5xD(71)(1) <= CNStageIntLLROutputS5xD(95)(1);
  VNStageIntLLRInputS5xD(156)(1) <= CNStageIntLLROutputS5xD(95)(2);
  VNStageIntLLRInputS5xD(207)(1) <= CNStageIntLLROutputS5xD(95)(3);
  VNStageIntLLRInputS5xD(262)(1) <= CNStageIntLLROutputS5xD(95)(4);
  VNStageIntLLRInputS5xD(356)(1) <= CNStageIntLLROutputS5xD(95)(5);
  VNStageIntLLRInputS5xD(60)(0) <= CNStageIntLLROutputS5xD(96)(0);
  VNStageIntLLRInputS5xD(91)(1) <= CNStageIntLLROutputS5xD(96)(1);
  VNStageIntLLRInputS5xD(142)(1) <= CNStageIntLLROutputS5xD(96)(2);
  VNStageIntLLRInputS5xD(197)(1) <= CNStageIntLLROutputS5xD(96)(3);
  VNStageIntLLRInputS5xD(291)(1) <= CNStageIntLLROutputS5xD(96)(4);
  VNStageIntLLRInputS5xD(339)(1) <= CNStageIntLLROutputS5xD(96)(5);
  VNStageIntLLRInputS5xD(58)(0) <= CNStageIntLLROutputS5xD(97)(0);
  VNStageIntLLRInputS5xD(67)(0) <= CNStageIntLLROutputS5xD(97)(1);
  VNStageIntLLRInputS5xD(161)(1) <= CNStageIntLLROutputS5xD(97)(2);
  VNStageIntLLRInputS5xD(209)(1) <= CNStageIntLLROutputS5xD(97)(3);
  VNStageIntLLRInputS5xD(304)(1) <= CNStageIntLLROutputS5xD(97)(4);
  VNStageIntLLRInputS5xD(329)(1) <= CNStageIntLLROutputS5xD(97)(5);
  VNStageIntLLRInputS5xD(57)(0) <= CNStageIntLLROutputS5xD(98)(0);
  VNStageIntLLRInputS5xD(96)(1) <= CNStageIntLLROutputS5xD(98)(1);
  VNStageIntLLRInputS5xD(144)(1) <= CNStageIntLLROutputS5xD(98)(2);
  VNStageIntLLRInputS5xD(239)(1) <= CNStageIntLLROutputS5xD(98)(3);
  VNStageIntLLRInputS5xD(264)(1) <= CNStageIntLLROutputS5xD(98)(4);
  VNStageIntLLRInputS5xD(365)(1) <= CNStageIntLLROutputS5xD(98)(5);
  VNStageIntLLRInputS5xD(56)(1) <= CNStageIntLLROutputS5xD(99)(0);
  VNStageIntLLRInputS5xD(79)(1) <= CNStageIntLLROutputS5xD(99)(1);
  VNStageIntLLRInputS5xD(174)(1) <= CNStageIntLLROutputS5xD(99)(2);
  VNStageIntLLRInputS5xD(199)(1) <= CNStageIntLLROutputS5xD(99)(3);
  VNStageIntLLRInputS5xD(300)(1) <= CNStageIntLLROutputS5xD(99)(4);
  VNStageIntLLRInputS5xD(349)(1) <= CNStageIntLLROutputS5xD(99)(5);
  VNStageIntLLRInputS5xD(55)(1) <= CNStageIntLLROutputS5xD(100)(0);
  VNStageIntLLRInputS5xD(109)(1) <= CNStageIntLLROutputS5xD(100)(1);
  VNStageIntLLRInputS5xD(134)(1) <= CNStageIntLLROutputS5xD(100)(2);
  VNStageIntLLRInputS5xD(235)(0) <= CNStageIntLLROutputS5xD(100)(3);
  VNStageIntLLRInputS5xD(284)(1) <= CNStageIntLLROutputS5xD(100)(4);
  VNStageIntLLRInputS5xD(352)(1) <= CNStageIntLLROutputS5xD(100)(5);
  VNStageIntLLRInputS5xD(54)(1) <= CNStageIntLLROutputS5xD(101)(0);
  VNStageIntLLRInputS5xD(69)(1) <= CNStageIntLLROutputS5xD(101)(1);
  VNStageIntLLRInputS5xD(170)(1) <= CNStageIntLLROutputS5xD(101)(2);
  VNStageIntLLRInputS5xD(219)(1) <= CNStageIntLLROutputS5xD(101)(3);
  VNStageIntLLRInputS5xD(287)(1) <= CNStageIntLLROutputS5xD(101)(4);
  VNStageIntLLRInputS5xD(330)(1) <= CNStageIntLLROutputS5xD(101)(5);
  VNStageIntLLRInputS5xD(52)(0) <= CNStageIntLLROutputS5xD(102)(0);
  VNStageIntLLRInputS5xD(89)(1) <= CNStageIntLLROutputS5xD(102)(1);
  VNStageIntLLRInputS5xD(157)(1) <= CNStageIntLLROutputS5xD(102)(2);
  VNStageIntLLRInputS5xD(200)(1) <= CNStageIntLLROutputS5xD(102)(3);
  VNStageIntLLRInputS5xD(303)(1) <= CNStageIntLLROutputS5xD(102)(4);
  VNStageIntLLRInputS5xD(366)(1) <= CNStageIntLLROutputS5xD(102)(5);
  VNStageIntLLRInputS5xD(51)(1) <= CNStageIntLLROutputS5xD(103)(0);
  VNStageIntLLRInputS5xD(92)(1) <= CNStageIntLLROutputS5xD(103)(1);
  VNStageIntLLRInputS5xD(135)(1) <= CNStageIntLLROutputS5xD(103)(2);
  VNStageIntLLRInputS5xD(238)(1) <= CNStageIntLLROutputS5xD(103)(3);
  VNStageIntLLRInputS5xD(301)(1) <= CNStageIntLLROutputS5xD(103)(4);
  VNStageIntLLRInputS5xD(328)(1) <= CNStageIntLLROutputS5xD(103)(5);
  VNStageIntLLRInputS5xD(50)(1) <= CNStageIntLLROutputS5xD(104)(0);
  VNStageIntLLRInputS5xD(70)(1) <= CNStageIntLLROutputS5xD(104)(1);
  VNStageIntLLRInputS5xD(173)(1) <= CNStageIntLLROutputS5xD(104)(2);
  VNStageIntLLRInputS5xD(236)(1) <= CNStageIntLLROutputS5xD(104)(3);
  VNStageIntLLRInputS5xD(263)(1) <= CNStageIntLLROutputS5xD(104)(4);
  VNStageIntLLRInputS5xD(336)(1) <= CNStageIntLLROutputS5xD(104)(5);
  VNStageIntLLRInputS5xD(49)(1) <= CNStageIntLLROutputS5xD(105)(0);
  VNStageIntLLRInputS5xD(108)(1) <= CNStageIntLLROutputS5xD(105)(1);
  VNStageIntLLRInputS5xD(171)(0) <= CNStageIntLLROutputS5xD(105)(2);
  VNStageIntLLRInputS5xD(198)(1) <= CNStageIntLLROutputS5xD(105)(3);
  VNStageIntLLRInputS5xD(271)(1) <= CNStageIntLLROutputS5xD(105)(4);
  VNStageIntLLRInputS5xD(379)(0) <= CNStageIntLLROutputS5xD(105)(5);
  VNStageIntLLRInputS5xD(46)(1) <= CNStageIntLLROutputS5xD(106)(0);
  VNStageIntLLRInputS5xD(76)(1) <= CNStageIntLLROutputS5xD(106)(1);
  VNStageIntLLRInputS5xD(184)(1) <= CNStageIntLLROutputS5xD(106)(2);
  VNStageIntLLRInputS5xD(243)(1) <= CNStageIntLLROutputS5xD(106)(3);
  VNStageIntLLRInputS5xD(256)(1) <= CNStageIntLLROutputS5xD(106)(4);
  VNStageIntLLRInputS5xD(372)(0) <= CNStageIntLLROutputS5xD(106)(5);
  VNStageIntLLRInputS5xD(45)(1) <= CNStageIntLLROutputS5xD(107)(0);
  VNStageIntLLRInputS5xD(119)(1) <= CNStageIntLLROutputS5xD(107)(1);
  VNStageIntLLRInputS5xD(178)(1) <= CNStageIntLLROutputS5xD(107)(2);
  VNStageIntLLRInputS5xD(192)(1) <= CNStageIntLLROutputS5xD(107)(3);
  VNStageIntLLRInputS5xD(307)(1) <= CNStageIntLLROutputS5xD(107)(4);
  VNStageIntLLRInputS5xD(377)(0) <= CNStageIntLLROutputS5xD(107)(5);
  VNStageIntLLRInputS5xD(44)(1) <= CNStageIntLLROutputS5xD(108)(0);
  VNStageIntLLRInputS5xD(113)(1) <= CNStageIntLLROutputS5xD(108)(1);
  VNStageIntLLRInputS5xD(128)(1) <= CNStageIntLLROutputS5xD(108)(2);
  VNStageIntLLRInputS5xD(242)(1) <= CNStageIntLLROutputS5xD(108)(3);
  VNStageIntLLRInputS5xD(312)(1) <= CNStageIntLLROutputS5xD(108)(4);
  VNStageIntLLRInputS5xD(333)(0) <= CNStageIntLLROutputS5xD(108)(5);
  VNStageIntLLRInputS5xD(43)(0) <= CNStageIntLLROutputS5xD(109)(0);
  VNStageIntLLRInputS5xD(64)(1) <= CNStageIntLLROutputS5xD(109)(1);
  VNStageIntLLRInputS5xD(177)(1) <= CNStageIntLLROutputS5xD(109)(2);
  VNStageIntLLRInputS5xD(247)(1) <= CNStageIntLLROutputS5xD(109)(3);
  VNStageIntLLRInputS5xD(268)(1) <= CNStageIntLLROutputS5xD(109)(4);
  VNStageIntLLRInputS5xD(324)(1) <= CNStageIntLLROutputS5xD(109)(5);
  VNStageIntLLRInputS5xD(0)(1) <= CNStageIntLLROutputS5xD(110)(0);
  VNStageIntLLRInputS5xD(107)(0) <= CNStageIntLLROutputS5xD(110)(1);
  VNStageIntLLRInputS5xD(172)(1) <= CNStageIntLLROutputS5xD(110)(2);
  VNStageIntLLRInputS5xD(237)(1) <= CNStageIntLLROutputS5xD(110)(3);
  VNStageIntLLRInputS5xD(302)(1) <= CNStageIntLLROutputS5xD(110)(4);
  VNStageIntLLRInputS5xD(367)(1) <= CNStageIntLLROutputS5xD(110)(5);
  VNStageIntLLRInputS5xD(32)(2) <= CNStageIntLLROutputS5xD(111)(0);
  VNStageIntLLRInputS5xD(117)(2) <= CNStageIntLLROutputS5xD(111)(1);
  VNStageIntLLRInputS5xD(136)(2) <= CNStageIntLLROutputS5xD(111)(2);
  VNStageIntLLRInputS5xD(198)(2) <= CNStageIntLLROutputS5xD(111)(3);
  VNStageIntLLRInputS5xD(297)(2) <= CNStageIntLLROutputS5xD(111)(4);
  VNStageIntLLRInputS5xD(382)(1) <= CNStageIntLLROutputS5xD(111)(5);
  VNStageIntLLRInputS5xD(30)(2) <= CNStageIntLLROutputS5xD(112)(0);
  VNStageIntLLRInputS5xD(68)(1) <= CNStageIntLLROutputS5xD(112)(1);
  VNStageIntLLRInputS5xD(167)(2) <= CNStageIntLLROutputS5xD(112)(2);
  VNStageIntLLRInputS5xD(252)(1) <= CNStageIntLLROutputS5xD(112)(3);
  VNStageIntLLRInputS5xD(303)(2) <= CNStageIntLLROutputS5xD(112)(4);
  VNStageIntLLRInputS5xD(358)(2) <= CNStageIntLLROutputS5xD(112)(5);
  VNStageIntLLRInputS5xD(29)(2) <= CNStageIntLLROutputS5xD(113)(0);
  VNStageIntLLRInputS5xD(102)(2) <= CNStageIntLLROutputS5xD(113)(1);
  VNStageIntLLRInputS5xD(187)(1) <= CNStageIntLLROutputS5xD(113)(2);
  VNStageIntLLRInputS5xD(238)(2) <= CNStageIntLLROutputS5xD(113)(3);
  VNStageIntLLRInputS5xD(293)(2) <= CNStageIntLLROutputS5xD(113)(4);
  VNStageIntLLRInputS5xD(324)(2) <= CNStageIntLLROutputS5xD(113)(5);
  VNStageIntLLRInputS5xD(28)(2) <= CNStageIntLLROutputS5xD(114)(0);
  VNStageIntLLRInputS5xD(122)(1) <= CNStageIntLLROutputS5xD(114)(1);
  VNStageIntLLRInputS5xD(173)(2) <= CNStageIntLLROutputS5xD(114)(2);
  VNStageIntLLRInputS5xD(228)(2) <= CNStageIntLLROutputS5xD(114)(3);
  VNStageIntLLRInputS5xD(259)(1) <= CNStageIntLLROutputS5xD(114)(4);
  VNStageIntLLRInputS5xD(370)(1) <= CNStageIntLLROutputS5xD(114)(5);
  VNStageIntLLRInputS5xD(27)(2) <= CNStageIntLLROutputS5xD(115)(0);
  VNStageIntLLRInputS5xD(108)(2) <= CNStageIntLLROutputS5xD(115)(1);
  VNStageIntLLRInputS5xD(163)(2) <= CNStageIntLLROutputS5xD(115)(2);
  VNStageIntLLRInputS5xD(194)(2) <= CNStageIntLLROutputS5xD(115)(3);
  VNStageIntLLRInputS5xD(305)(2) <= CNStageIntLLROutputS5xD(115)(4);
  VNStageIntLLRInputS5xD(337)(2) <= CNStageIntLLROutputS5xD(115)(5);
  VNStageIntLLRInputS5xD(26)(2) <= CNStageIntLLROutputS5xD(116)(0);
  VNStageIntLLRInputS5xD(98)(1) <= CNStageIntLLROutputS5xD(116)(1);
  VNStageIntLLRInputS5xD(129)(2) <= CNStageIntLLROutputS5xD(116)(2);
  VNStageIntLLRInputS5xD(240)(2) <= CNStageIntLLROutputS5xD(116)(3);
  VNStageIntLLRInputS5xD(272)(2) <= CNStageIntLLROutputS5xD(116)(4);
  VNStageIntLLRInputS5xD(360)(2) <= CNStageIntLLROutputS5xD(116)(5);
  VNStageIntLLRInputS5xD(25)(2) <= CNStageIntLLROutputS5xD(117)(0);
  VNStageIntLLRInputS5xD(127)(2) <= CNStageIntLLROutputS5xD(117)(1);
  VNStageIntLLRInputS5xD(175)(2) <= CNStageIntLLROutputS5xD(117)(2);
  VNStageIntLLRInputS5xD(207)(2) <= CNStageIntLLROutputS5xD(117)(3);
  VNStageIntLLRInputS5xD(295)(2) <= CNStageIntLLROutputS5xD(117)(4);
  VNStageIntLLRInputS5xD(333)(1) <= CNStageIntLLROutputS5xD(117)(5);
  VNStageIntLLRInputS5xD(24)(2) <= CNStageIntLLROutputS5xD(118)(0);
  VNStageIntLLRInputS5xD(110)(2) <= CNStageIntLLROutputS5xD(118)(1);
  VNStageIntLLRInputS5xD(142)(2) <= CNStageIntLLROutputS5xD(118)(2);
  VNStageIntLLRInputS5xD(230)(1) <= CNStageIntLLROutputS5xD(118)(3);
  VNStageIntLLRInputS5xD(268)(2) <= CNStageIntLLROutputS5xD(118)(4);
  VNStageIntLLRInputS5xD(380)(1) <= CNStageIntLLROutputS5xD(118)(5);
  VNStageIntLLRInputS5xD(23)(2) <= CNStageIntLLROutputS5xD(119)(0);
  VNStageIntLLRInputS5xD(77)(0) <= CNStageIntLLROutputS5xD(119)(1);
  VNStageIntLLRInputS5xD(165)(2) <= CNStageIntLLROutputS5xD(119)(2);
  VNStageIntLLRInputS5xD(203)(2) <= CNStageIntLLROutputS5xD(119)(3);
  VNStageIntLLRInputS5xD(315)(1) <= CNStageIntLLROutputS5xD(119)(4);
  VNStageIntLLRInputS5xD(383)(2) <= CNStageIntLLROutputS5xD(119)(5);
  VNStageIntLLRInputS5xD(22)(2) <= CNStageIntLLROutputS5xD(120)(0);
  VNStageIntLLRInputS5xD(100)(2) <= CNStageIntLLROutputS5xD(120)(1);
  VNStageIntLLRInputS5xD(138)(2) <= CNStageIntLLROutputS5xD(120)(2);
  VNStageIntLLRInputS5xD(250)(1) <= CNStageIntLLROutputS5xD(120)(3);
  VNStageIntLLRInputS5xD(318)(0) <= CNStageIntLLROutputS5xD(120)(4);
  VNStageIntLLRInputS5xD(361)(2) <= CNStageIntLLROutputS5xD(120)(5);
  VNStageIntLLRInputS5xD(21)(2) <= CNStageIntLLROutputS5xD(121)(0);
  VNStageIntLLRInputS5xD(73)(2) <= CNStageIntLLROutputS5xD(121)(1);
  VNStageIntLLRInputS5xD(185)(0) <= CNStageIntLLROutputS5xD(121)(2);
  VNStageIntLLRInputS5xD(253)(1) <= CNStageIntLLROutputS5xD(121)(3);
  VNStageIntLLRInputS5xD(296)(2) <= CNStageIntLLROutputS5xD(121)(4);
  VNStageIntLLRInputS5xD(336)(2) <= CNStageIntLLROutputS5xD(121)(5);
  VNStageIntLLRInputS5xD(19)(2) <= CNStageIntLLROutputS5xD(122)(0);
  VNStageIntLLRInputS5xD(123)(1) <= CNStageIntLLROutputS5xD(122)(1);
  VNStageIntLLRInputS5xD(166)(2) <= CNStageIntLLROutputS5xD(122)(2);
  VNStageIntLLRInputS5xD(206)(1) <= CNStageIntLLROutputS5xD(122)(3);
  VNStageIntLLRInputS5xD(269)(1) <= CNStageIntLLROutputS5xD(122)(4);
  VNStageIntLLRInputS5xD(359)(2) <= CNStageIntLLROutputS5xD(122)(5);
  VNStageIntLLRInputS5xD(18)(2) <= CNStageIntLLROutputS5xD(123)(0);
  VNStageIntLLRInputS5xD(101)(2) <= CNStageIntLLROutputS5xD(123)(1);
  VNStageIntLLRInputS5xD(141)(0) <= CNStageIntLLROutputS5xD(123)(2);
  VNStageIntLLRInputS5xD(204)(2) <= CNStageIntLLROutputS5xD(123)(3);
  VNStageIntLLRInputS5xD(294)(2) <= CNStageIntLLROutputS5xD(123)(4);
  VNStageIntLLRInputS5xD(367)(2) <= CNStageIntLLROutputS5xD(123)(5);
  VNStageIntLLRInputS5xD(17)(2) <= CNStageIntLLROutputS5xD(124)(0);
  VNStageIntLLRInputS5xD(76)(2) <= CNStageIntLLROutputS5xD(124)(1);
  VNStageIntLLRInputS5xD(139)(2) <= CNStageIntLLROutputS5xD(124)(2);
  VNStageIntLLRInputS5xD(229)(2) <= CNStageIntLLROutputS5xD(124)(3);
  VNStageIntLLRInputS5xD(302)(2) <= CNStageIntLLROutputS5xD(124)(4);
  VNStageIntLLRInputS5xD(347)(2) <= CNStageIntLLROutputS5xD(124)(5);
  VNStageIntLLRInputS5xD(16)(1) <= CNStageIntLLROutputS5xD(125)(0);
  VNStageIntLLRInputS5xD(74)(2) <= CNStageIntLLROutputS5xD(125)(1);
  VNStageIntLLRInputS5xD(164)(2) <= CNStageIntLLROutputS5xD(125)(2);
  VNStageIntLLRInputS5xD(237)(2) <= CNStageIntLLROutputS5xD(125)(3);
  VNStageIntLLRInputS5xD(282)(2) <= CNStageIntLLROutputS5xD(125)(4);
  VNStageIntLLRInputS5xD(341)(2) <= CNStageIntLLROutputS5xD(125)(5);
  VNStageIntLLRInputS5xD(15)(2) <= CNStageIntLLROutputS5xD(126)(0);
  VNStageIntLLRInputS5xD(99)(2) <= CNStageIntLLROutputS5xD(126)(1);
  VNStageIntLLRInputS5xD(172)(2) <= CNStageIntLLROutputS5xD(126)(2);
  VNStageIntLLRInputS5xD(217)(2) <= CNStageIntLLROutputS5xD(126)(3);
  VNStageIntLLRInputS5xD(276)(2) <= CNStageIntLLROutputS5xD(126)(4);
  VNStageIntLLRInputS5xD(320)(1) <= CNStageIntLLROutputS5xD(126)(5);
  VNStageIntLLRInputS5xD(14)(2) <= CNStageIntLLROutputS5xD(127)(0);
  VNStageIntLLRInputS5xD(107)(1) <= CNStageIntLLROutputS5xD(127)(1);
  VNStageIntLLRInputS5xD(152)(2) <= CNStageIntLLROutputS5xD(127)(2);
  VNStageIntLLRInputS5xD(211)(2) <= CNStageIntLLROutputS5xD(127)(3);
  VNStageIntLLRInputS5xD(256)(2) <= CNStageIntLLROutputS5xD(127)(4);
  VNStageIntLLRInputS5xD(340)(2) <= CNStageIntLLROutputS5xD(127)(5);
  VNStageIntLLRInputS5xD(13)(1) <= CNStageIntLLROutputS5xD(128)(0);
  VNStageIntLLRInputS5xD(87)(2) <= CNStageIntLLROutputS5xD(128)(1);
  VNStageIntLLRInputS5xD(146)(2) <= CNStageIntLLROutputS5xD(128)(2);
  VNStageIntLLRInputS5xD(192)(2) <= CNStageIntLLROutputS5xD(128)(3);
  VNStageIntLLRInputS5xD(275)(2) <= CNStageIntLLROutputS5xD(128)(4);
  VNStageIntLLRInputS5xD(345)(2) <= CNStageIntLLROutputS5xD(128)(5);
  VNStageIntLLRInputS5xD(12)(2) <= CNStageIntLLROutputS5xD(129)(0);
  VNStageIntLLRInputS5xD(81)(2) <= CNStageIntLLROutputS5xD(129)(1);
  VNStageIntLLRInputS5xD(128)(2) <= CNStageIntLLROutputS5xD(129)(2);
  VNStageIntLLRInputS5xD(210)(2) <= CNStageIntLLROutputS5xD(129)(3);
  VNStageIntLLRInputS5xD(280)(2) <= CNStageIntLLROutputS5xD(129)(4);
  VNStageIntLLRInputS5xD(364)(2) <= CNStageIntLLROutputS5xD(129)(5);
  VNStageIntLLRInputS5xD(11)(2) <= CNStageIntLLROutputS5xD(130)(0);
  VNStageIntLLRInputS5xD(64)(2) <= CNStageIntLLROutputS5xD(130)(1);
  VNStageIntLLRInputS5xD(145)(2) <= CNStageIntLLROutputS5xD(130)(2);
  VNStageIntLLRInputS5xD(215)(2) <= CNStageIntLLROutputS5xD(130)(3);
  VNStageIntLLRInputS5xD(299)(1) <= CNStageIntLLROutputS5xD(130)(4);
  VNStageIntLLRInputS5xD(355)(2) <= CNStageIntLLROutputS5xD(130)(5);
  VNStageIntLLRInputS5xD(10)(2) <= CNStageIntLLROutputS5xD(131)(0);
  VNStageIntLLRInputS5xD(80)(2) <= CNStageIntLLROutputS5xD(131)(1);
  VNStageIntLLRInputS5xD(150)(2) <= CNStageIntLLROutputS5xD(131)(2);
  VNStageIntLLRInputS5xD(234)(2) <= CNStageIntLLROutputS5xD(131)(3);
  VNStageIntLLRInputS5xD(290)(2) <= CNStageIntLLROutputS5xD(131)(4);
  VNStageIntLLRInputS5xD(329)(2) <= CNStageIntLLROutputS5xD(131)(5);
  VNStageIntLLRInputS5xD(9)(2) <= CNStageIntLLROutputS5xD(132)(0);
  VNStageIntLLRInputS5xD(85)(1) <= CNStageIntLLROutputS5xD(132)(1);
  VNStageIntLLRInputS5xD(169)(2) <= CNStageIntLLROutputS5xD(132)(2);
  VNStageIntLLRInputS5xD(225)(2) <= CNStageIntLLROutputS5xD(132)(3);
  VNStageIntLLRInputS5xD(264)(2) <= CNStageIntLLROutputS5xD(132)(4);
  VNStageIntLLRInputS5xD(330)(2) <= CNStageIntLLROutputS5xD(132)(5);
  VNStageIntLLRInputS5xD(8)(1) <= CNStageIntLLROutputS5xD(133)(0);
  VNStageIntLLRInputS5xD(104)(2) <= CNStageIntLLROutputS5xD(133)(1);
  VNStageIntLLRInputS5xD(160)(2) <= CNStageIntLLROutputS5xD(133)(2);
  VNStageIntLLRInputS5xD(199)(2) <= CNStageIntLLROutputS5xD(133)(3);
  VNStageIntLLRInputS5xD(265)(1) <= CNStageIntLLROutputS5xD(133)(4);
  VNStageIntLLRInputS5xD(354)(2) <= CNStageIntLLROutputS5xD(133)(5);
  VNStageIntLLRInputS5xD(7)(2) <= CNStageIntLLROutputS5xD(134)(0);
  VNStageIntLLRInputS5xD(95)(2) <= CNStageIntLLROutputS5xD(134)(1);
  VNStageIntLLRInputS5xD(134)(2) <= CNStageIntLLROutputS5xD(134)(2);
  VNStageIntLLRInputS5xD(200)(2) <= CNStageIntLLROutputS5xD(134)(3);
  VNStageIntLLRInputS5xD(289)(2) <= CNStageIntLLROutputS5xD(134)(4);
  VNStageIntLLRInputS5xD(375)(2) <= CNStageIntLLROutputS5xD(134)(5);
  VNStageIntLLRInputS5xD(6)(2) <= CNStageIntLLROutputS5xD(135)(0);
  VNStageIntLLRInputS5xD(69)(2) <= CNStageIntLLROutputS5xD(135)(1);
  VNStageIntLLRInputS5xD(135)(2) <= CNStageIntLLROutputS5xD(135)(2);
  VNStageIntLLRInputS5xD(224)(2) <= CNStageIntLLROutputS5xD(135)(3);
  VNStageIntLLRInputS5xD(310)(2) <= CNStageIntLLROutputS5xD(135)(4);
  VNStageIntLLRInputS5xD(371)(1) <= CNStageIntLLROutputS5xD(135)(5);
  VNStageIntLLRInputS5xD(5)(2) <= CNStageIntLLROutputS5xD(136)(0);
  VNStageIntLLRInputS5xD(70)(2) <= CNStageIntLLROutputS5xD(136)(1);
  VNStageIntLLRInputS5xD(159)(2) <= CNStageIntLLROutputS5xD(136)(2);
  VNStageIntLLRInputS5xD(245)(2) <= CNStageIntLLROutputS5xD(136)(3);
  VNStageIntLLRInputS5xD(306)(2) <= CNStageIntLLROutputS5xD(136)(4);
  VNStageIntLLRInputS5xD(323)(1) <= CNStageIntLLROutputS5xD(136)(5);
  VNStageIntLLRInputS5xD(3)(1) <= CNStageIntLLROutputS5xD(137)(0);
  VNStageIntLLRInputS5xD(115)(2) <= CNStageIntLLROutputS5xD(137)(1);
  VNStageIntLLRInputS5xD(176)(2) <= CNStageIntLLROutputS5xD(137)(2);
  VNStageIntLLRInputS5xD(193)(2) <= CNStageIntLLROutputS5xD(137)(3);
  VNStageIntLLRInputS5xD(284)(2) <= CNStageIntLLROutputS5xD(137)(4);
  VNStageIntLLRInputS5xD(325)(2) <= CNStageIntLLROutputS5xD(137)(5);
  VNStageIntLLRInputS5xD(2)(2) <= CNStageIntLLROutputS5xD(138)(0);
  VNStageIntLLRInputS5xD(111)(2) <= CNStageIntLLROutputS5xD(138)(1);
  VNStageIntLLRInputS5xD(191)(2) <= CNStageIntLLROutputS5xD(138)(2);
  VNStageIntLLRInputS5xD(219)(2) <= CNStageIntLLROutputS5xD(138)(3);
  VNStageIntLLRInputS5xD(260)(2) <= CNStageIntLLROutputS5xD(138)(4);
  VNStageIntLLRInputS5xD(357)(2) <= CNStageIntLLROutputS5xD(138)(5);
  VNStageIntLLRInputS5xD(1)(1) <= CNStageIntLLROutputS5xD(139)(0);
  VNStageIntLLRInputS5xD(126)(1) <= CNStageIntLLROutputS5xD(139)(1);
  VNStageIntLLRInputS5xD(154)(1) <= CNStageIntLLROutputS5xD(139)(2);
  VNStageIntLLRInputS5xD(195)(1) <= CNStageIntLLROutputS5xD(139)(3);
  VNStageIntLLRInputS5xD(292)(2) <= CNStageIntLLROutputS5xD(139)(4);
  VNStageIntLLRInputS5xD(373)(1) <= CNStageIntLLROutputS5xD(139)(5);
  VNStageIntLLRInputS5xD(63)(2) <= CNStageIntLLROutputS5xD(140)(0);
  VNStageIntLLRInputS5xD(89)(2) <= CNStageIntLLROutputS5xD(140)(1);
  VNStageIntLLRInputS5xD(130)(2) <= CNStageIntLLROutputS5xD(140)(2);
  VNStageIntLLRInputS5xD(227)(2) <= CNStageIntLLROutputS5xD(140)(3);
  VNStageIntLLRInputS5xD(308)(0) <= CNStageIntLLROutputS5xD(140)(4);
  VNStageIntLLRInputS5xD(343)(2) <= CNStageIntLLROutputS5xD(140)(5);
  VNStageIntLLRInputS5xD(62)(1) <= CNStageIntLLROutputS5xD(141)(0);
  VNStageIntLLRInputS5xD(65)(2) <= CNStageIntLLROutputS5xD(141)(1);
  VNStageIntLLRInputS5xD(162)(2) <= CNStageIntLLROutputS5xD(141)(2);
  VNStageIntLLRInputS5xD(243)(2) <= CNStageIntLLROutputS5xD(141)(3);
  VNStageIntLLRInputS5xD(278)(2) <= CNStageIntLLROutputS5xD(141)(4);
  VNStageIntLLRInputS5xD(352)(2) <= CNStageIntLLROutputS5xD(141)(5);
  VNStageIntLLRInputS5xD(61)(1) <= CNStageIntLLROutputS5xD(142)(0);
  VNStageIntLLRInputS5xD(97)(2) <= CNStageIntLLROutputS5xD(142)(1);
  VNStageIntLLRInputS5xD(178)(2) <= CNStageIntLLROutputS5xD(142)(2);
  VNStageIntLLRInputS5xD(213)(2) <= CNStageIntLLROutputS5xD(142)(3);
  VNStageIntLLRInputS5xD(287)(2) <= CNStageIntLLROutputS5xD(142)(4);
  VNStageIntLLRInputS5xD(365)(2) <= CNStageIntLLROutputS5xD(142)(5);
  VNStageIntLLRInputS5xD(60)(1) <= CNStageIntLLROutputS5xD(143)(0);
  VNStageIntLLRInputS5xD(113)(2) <= CNStageIntLLROutputS5xD(143)(1);
  VNStageIntLLRInputS5xD(148)(2) <= CNStageIntLLROutputS5xD(143)(2);
  VNStageIntLLRInputS5xD(222)(1) <= CNStageIntLLROutputS5xD(143)(3);
  VNStageIntLLRInputS5xD(300)(2) <= CNStageIntLLROutputS5xD(143)(4);
  VNStageIntLLRInputS5xD(344)(2) <= CNStageIntLLROutputS5xD(143)(5);
  VNStageIntLLRInputS5xD(59)(0) <= CNStageIntLLROutputS5xD(144)(0);
  VNStageIntLLRInputS5xD(83)(2) <= CNStageIntLLROutputS5xD(144)(1);
  VNStageIntLLRInputS5xD(157)(2) <= CNStageIntLLROutputS5xD(144)(2);
  VNStageIntLLRInputS5xD(235)(1) <= CNStageIntLLROutputS5xD(144)(3);
  VNStageIntLLRInputS5xD(279)(2) <= CNStageIntLLROutputS5xD(144)(4);
  VNStageIntLLRInputS5xD(372)(1) <= CNStageIntLLROutputS5xD(144)(5);
  VNStageIntLLRInputS5xD(58)(1) <= CNStageIntLLROutputS5xD(145)(0);
  VNStageIntLLRInputS5xD(92)(2) <= CNStageIntLLROutputS5xD(145)(1);
  VNStageIntLLRInputS5xD(170)(2) <= CNStageIntLLROutputS5xD(145)(2);
  VNStageIntLLRInputS5xD(214)(2) <= CNStageIntLLROutputS5xD(145)(3);
  VNStageIntLLRInputS5xD(307)(2) <= CNStageIntLLROutputS5xD(145)(4);
  VNStageIntLLRInputS5xD(374)(2) <= CNStageIntLLROutputS5xD(145)(5);
  VNStageIntLLRInputS5xD(57)(1) <= CNStageIntLLROutputS5xD(146)(0);
  VNStageIntLLRInputS5xD(105)(1) <= CNStageIntLLROutputS5xD(146)(1);
  VNStageIntLLRInputS5xD(149)(2) <= CNStageIntLLROutputS5xD(146)(2);
  VNStageIntLLRInputS5xD(242)(2) <= CNStageIntLLROutputS5xD(146)(3);
  VNStageIntLLRInputS5xD(309)(2) <= CNStageIntLLROutputS5xD(146)(4);
  VNStageIntLLRInputS5xD(356)(2) <= CNStageIntLLROutputS5xD(146)(5);
  VNStageIntLLRInputS5xD(56)(2) <= CNStageIntLLROutputS5xD(147)(0);
  VNStageIntLLRInputS5xD(84)(2) <= CNStageIntLLROutputS5xD(147)(1);
  VNStageIntLLRInputS5xD(177)(2) <= CNStageIntLLROutputS5xD(147)(2);
  VNStageIntLLRInputS5xD(244)(0) <= CNStageIntLLROutputS5xD(147)(3);
  VNStageIntLLRInputS5xD(291)(2) <= CNStageIntLLROutputS5xD(147)(4);
  VNStageIntLLRInputS5xD(363)(1) <= CNStageIntLLROutputS5xD(147)(5);
  VNStageIntLLRInputS5xD(55)(2) <= CNStageIntLLROutputS5xD(148)(0);
  VNStageIntLLRInputS5xD(112)(2) <= CNStageIntLLROutputS5xD(148)(1);
  VNStageIntLLRInputS5xD(179)(2) <= CNStageIntLLROutputS5xD(148)(2);
  VNStageIntLLRInputS5xD(226)(1) <= CNStageIntLLROutputS5xD(148)(3);
  VNStageIntLLRInputS5xD(298)(2) <= CNStageIntLLROutputS5xD(148)(4);
  VNStageIntLLRInputS5xD(327)(2) <= CNStageIntLLROutputS5xD(148)(5);
  VNStageIntLLRInputS5xD(54)(2) <= CNStageIntLLROutputS5xD(149)(0);
  VNStageIntLLRInputS5xD(114)(2) <= CNStageIntLLROutputS5xD(149)(1);
  VNStageIntLLRInputS5xD(161)(2) <= CNStageIntLLROutputS5xD(149)(2);
  VNStageIntLLRInputS5xD(233)(2) <= CNStageIntLLROutputS5xD(149)(3);
  VNStageIntLLRInputS5xD(262)(2) <= CNStageIntLLROutputS5xD(149)(4);
  VNStageIntLLRInputS5xD(378)(1) <= CNStageIntLLROutputS5xD(149)(5);
  VNStageIntLLRInputS5xD(53)(1) <= CNStageIntLLROutputS5xD(150)(0);
  VNStageIntLLRInputS5xD(96)(2) <= CNStageIntLLROutputS5xD(150)(1);
  VNStageIntLLRInputS5xD(168)(1) <= CNStageIntLLROutputS5xD(150)(2);
  VNStageIntLLRInputS5xD(197)(2) <= CNStageIntLLROutputS5xD(150)(3);
  VNStageIntLLRInputS5xD(313)(0) <= CNStageIntLLROutputS5xD(150)(4);
  VNStageIntLLRInputS5xD(321)(2) <= CNStageIntLLROutputS5xD(150)(5);
  VNStageIntLLRInputS5xD(52)(1) <= CNStageIntLLROutputS5xD(151)(0);
  VNStageIntLLRInputS5xD(103)(2) <= CNStageIntLLROutputS5xD(151)(1);
  VNStageIntLLRInputS5xD(132)(1) <= CNStageIntLLROutputS5xD(151)(2);
  VNStageIntLLRInputS5xD(248)(2) <= CNStageIntLLROutputS5xD(151)(3);
  VNStageIntLLRInputS5xD(319)(2) <= CNStageIntLLROutputS5xD(151)(4);
  VNStageIntLLRInputS5xD(379)(1) <= CNStageIntLLROutputS5xD(151)(5);
  VNStageIntLLRInputS5xD(50)(2) <= CNStageIntLLROutputS5xD(152)(0);
  VNStageIntLLRInputS5xD(118)(2) <= CNStageIntLLROutputS5xD(152)(1);
  VNStageIntLLRInputS5xD(189)(1) <= CNStageIntLLROutputS5xD(152)(2);
  VNStageIntLLRInputS5xD(249)(0) <= CNStageIntLLROutputS5xD(152)(3);
  VNStageIntLLRInputS5xD(261)(2) <= CNStageIntLLROutputS5xD(152)(4);
  VNStageIntLLRInputS5xD(348)(2) <= CNStageIntLLROutputS5xD(152)(5);
  VNStageIntLLRInputS5xD(49)(2) <= CNStageIntLLROutputS5xD(153)(0);
  VNStageIntLLRInputS5xD(124)(1) <= CNStageIntLLROutputS5xD(153)(1);
  VNStageIntLLRInputS5xD(184)(2) <= CNStageIntLLROutputS5xD(153)(2);
  VNStageIntLLRInputS5xD(196)(2) <= CNStageIntLLROutputS5xD(153)(3);
  VNStageIntLLRInputS5xD(283)(2) <= CNStageIntLLROutputS5xD(153)(4);
  VNStageIntLLRInputS5xD(366)(2) <= CNStageIntLLROutputS5xD(153)(5);
  VNStageIntLLRInputS5xD(48)(1) <= CNStageIntLLROutputS5xD(154)(0);
  VNStageIntLLRInputS5xD(119)(2) <= CNStageIntLLROutputS5xD(154)(1);
  VNStageIntLLRInputS5xD(131)(1) <= CNStageIntLLROutputS5xD(154)(2);
  VNStageIntLLRInputS5xD(218)(2) <= CNStageIntLLROutputS5xD(154)(3);
  VNStageIntLLRInputS5xD(301)(2) <= CNStageIntLLROutputS5xD(154)(4);
  VNStageIntLLRInputS5xD(351)(1) <= CNStageIntLLROutputS5xD(154)(5);
  VNStageIntLLRInputS5xD(47)(1) <= CNStageIntLLROutputS5xD(155)(0);
  VNStageIntLLRInputS5xD(66)(2) <= CNStageIntLLROutputS5xD(155)(1);
  VNStageIntLLRInputS5xD(153)(2) <= CNStageIntLLROutputS5xD(155)(2);
  VNStageIntLLRInputS5xD(236)(2) <= CNStageIntLLROutputS5xD(155)(3);
  VNStageIntLLRInputS5xD(286)(2) <= CNStageIntLLROutputS5xD(155)(4);
  VNStageIntLLRInputS5xD(338)(2) <= CNStageIntLLROutputS5xD(155)(5);
  VNStageIntLLRInputS5xD(46)(2) <= CNStageIntLLROutputS5xD(156)(0);
  VNStageIntLLRInputS5xD(88)(2) <= CNStageIntLLROutputS5xD(156)(1);
  VNStageIntLLRInputS5xD(171)(1) <= CNStageIntLLROutputS5xD(156)(2);
  VNStageIntLLRInputS5xD(221)(2) <= CNStageIntLLROutputS5xD(156)(3);
  VNStageIntLLRInputS5xD(273)(2) <= CNStageIntLLROutputS5xD(156)(4);
  VNStageIntLLRInputS5xD(369)(1) <= CNStageIntLLROutputS5xD(156)(5);
  VNStageIntLLRInputS5xD(45)(2) <= CNStageIntLLROutputS5xD(157)(0);
  VNStageIntLLRInputS5xD(106)(1) <= CNStageIntLLROutputS5xD(157)(1);
  VNStageIntLLRInputS5xD(156)(2) <= CNStageIntLLROutputS5xD(157)(2);
  VNStageIntLLRInputS5xD(208)(2) <= CNStageIntLLROutputS5xD(157)(3);
  VNStageIntLLRInputS5xD(304)(2) <= CNStageIntLLROutputS5xD(157)(4);
  VNStageIntLLRInputS5xD(381)(1) <= CNStageIntLLROutputS5xD(157)(5);
  VNStageIntLLRInputS5xD(44)(2) <= CNStageIntLLROutputS5xD(158)(0);
  VNStageIntLLRInputS5xD(91)(2) <= CNStageIntLLROutputS5xD(158)(1);
  VNStageIntLLRInputS5xD(143)(2) <= CNStageIntLLROutputS5xD(158)(2);
  VNStageIntLLRInputS5xD(239)(2) <= CNStageIntLLROutputS5xD(158)(3);
  VNStageIntLLRInputS5xD(316)(1) <= CNStageIntLLROutputS5xD(158)(4);
  VNStageIntLLRInputS5xD(332)(2) <= CNStageIntLLROutputS5xD(158)(5);
  VNStageIntLLRInputS5xD(43)(1) <= CNStageIntLLROutputS5xD(159)(0);
  VNStageIntLLRInputS5xD(78)(2) <= CNStageIntLLROutputS5xD(159)(1);
  VNStageIntLLRInputS5xD(174)(2) <= CNStageIntLLROutputS5xD(159)(2);
  VNStageIntLLRInputS5xD(251)(1) <= CNStageIntLLROutputS5xD(159)(3);
  VNStageIntLLRInputS5xD(267)(2) <= CNStageIntLLROutputS5xD(159)(4);
  VNStageIntLLRInputS5xD(376)(2) <= CNStageIntLLROutputS5xD(159)(5);
  VNStageIntLLRInputS5xD(42)(2) <= CNStageIntLLROutputS5xD(160)(0);
  VNStageIntLLRInputS5xD(109)(2) <= CNStageIntLLROutputS5xD(160)(1);
  VNStageIntLLRInputS5xD(186)(1) <= CNStageIntLLROutputS5xD(160)(2);
  VNStageIntLLRInputS5xD(202)(2) <= CNStageIntLLROutputS5xD(160)(3);
  VNStageIntLLRInputS5xD(311)(2) <= CNStageIntLLROutputS5xD(160)(4);
  VNStageIntLLRInputS5xD(353)(2) <= CNStageIntLLROutputS5xD(160)(5);
  VNStageIntLLRInputS5xD(41)(2) <= CNStageIntLLROutputS5xD(161)(0);
  VNStageIntLLRInputS5xD(121)(1) <= CNStageIntLLROutputS5xD(161)(1);
  VNStageIntLLRInputS5xD(137)(2) <= CNStageIntLLROutputS5xD(161)(2);
  VNStageIntLLRInputS5xD(246)(2) <= CNStageIntLLROutputS5xD(161)(3);
  VNStageIntLLRInputS5xD(288)(2) <= CNStageIntLLROutputS5xD(161)(4);
  VNStageIntLLRInputS5xD(342)(2) <= CNStageIntLLROutputS5xD(161)(5);
  VNStageIntLLRInputS5xD(40)(2) <= CNStageIntLLROutputS5xD(162)(0);
  VNStageIntLLRInputS5xD(72)(2) <= CNStageIntLLROutputS5xD(162)(1);
  VNStageIntLLRInputS5xD(181)(2) <= CNStageIntLLROutputS5xD(162)(2);
  VNStageIntLLRInputS5xD(223)(2) <= CNStageIntLLROutputS5xD(162)(3);
  VNStageIntLLRInputS5xD(277)(2) <= CNStageIntLLROutputS5xD(162)(4);
  VNStageIntLLRInputS5xD(346)(2) <= CNStageIntLLROutputS5xD(162)(5);
  VNStageIntLLRInputS5xD(39)(2) <= CNStageIntLLROutputS5xD(163)(0);
  VNStageIntLLRInputS5xD(116)(1) <= CNStageIntLLROutputS5xD(163)(1);
  VNStageIntLLRInputS5xD(158)(2) <= CNStageIntLLROutputS5xD(163)(2);
  VNStageIntLLRInputS5xD(212)(2) <= CNStageIntLLROutputS5xD(163)(3);
  VNStageIntLLRInputS5xD(281)(2) <= CNStageIntLLROutputS5xD(163)(4);
  VNStageIntLLRInputS5xD(339)(2) <= CNStageIntLLROutputS5xD(163)(5);
  VNStageIntLLRInputS5xD(38)(2) <= CNStageIntLLROutputS5xD(164)(0);
  VNStageIntLLRInputS5xD(93)(2) <= CNStageIntLLROutputS5xD(164)(1);
  VNStageIntLLRInputS5xD(147)(2) <= CNStageIntLLROutputS5xD(164)(2);
  VNStageIntLLRInputS5xD(216)(2) <= CNStageIntLLROutputS5xD(164)(3);
  VNStageIntLLRInputS5xD(274)(1) <= CNStageIntLLROutputS5xD(164)(4);
  VNStageIntLLRInputS5xD(350)(2) <= CNStageIntLLROutputS5xD(164)(5);
  VNStageIntLLRInputS5xD(37)(2) <= CNStageIntLLROutputS5xD(165)(0);
  VNStageIntLLRInputS5xD(82)(2) <= CNStageIntLLROutputS5xD(165)(1);
  VNStageIntLLRInputS5xD(151)(2) <= CNStageIntLLROutputS5xD(165)(2);
  VNStageIntLLRInputS5xD(209)(2) <= CNStageIntLLROutputS5xD(165)(3);
  VNStageIntLLRInputS5xD(285)(2) <= CNStageIntLLROutputS5xD(165)(4);
  VNStageIntLLRInputS5xD(322)(2) <= CNStageIntLLROutputS5xD(165)(5);
  VNStageIntLLRInputS5xD(36)(2) <= CNStageIntLLROutputS5xD(166)(0);
  VNStageIntLLRInputS5xD(86)(1) <= CNStageIntLLROutputS5xD(166)(1);
  VNStageIntLLRInputS5xD(144)(2) <= CNStageIntLLROutputS5xD(166)(2);
  VNStageIntLLRInputS5xD(220)(2) <= CNStageIntLLROutputS5xD(166)(3);
  VNStageIntLLRInputS5xD(257)(2) <= CNStageIntLLROutputS5xD(166)(4);
  VNStageIntLLRInputS5xD(377)(1) <= CNStageIntLLROutputS5xD(166)(5);
  VNStageIntLLRInputS5xD(35)(2) <= CNStageIntLLROutputS5xD(167)(0);
  VNStageIntLLRInputS5xD(79)(2) <= CNStageIntLLROutputS5xD(167)(1);
  VNStageIntLLRInputS5xD(155)(2) <= CNStageIntLLROutputS5xD(167)(2);
  VNStageIntLLRInputS5xD(255)(2) <= CNStageIntLLROutputS5xD(167)(3);
  VNStageIntLLRInputS5xD(312)(2) <= CNStageIntLLROutputS5xD(167)(4);
  VNStageIntLLRInputS5xD(331)(2) <= CNStageIntLLROutputS5xD(167)(5);
  VNStageIntLLRInputS5xD(34)(2) <= CNStageIntLLROutputS5xD(168)(0);
  VNStageIntLLRInputS5xD(90)(2) <= CNStageIntLLROutputS5xD(168)(1);
  VNStageIntLLRInputS5xD(190)(0) <= CNStageIntLLROutputS5xD(168)(2);
  VNStageIntLLRInputS5xD(247)(2) <= CNStageIntLLROutputS5xD(168)(3);
  VNStageIntLLRInputS5xD(266)(1) <= CNStageIntLLROutputS5xD(168)(4);
  VNStageIntLLRInputS5xD(328)(2) <= CNStageIntLLROutputS5xD(168)(5);
  VNStageIntLLRInputS5xD(33)(2) <= CNStageIntLLROutputS5xD(169)(0);
  VNStageIntLLRInputS5xD(125)(1) <= CNStageIntLLROutputS5xD(169)(1);
  VNStageIntLLRInputS5xD(182)(2) <= CNStageIntLLROutputS5xD(169)(2);
  VNStageIntLLRInputS5xD(201)(2) <= CNStageIntLLROutputS5xD(169)(3);
  VNStageIntLLRInputS5xD(263)(2) <= CNStageIntLLROutputS5xD(169)(4);
  VNStageIntLLRInputS5xD(362)(2) <= CNStageIntLLROutputS5xD(169)(5);
  VNStageIntLLRInputS5xD(0)(2) <= CNStageIntLLROutputS5xD(170)(0);
  VNStageIntLLRInputS5xD(75)(2) <= CNStageIntLLROutputS5xD(170)(1);
  VNStageIntLLRInputS5xD(140)(2) <= CNStageIntLLROutputS5xD(170)(2);
  VNStageIntLLRInputS5xD(205)(0) <= CNStageIntLLROutputS5xD(170)(3);
  VNStageIntLLRInputS5xD(270)(2) <= CNStageIntLLROutputS5xD(170)(4);
  VNStageIntLLRInputS5xD(335)(2) <= CNStageIntLLROutputS5xD(170)(5);
  VNStageIntLLRInputS5xD(62)(2) <= CNStageIntLLROutputS5xD(171)(0);
  VNStageIntLLRInputS5xD(109)(3) <= CNStageIntLLROutputS5xD(171)(1);
  VNStageIntLLRInputS5xD(161)(3) <= CNStageIntLLROutputS5xD(171)(2);
  VNStageIntLLRInputS5xD(194)(3) <= CNStageIntLLROutputS5xD(171)(3);
  VNStageIntLLRInputS5xD(271)(2) <= CNStageIntLLROutputS5xD(171)(4);
  VNStageIntLLRInputS5xD(350)(3) <= CNStageIntLLROutputS5xD(171)(5);
  VNStageIntLLRInputS5xD(61)(2) <= CNStageIntLLROutputS5xD(172)(0);
  VNStageIntLLRInputS5xD(96)(3) <= CNStageIntLLROutputS5xD(172)(1);
  VNStageIntLLRInputS5xD(129)(3) <= CNStageIntLLROutputS5xD(172)(2);
  VNStageIntLLRInputS5xD(206)(2) <= CNStageIntLLROutputS5xD(172)(3);
  VNStageIntLLRInputS5xD(285)(3) <= CNStageIntLLROutputS5xD(172)(4);
  VNStageIntLLRInputS5xD(331)(3) <= CNStageIntLLROutputS5xD(172)(5);
  VNStageIntLLRInputS5xD(60)(2) <= CNStageIntLLROutputS5xD(173)(0);
  VNStageIntLLRInputS5xD(127)(3) <= CNStageIntLLROutputS5xD(173)(1);
  VNStageIntLLRInputS5xD(141)(1) <= CNStageIntLLROutputS5xD(173)(2);
  VNStageIntLLRInputS5xD(220)(3) <= CNStageIntLLROutputS5xD(173)(3);
  VNStageIntLLRInputS5xD(266)(2) <= CNStageIntLLROutputS5xD(173)(4);
  VNStageIntLLRInputS5xD(371)(2) <= CNStageIntLLROutputS5xD(173)(5);
  VNStageIntLLRInputS5xD(59)(1) <= CNStageIntLLROutputS5xD(174)(0);
  VNStageIntLLRInputS5xD(76)(3) <= CNStageIntLLROutputS5xD(174)(1);
  VNStageIntLLRInputS5xD(155)(3) <= CNStageIntLLROutputS5xD(174)(2);
  VNStageIntLLRInputS5xD(201)(3) <= CNStageIntLLROutputS5xD(174)(3);
  VNStageIntLLRInputS5xD(306)(3) <= CNStageIntLLROutputS5xD(174)(4);
  VNStageIntLLRInputS5xD(360)(3) <= CNStageIntLLROutputS5xD(174)(5);
  VNStageIntLLRInputS5xD(58)(2) <= CNStageIntLLROutputS5xD(175)(0);
  VNStageIntLLRInputS5xD(90)(3) <= CNStageIntLLROutputS5xD(175)(1);
  VNStageIntLLRInputS5xD(136)(3) <= CNStageIntLLROutputS5xD(175)(2);
  VNStageIntLLRInputS5xD(241)(2) <= CNStageIntLLROutputS5xD(175)(3);
  VNStageIntLLRInputS5xD(295)(3) <= CNStageIntLLROutputS5xD(175)(4);
  VNStageIntLLRInputS5xD(364)(3) <= CNStageIntLLROutputS5xD(175)(5);
  VNStageIntLLRInputS5xD(57)(2) <= CNStageIntLLROutputS5xD(176)(0);
  VNStageIntLLRInputS5xD(71)(2) <= CNStageIntLLROutputS5xD(176)(1);
  VNStageIntLLRInputS5xD(176)(3) <= CNStageIntLLROutputS5xD(176)(2);
  VNStageIntLLRInputS5xD(230)(2) <= CNStageIntLLROutputS5xD(176)(3);
  VNStageIntLLRInputS5xD(299)(2) <= CNStageIntLLROutputS5xD(176)(4);
  VNStageIntLLRInputS5xD(357)(3) <= CNStageIntLLROutputS5xD(176)(5);
  VNStageIntLLRInputS5xD(56)(3) <= CNStageIntLLROutputS5xD(177)(0);
  VNStageIntLLRInputS5xD(111)(3) <= CNStageIntLLROutputS5xD(177)(1);
  VNStageIntLLRInputS5xD(165)(3) <= CNStageIntLLROutputS5xD(177)(2);
  VNStageIntLLRInputS5xD(234)(3) <= CNStageIntLLROutputS5xD(177)(3);
  VNStageIntLLRInputS5xD(292)(3) <= CNStageIntLLROutputS5xD(177)(4);
  VNStageIntLLRInputS5xD(368)(1) <= CNStageIntLLROutputS5xD(177)(5);
  VNStageIntLLRInputS5xD(55)(3) <= CNStageIntLLROutputS5xD(178)(0);
  VNStageIntLLRInputS5xD(100)(3) <= CNStageIntLLROutputS5xD(178)(1);
  VNStageIntLLRInputS5xD(169)(3) <= CNStageIntLLROutputS5xD(178)(2);
  VNStageIntLLRInputS5xD(227)(3) <= CNStageIntLLROutputS5xD(178)(3);
  VNStageIntLLRInputS5xD(303)(3) <= CNStageIntLLROutputS5xD(178)(4);
  VNStageIntLLRInputS5xD(340)(3) <= CNStageIntLLROutputS5xD(178)(5);
  VNStageIntLLRInputS5xD(54)(3) <= CNStageIntLLROutputS5xD(179)(0);
  VNStageIntLLRInputS5xD(104)(3) <= CNStageIntLLROutputS5xD(179)(1);
  VNStageIntLLRInputS5xD(162)(3) <= CNStageIntLLROutputS5xD(179)(2);
  VNStageIntLLRInputS5xD(238)(3) <= CNStageIntLLROutputS5xD(179)(3);
  VNStageIntLLRInputS5xD(275)(3) <= CNStageIntLLROutputS5xD(179)(4);
  VNStageIntLLRInputS5xD(332)(3) <= CNStageIntLLROutputS5xD(179)(5);
  VNStageIntLLRInputS5xD(53)(2) <= CNStageIntLLROutputS5xD(180)(0);
  VNStageIntLLRInputS5xD(97)(3) <= CNStageIntLLROutputS5xD(180)(1);
  VNStageIntLLRInputS5xD(173)(3) <= CNStageIntLLROutputS5xD(180)(2);
  VNStageIntLLRInputS5xD(210)(3) <= CNStageIntLLROutputS5xD(180)(3);
  VNStageIntLLRInputS5xD(267)(3) <= CNStageIntLLROutputS5xD(180)(4);
  VNStageIntLLRInputS5xD(349)(2) <= CNStageIntLLROutputS5xD(180)(5);
  VNStageIntLLRInputS5xD(52)(2) <= CNStageIntLLROutputS5xD(181)(0);
  VNStageIntLLRInputS5xD(108)(3) <= CNStageIntLLROutputS5xD(181)(1);
  VNStageIntLLRInputS5xD(145)(3) <= CNStageIntLLROutputS5xD(181)(2);
  VNStageIntLLRInputS5xD(202)(3) <= CNStageIntLLROutputS5xD(181)(3);
  VNStageIntLLRInputS5xD(284)(3) <= CNStageIntLLROutputS5xD(181)(4);
  VNStageIntLLRInputS5xD(346)(3) <= CNStageIntLLROutputS5xD(181)(5);
  VNStageIntLLRInputS5xD(51)(2) <= CNStageIntLLROutputS5xD(182)(0);
  VNStageIntLLRInputS5xD(80)(3) <= CNStageIntLLROutputS5xD(182)(1);
  VNStageIntLLRInputS5xD(137)(3) <= CNStageIntLLROutputS5xD(182)(2);
  VNStageIntLLRInputS5xD(219)(3) <= CNStageIntLLROutputS5xD(182)(3);
  VNStageIntLLRInputS5xD(281)(3) <= CNStageIntLLROutputS5xD(182)(4);
  VNStageIntLLRInputS5xD(380)(2) <= CNStageIntLLROutputS5xD(182)(5);
  VNStageIntLLRInputS5xD(50)(3) <= CNStageIntLLROutputS5xD(183)(0);
  VNStageIntLLRInputS5xD(72)(3) <= CNStageIntLLROutputS5xD(183)(1);
  VNStageIntLLRInputS5xD(154)(2) <= CNStageIntLLROutputS5xD(183)(2);
  VNStageIntLLRInputS5xD(216)(3) <= CNStageIntLLROutputS5xD(183)(3);
  VNStageIntLLRInputS5xD(315)(2) <= CNStageIntLLROutputS5xD(183)(4);
  VNStageIntLLRInputS5xD(337)(3) <= CNStageIntLLROutputS5xD(183)(5);
  VNStageIntLLRInputS5xD(49)(3) <= CNStageIntLLROutputS5xD(184)(0);
  VNStageIntLLRInputS5xD(89)(3) <= CNStageIntLLROutputS5xD(184)(1);
  VNStageIntLLRInputS5xD(151)(3) <= CNStageIntLLROutputS5xD(184)(2);
  VNStageIntLLRInputS5xD(250)(2) <= CNStageIntLLROutputS5xD(184)(3);
  VNStageIntLLRInputS5xD(272)(3) <= CNStageIntLLROutputS5xD(184)(4);
  VNStageIntLLRInputS5xD(323)(2) <= CNStageIntLLROutputS5xD(184)(5);
  VNStageIntLLRInputS5xD(46)(3) <= CNStageIntLLROutputS5xD(185)(0);
  VNStageIntLLRInputS5xD(77)(1) <= CNStageIntLLROutputS5xD(185)(1);
  VNStageIntLLRInputS5xD(191)(3) <= CNStageIntLLROutputS5xD(185)(2);
  VNStageIntLLRInputS5xD(246)(3) <= CNStageIntLLROutputS5xD(185)(3);
  VNStageIntLLRInputS5xD(277)(3) <= CNStageIntLLROutputS5xD(185)(4);
  VNStageIntLLRInputS5xD(325)(3) <= CNStageIntLLROutputS5xD(185)(5);
  VNStageIntLLRInputS5xD(45)(3) <= CNStageIntLLROutputS5xD(186)(0);
  VNStageIntLLRInputS5xD(126)(2) <= CNStageIntLLROutputS5xD(186)(1);
  VNStageIntLLRInputS5xD(181)(3) <= CNStageIntLLROutputS5xD(186)(2);
  VNStageIntLLRInputS5xD(212)(3) <= CNStageIntLLROutputS5xD(186)(3);
  VNStageIntLLRInputS5xD(260)(3) <= CNStageIntLLROutputS5xD(186)(4);
  VNStageIntLLRInputS5xD(355)(3) <= CNStageIntLLROutputS5xD(186)(5);
  VNStageIntLLRInputS5xD(44)(3) <= CNStageIntLLROutputS5xD(187)(0);
  VNStageIntLLRInputS5xD(116)(2) <= CNStageIntLLROutputS5xD(187)(1);
  VNStageIntLLRInputS5xD(147)(3) <= CNStageIntLLROutputS5xD(187)(2);
  VNStageIntLLRInputS5xD(195)(2) <= CNStageIntLLROutputS5xD(187)(3);
  VNStageIntLLRInputS5xD(290)(3) <= CNStageIntLLROutputS5xD(187)(4);
  VNStageIntLLRInputS5xD(378)(2) <= CNStageIntLLROutputS5xD(187)(5);
  VNStageIntLLRInputS5xD(43)(2) <= CNStageIntLLROutputS5xD(188)(0);
  VNStageIntLLRInputS5xD(82)(3) <= CNStageIntLLROutputS5xD(188)(1);
  VNStageIntLLRInputS5xD(130)(3) <= CNStageIntLLROutputS5xD(188)(2);
  VNStageIntLLRInputS5xD(225)(3) <= CNStageIntLLROutputS5xD(188)(3);
  VNStageIntLLRInputS5xD(313)(1) <= CNStageIntLLROutputS5xD(188)(4);
  VNStageIntLLRInputS5xD(351)(2) <= CNStageIntLLROutputS5xD(188)(5);
  VNStageIntLLRInputS5xD(42)(3) <= CNStageIntLLROutputS5xD(189)(0);
  VNStageIntLLRInputS5xD(65)(3) <= CNStageIntLLROutputS5xD(189)(1);
  VNStageIntLLRInputS5xD(160)(3) <= CNStageIntLLROutputS5xD(189)(2);
  VNStageIntLLRInputS5xD(248)(3) <= CNStageIntLLROutputS5xD(189)(3);
  VNStageIntLLRInputS5xD(286)(3) <= CNStageIntLLROutputS5xD(189)(4);
  VNStageIntLLRInputS5xD(335)(3) <= CNStageIntLLROutputS5xD(189)(5);
  VNStageIntLLRInputS5xD(41)(3) <= CNStageIntLLROutputS5xD(190)(0);
  VNStageIntLLRInputS5xD(95)(3) <= CNStageIntLLROutputS5xD(190)(1);
  VNStageIntLLRInputS5xD(183)(2) <= CNStageIntLLROutputS5xD(190)(2);
  VNStageIntLLRInputS5xD(221)(3) <= CNStageIntLLROutputS5xD(190)(3);
  VNStageIntLLRInputS5xD(270)(3) <= CNStageIntLLROutputS5xD(190)(4);
  VNStageIntLLRInputS5xD(338)(3) <= CNStageIntLLROutputS5xD(190)(5);
  VNStageIntLLRInputS5xD(39)(3) <= CNStageIntLLROutputS5xD(191)(0);
  VNStageIntLLRInputS5xD(91)(3) <= CNStageIntLLROutputS5xD(191)(1);
  VNStageIntLLRInputS5xD(140)(3) <= CNStageIntLLROutputS5xD(191)(2);
  VNStageIntLLRInputS5xD(208)(3) <= CNStageIntLLROutputS5xD(191)(3);
  VNStageIntLLRInputS5xD(314)(0) <= CNStageIntLLROutputS5xD(191)(4);
  VNStageIntLLRInputS5xD(354)(3) <= CNStageIntLLROutputS5xD(191)(5);
  VNStageIntLLRInputS5xD(38)(3) <= CNStageIntLLROutputS5xD(192)(0);
  VNStageIntLLRInputS5xD(75)(3) <= CNStageIntLLROutputS5xD(192)(1);
  VNStageIntLLRInputS5xD(143)(3) <= CNStageIntLLROutputS5xD(192)(2);
  VNStageIntLLRInputS5xD(249)(1) <= CNStageIntLLROutputS5xD(192)(3);
  VNStageIntLLRInputS5xD(289)(3) <= CNStageIntLLROutputS5xD(192)(4);
  VNStageIntLLRInputS5xD(352)(3) <= CNStageIntLLROutputS5xD(192)(5);
  VNStageIntLLRInputS5xD(37)(3) <= CNStageIntLLROutputS5xD(193)(0);
  VNStageIntLLRInputS5xD(78)(3) <= CNStageIntLLROutputS5xD(193)(1);
  VNStageIntLLRInputS5xD(184)(3) <= CNStageIntLLROutputS5xD(193)(2);
  VNStageIntLLRInputS5xD(224)(3) <= CNStageIntLLROutputS5xD(193)(3);
  VNStageIntLLRInputS5xD(287)(3) <= CNStageIntLLROutputS5xD(193)(4);
  VNStageIntLLRInputS5xD(377)(2) <= CNStageIntLLROutputS5xD(193)(5);
  VNStageIntLLRInputS5xD(35)(3) <= CNStageIntLLROutputS5xD(194)(0);
  VNStageIntLLRInputS5xD(94)(2) <= CNStageIntLLROutputS5xD(194)(1);
  VNStageIntLLRInputS5xD(157)(3) <= CNStageIntLLROutputS5xD(194)(2);
  VNStageIntLLRInputS5xD(247)(3) <= CNStageIntLLROutputS5xD(194)(3);
  VNStageIntLLRInputS5xD(257)(3) <= CNStageIntLLROutputS5xD(194)(4);
  VNStageIntLLRInputS5xD(365)(3) <= CNStageIntLLROutputS5xD(194)(5);
  VNStageIntLLRInputS5xD(34)(3) <= CNStageIntLLROutputS5xD(195)(0);
  VNStageIntLLRInputS5xD(92)(3) <= CNStageIntLLROutputS5xD(195)(1);
  VNStageIntLLRInputS5xD(182)(3) <= CNStageIntLLROutputS5xD(195)(2);
  VNStageIntLLRInputS5xD(255)(3) <= CNStageIntLLROutputS5xD(195)(3);
  VNStageIntLLRInputS5xD(300)(3) <= CNStageIntLLROutputS5xD(195)(4);
  VNStageIntLLRInputS5xD(359)(3) <= CNStageIntLLROutputS5xD(195)(5);
  VNStageIntLLRInputS5xD(33)(3) <= CNStageIntLLROutputS5xD(196)(0);
  VNStageIntLLRInputS5xD(117)(3) <= CNStageIntLLROutputS5xD(196)(1);
  VNStageIntLLRInputS5xD(190)(1) <= CNStageIntLLROutputS5xD(196)(2);
  VNStageIntLLRInputS5xD(235)(2) <= CNStageIntLLROutputS5xD(196)(3);
  VNStageIntLLRInputS5xD(294)(3) <= CNStageIntLLROutputS5xD(196)(4);
  VNStageIntLLRInputS5xD(320)(2) <= CNStageIntLLROutputS5xD(196)(5);
  VNStageIntLLRInputS5xD(31)(2) <= CNStageIntLLROutputS5xD(197)(0);
  VNStageIntLLRInputS5xD(105)(2) <= CNStageIntLLROutputS5xD(197)(1);
  VNStageIntLLRInputS5xD(164)(3) <= CNStageIntLLROutputS5xD(197)(2);
  VNStageIntLLRInputS5xD(192)(3) <= CNStageIntLLROutputS5xD(197)(3);
  VNStageIntLLRInputS5xD(293)(3) <= CNStageIntLLROutputS5xD(197)(4);
  VNStageIntLLRInputS5xD(363)(2) <= CNStageIntLLROutputS5xD(197)(5);
  VNStageIntLLRInputS5xD(30)(3) <= CNStageIntLLROutputS5xD(198)(0);
  VNStageIntLLRInputS5xD(99)(3) <= CNStageIntLLROutputS5xD(198)(1);
  VNStageIntLLRInputS5xD(128)(3) <= CNStageIntLLROutputS5xD(198)(2);
  VNStageIntLLRInputS5xD(228)(3) <= CNStageIntLLROutputS5xD(198)(3);
  VNStageIntLLRInputS5xD(298)(3) <= CNStageIntLLROutputS5xD(198)(4);
  VNStageIntLLRInputS5xD(382)(2) <= CNStageIntLLROutputS5xD(198)(5);
  VNStageIntLLRInputS5xD(28)(3) <= CNStageIntLLROutputS5xD(199)(0);
  VNStageIntLLRInputS5xD(98)(2) <= CNStageIntLLROutputS5xD(199)(1);
  VNStageIntLLRInputS5xD(168)(2) <= CNStageIntLLROutputS5xD(199)(2);
  VNStageIntLLRInputS5xD(252)(2) <= CNStageIntLLROutputS5xD(199)(3);
  VNStageIntLLRInputS5xD(308)(1) <= CNStageIntLLROutputS5xD(199)(4);
  VNStageIntLLRInputS5xD(347)(3) <= CNStageIntLLROutputS5xD(199)(5);
  VNStageIntLLRInputS5xD(27)(3) <= CNStageIntLLROutputS5xD(200)(0);
  VNStageIntLLRInputS5xD(103)(3) <= CNStageIntLLROutputS5xD(200)(1);
  VNStageIntLLRInputS5xD(187)(2) <= CNStageIntLLROutputS5xD(200)(2);
  VNStageIntLLRInputS5xD(243)(3) <= CNStageIntLLROutputS5xD(200)(3);
  VNStageIntLLRInputS5xD(282)(3) <= CNStageIntLLROutputS5xD(200)(4);
  VNStageIntLLRInputS5xD(348)(3) <= CNStageIntLLROutputS5xD(200)(5);
  VNStageIntLLRInputS5xD(26)(3) <= CNStageIntLLROutputS5xD(201)(0);
  VNStageIntLLRInputS5xD(122)(2) <= CNStageIntLLROutputS5xD(201)(1);
  VNStageIntLLRInputS5xD(178)(3) <= CNStageIntLLROutputS5xD(201)(2);
  VNStageIntLLRInputS5xD(217)(3) <= CNStageIntLLROutputS5xD(201)(3);
  VNStageIntLLRInputS5xD(283)(3) <= CNStageIntLLROutputS5xD(201)(4);
  VNStageIntLLRInputS5xD(372)(2) <= CNStageIntLLROutputS5xD(201)(5);
  VNStageIntLLRInputS5xD(25)(3) <= CNStageIntLLROutputS5xD(202)(0);
  VNStageIntLLRInputS5xD(113)(3) <= CNStageIntLLROutputS5xD(202)(1);
  VNStageIntLLRInputS5xD(152)(3) <= CNStageIntLLROutputS5xD(202)(2);
  VNStageIntLLRInputS5xD(218)(3) <= CNStageIntLLROutputS5xD(202)(3);
  VNStageIntLLRInputS5xD(307)(3) <= CNStageIntLLROutputS5xD(202)(4);
  VNStageIntLLRInputS5xD(330)(3) <= CNStageIntLLROutputS5xD(202)(5);
  VNStageIntLLRInputS5xD(24)(3) <= CNStageIntLLROutputS5xD(203)(0);
  VNStageIntLLRInputS5xD(87)(3) <= CNStageIntLLROutputS5xD(203)(1);
  VNStageIntLLRInputS5xD(153)(3) <= CNStageIntLLROutputS5xD(203)(2);
  VNStageIntLLRInputS5xD(242)(3) <= CNStageIntLLROutputS5xD(203)(3);
  VNStageIntLLRInputS5xD(265)(2) <= CNStageIntLLROutputS5xD(203)(4);
  VNStageIntLLRInputS5xD(326)(2) <= CNStageIntLLROutputS5xD(203)(5);
  VNStageIntLLRInputS5xD(23)(3) <= CNStageIntLLROutputS5xD(204)(0);
  VNStageIntLLRInputS5xD(88)(3) <= CNStageIntLLROutputS5xD(204)(1);
  VNStageIntLLRInputS5xD(177)(3) <= CNStageIntLLROutputS5xD(204)(2);
  VNStageIntLLRInputS5xD(200)(3) <= CNStageIntLLROutputS5xD(204)(3);
  VNStageIntLLRInputS5xD(261)(3) <= CNStageIntLLROutputS5xD(204)(4);
  VNStageIntLLRInputS5xD(341)(3) <= CNStageIntLLROutputS5xD(204)(5);
  VNStageIntLLRInputS5xD(22)(3) <= CNStageIntLLROutputS5xD(205)(0);
  VNStageIntLLRInputS5xD(112)(3) <= CNStageIntLLROutputS5xD(205)(1);
  VNStageIntLLRInputS5xD(135)(3) <= CNStageIntLLROutputS5xD(205)(2);
  VNStageIntLLRInputS5xD(196)(3) <= CNStageIntLLROutputS5xD(205)(3);
  VNStageIntLLRInputS5xD(276)(3) <= CNStageIntLLROutputS5xD(205)(4);
  VNStageIntLLRInputS5xD(367)(3) <= CNStageIntLLROutputS5xD(205)(5);
  VNStageIntLLRInputS5xD(21)(3) <= CNStageIntLLROutputS5xD(206)(0);
  VNStageIntLLRInputS5xD(70)(3) <= CNStageIntLLROutputS5xD(206)(1);
  VNStageIntLLRInputS5xD(131)(2) <= CNStageIntLLROutputS5xD(206)(2);
  VNStageIntLLRInputS5xD(211)(3) <= CNStageIntLLROutputS5xD(206)(3);
  VNStageIntLLRInputS5xD(302)(3) <= CNStageIntLLROutputS5xD(206)(4);
  VNStageIntLLRInputS5xD(343)(3) <= CNStageIntLLROutputS5xD(206)(5);
  VNStageIntLLRInputS5xD(18)(3) <= CNStageIntLLROutputS5xD(207)(0);
  VNStageIntLLRInputS5xD(107)(2) <= CNStageIntLLROutputS5xD(207)(1);
  VNStageIntLLRInputS5xD(148)(3) <= CNStageIntLLROutputS5xD(207)(2);
  VNStageIntLLRInputS5xD(245)(3) <= CNStageIntLLROutputS5xD(207)(3);
  VNStageIntLLRInputS5xD(263)(3) <= CNStageIntLLROutputS5xD(207)(4);
  VNStageIntLLRInputS5xD(361)(3) <= CNStageIntLLROutputS5xD(207)(5);
  VNStageIntLLRInputS5xD(17)(3) <= CNStageIntLLROutputS5xD(208)(0);
  VNStageIntLLRInputS5xD(83)(3) <= CNStageIntLLROutputS5xD(208)(1);
  VNStageIntLLRInputS5xD(180)(1) <= CNStageIntLLROutputS5xD(208)(2);
  VNStageIntLLRInputS5xD(198)(3) <= CNStageIntLLROutputS5xD(208)(3);
  VNStageIntLLRInputS5xD(296)(3) <= CNStageIntLLROutputS5xD(208)(4);
  VNStageIntLLRInputS5xD(370)(2) <= CNStageIntLLROutputS5xD(208)(5);
  VNStageIntLLRInputS5xD(16)(2) <= CNStageIntLLROutputS5xD(209)(0);
  VNStageIntLLRInputS5xD(115)(3) <= CNStageIntLLROutputS5xD(209)(1);
  VNStageIntLLRInputS5xD(133)(1) <= CNStageIntLLROutputS5xD(209)(2);
  VNStageIntLLRInputS5xD(231)(2) <= CNStageIntLLROutputS5xD(209)(3);
  VNStageIntLLRInputS5xD(305)(3) <= CNStageIntLLROutputS5xD(209)(4);
  VNStageIntLLRInputS5xD(383)(3) <= CNStageIntLLROutputS5xD(209)(5);
  VNStageIntLLRInputS5xD(15)(3) <= CNStageIntLLROutputS5xD(210)(0);
  VNStageIntLLRInputS5xD(68)(2) <= CNStageIntLLROutputS5xD(210)(1);
  VNStageIntLLRInputS5xD(166)(3) <= CNStageIntLLROutputS5xD(210)(2);
  VNStageIntLLRInputS5xD(240)(3) <= CNStageIntLLROutputS5xD(210)(3);
  VNStageIntLLRInputS5xD(318)(1) <= CNStageIntLLROutputS5xD(210)(4);
  VNStageIntLLRInputS5xD(362)(3) <= CNStageIntLLROutputS5xD(210)(5);
  VNStageIntLLRInputS5xD(14)(3) <= CNStageIntLLROutputS5xD(211)(0);
  VNStageIntLLRInputS5xD(101)(3) <= CNStageIntLLROutputS5xD(211)(1);
  VNStageIntLLRInputS5xD(175)(3) <= CNStageIntLLROutputS5xD(211)(2);
  VNStageIntLLRInputS5xD(253)(2) <= CNStageIntLLROutputS5xD(211)(3);
  VNStageIntLLRInputS5xD(297)(3) <= CNStageIntLLROutputS5xD(211)(4);
  VNStageIntLLRInputS5xD(327)(3) <= CNStageIntLLROutputS5xD(211)(5);
  VNStageIntLLRInputS5xD(13)(2) <= CNStageIntLLROutputS5xD(212)(0);
  VNStageIntLLRInputS5xD(110)(3) <= CNStageIntLLROutputS5xD(212)(1);
  VNStageIntLLRInputS5xD(188)(1) <= CNStageIntLLROutputS5xD(212)(2);
  VNStageIntLLRInputS5xD(232)(2) <= CNStageIntLLROutputS5xD(212)(3);
  VNStageIntLLRInputS5xD(262)(3) <= CNStageIntLLROutputS5xD(212)(4);
  VNStageIntLLRInputS5xD(329)(3) <= CNStageIntLLROutputS5xD(212)(5);
  VNStageIntLLRInputS5xD(12)(3) <= CNStageIntLLROutputS5xD(213)(0);
  VNStageIntLLRInputS5xD(123)(2) <= CNStageIntLLROutputS5xD(213)(1);
  VNStageIntLLRInputS5xD(167)(3) <= CNStageIntLLROutputS5xD(213)(2);
  VNStageIntLLRInputS5xD(197)(3) <= CNStageIntLLROutputS5xD(213)(3);
  VNStageIntLLRInputS5xD(264)(3) <= CNStageIntLLROutputS5xD(213)(4);
  VNStageIntLLRInputS5xD(374)(3) <= CNStageIntLLROutputS5xD(213)(5);
  VNStageIntLLRInputS5xD(11)(3) <= CNStageIntLLROutputS5xD(214)(0);
  VNStageIntLLRInputS5xD(102)(3) <= CNStageIntLLROutputS5xD(214)(1);
  VNStageIntLLRInputS5xD(132)(2) <= CNStageIntLLROutputS5xD(214)(2);
  VNStageIntLLRInputS5xD(199)(3) <= CNStageIntLLROutputS5xD(214)(3);
  VNStageIntLLRInputS5xD(309)(3) <= CNStageIntLLROutputS5xD(214)(4);
  VNStageIntLLRInputS5xD(381)(2) <= CNStageIntLLROutputS5xD(214)(5);
  VNStageIntLLRInputS5xD(9)(3) <= CNStageIntLLROutputS5xD(215)(0);
  VNStageIntLLRInputS5xD(69)(3) <= CNStageIntLLROutputS5xD(215)(1);
  VNStageIntLLRInputS5xD(179)(3) <= CNStageIntLLROutputS5xD(215)(2);
  VNStageIntLLRInputS5xD(251)(2) <= CNStageIntLLROutputS5xD(215)(3);
  VNStageIntLLRInputS5xD(280)(3) <= CNStageIntLLROutputS5xD(215)(4);
  VNStageIntLLRInputS5xD(333)(2) <= CNStageIntLLROutputS5xD(215)(5);
  VNStageIntLLRInputS5xD(8)(2) <= CNStageIntLLROutputS5xD(216)(0);
  VNStageIntLLRInputS5xD(114)(3) <= CNStageIntLLROutputS5xD(216)(1);
  VNStageIntLLRInputS5xD(186)(2) <= CNStageIntLLROutputS5xD(216)(2);
  VNStageIntLLRInputS5xD(215)(3) <= CNStageIntLLROutputS5xD(216)(3);
  VNStageIntLLRInputS5xD(268)(3) <= CNStageIntLLROutputS5xD(216)(4);
  VNStageIntLLRInputS5xD(339)(3) <= CNStageIntLLROutputS5xD(216)(5);
  VNStageIntLLRInputS5xD(7)(3) <= CNStageIntLLROutputS5xD(217)(0);
  VNStageIntLLRInputS5xD(121)(2) <= CNStageIntLLROutputS5xD(217)(1);
  VNStageIntLLRInputS5xD(150)(3) <= CNStageIntLLROutputS5xD(217)(2);
  VNStageIntLLRInputS5xD(203)(3) <= CNStageIntLLROutputS5xD(217)(3);
  VNStageIntLLRInputS5xD(274)(2) <= CNStageIntLLROutputS5xD(217)(4);
  VNStageIntLLRInputS5xD(334)(2) <= CNStageIntLLROutputS5xD(217)(5);
  VNStageIntLLRInputS5xD(6)(3) <= CNStageIntLLROutputS5xD(218)(0);
  VNStageIntLLRInputS5xD(85)(2) <= CNStageIntLLROutputS5xD(218)(1);
  VNStageIntLLRInputS5xD(138)(3) <= CNStageIntLLROutputS5xD(218)(2);
  VNStageIntLLRInputS5xD(209)(3) <= CNStageIntLLROutputS5xD(218)(3);
  VNStageIntLLRInputS5xD(269)(2) <= CNStageIntLLROutputS5xD(218)(4);
  VNStageIntLLRInputS5xD(344)(3) <= CNStageIntLLROutputS5xD(218)(5);
  VNStageIntLLRInputS5xD(5)(3) <= CNStageIntLLROutputS5xD(219)(0);
  VNStageIntLLRInputS5xD(73)(3) <= CNStageIntLLROutputS5xD(219)(1);
  VNStageIntLLRInputS5xD(144)(3) <= CNStageIntLLROutputS5xD(219)(2);
  VNStageIntLLRInputS5xD(204)(3) <= CNStageIntLLROutputS5xD(219)(3);
  VNStageIntLLRInputS5xD(279)(3) <= CNStageIntLLROutputS5xD(219)(4);
  VNStageIntLLRInputS5xD(366)(3) <= CNStageIntLLROutputS5xD(219)(5);
  VNStageIntLLRInputS5xD(4)(2) <= CNStageIntLLROutputS5xD(220)(0);
  VNStageIntLLRInputS5xD(79)(3) <= CNStageIntLLROutputS5xD(220)(1);
  VNStageIntLLRInputS5xD(139)(3) <= CNStageIntLLROutputS5xD(220)(2);
  VNStageIntLLRInputS5xD(214)(3) <= CNStageIntLLROutputS5xD(220)(3);
  VNStageIntLLRInputS5xD(301)(3) <= CNStageIntLLROutputS5xD(220)(4);
  VNStageIntLLRInputS5xD(321)(3) <= CNStageIntLLROutputS5xD(220)(5);
  VNStageIntLLRInputS5xD(3)(2) <= CNStageIntLLROutputS5xD(221)(0);
  VNStageIntLLRInputS5xD(74)(3) <= CNStageIntLLROutputS5xD(221)(1);
  VNStageIntLLRInputS5xD(149)(3) <= CNStageIntLLROutputS5xD(221)(2);
  VNStageIntLLRInputS5xD(236)(3) <= CNStageIntLLROutputS5xD(221)(3);
  VNStageIntLLRInputS5xD(319)(3) <= CNStageIntLLROutputS5xD(221)(4);
  VNStageIntLLRInputS5xD(369)(2) <= CNStageIntLLROutputS5xD(221)(5);
  VNStageIntLLRInputS5xD(2)(3) <= CNStageIntLLROutputS5xD(222)(0);
  VNStageIntLLRInputS5xD(84)(3) <= CNStageIntLLROutputS5xD(222)(1);
  VNStageIntLLRInputS5xD(171)(2) <= CNStageIntLLROutputS5xD(222)(2);
  VNStageIntLLRInputS5xD(254)(1) <= CNStageIntLLROutputS5xD(222)(3);
  VNStageIntLLRInputS5xD(304)(3) <= CNStageIntLLROutputS5xD(222)(4);
  VNStageIntLLRInputS5xD(356)(3) <= CNStageIntLLROutputS5xD(222)(5);
  VNStageIntLLRInputS5xD(1)(2) <= CNStageIntLLROutputS5xD(223)(0);
  VNStageIntLLRInputS5xD(106)(2) <= CNStageIntLLROutputS5xD(223)(1);
  VNStageIntLLRInputS5xD(189)(2) <= CNStageIntLLROutputS5xD(223)(2);
  VNStageIntLLRInputS5xD(239)(3) <= CNStageIntLLROutputS5xD(223)(3);
  VNStageIntLLRInputS5xD(291)(3) <= CNStageIntLLROutputS5xD(223)(4);
  VNStageIntLLRInputS5xD(324)(3) <= CNStageIntLLROutputS5xD(223)(5);
  VNStageIntLLRInputS5xD(0)(3) <= CNStageIntLLROutputS5xD(224)(0);
  VNStageIntLLRInputS5xD(93)(3) <= CNStageIntLLROutputS5xD(224)(1);
  VNStageIntLLRInputS5xD(158)(3) <= CNStageIntLLROutputS5xD(224)(2);
  VNStageIntLLRInputS5xD(223)(3) <= CNStageIntLLROutputS5xD(224)(3);
  VNStageIntLLRInputS5xD(288)(3) <= CNStageIntLLROutputS5xD(224)(4);
  VNStageIntLLRInputS5xD(353)(3) <= CNStageIntLLROutputS5xD(224)(5);
  VNStageIntLLRInputS5xD(18)(4) <= CNStageIntLLROutputS5xD(225)(0);
  VNStageIntLLRInputS5xD(110)(4) <= CNStageIntLLROutputS5xD(225)(1);
  VNStageIntLLRInputS5xD(167)(4) <= CNStageIntLLROutputS5xD(225)(2);
  VNStageIntLLRInputS5xD(249)(2) <= CNStageIntLLROutputS5xD(225)(3);
  VNStageIntLLRInputS5xD(311)(3) <= CNStageIntLLROutputS5xD(225)(4);
  VNStageIntLLRInputS5xD(347)(4) <= CNStageIntLLROutputS5xD(225)(5);
  VNStageIntLLRInputS5xD(17)(4) <= CNStageIntLLROutputS5xD(226)(0);
  VNStageIntLLRInputS5xD(102)(4) <= CNStageIntLLROutputS5xD(226)(1);
  VNStageIntLLRInputS5xD(184)(4) <= CNStageIntLLROutputS5xD(226)(2);
  VNStageIntLLRInputS5xD(246)(4) <= CNStageIntLLROutputS5xD(226)(3);
  VNStageIntLLRInputS5xD(282)(4) <= CNStageIntLLROutputS5xD(226)(4);
  VNStageIntLLRInputS5xD(367)(4) <= CNStageIntLLROutputS5xD(226)(5);
  VNStageIntLLRInputS5xD(16)(3) <= CNStageIntLLROutputS5xD(227)(0);
  VNStageIntLLRInputS5xD(119)(3) <= CNStageIntLLROutputS5xD(227)(1);
  VNStageIntLLRInputS5xD(181)(4) <= CNStageIntLLROutputS5xD(227)(2);
  VNStageIntLLRInputS5xD(217)(4) <= CNStageIntLLROutputS5xD(227)(3);
  VNStageIntLLRInputS5xD(302)(4) <= CNStageIntLLROutputS5xD(227)(4);
  VNStageIntLLRInputS5xD(353)(4) <= CNStageIntLLROutputS5xD(227)(5);
  VNStageIntLLRInputS5xD(15)(4) <= CNStageIntLLROutputS5xD(228)(0);
  VNStageIntLLRInputS5xD(116)(3) <= CNStageIntLLROutputS5xD(228)(1);
  VNStageIntLLRInputS5xD(152)(4) <= CNStageIntLLROutputS5xD(228)(2);
  VNStageIntLLRInputS5xD(237)(3) <= CNStageIntLLROutputS5xD(228)(3);
  VNStageIntLLRInputS5xD(288)(4) <= CNStageIntLLROutputS5xD(228)(4);
  VNStageIntLLRInputS5xD(343)(4) <= CNStageIntLLROutputS5xD(228)(5);
  VNStageIntLLRInputS5xD(14)(4) <= CNStageIntLLROutputS5xD(229)(0);
  VNStageIntLLRInputS5xD(87)(4) <= CNStageIntLLROutputS5xD(229)(1);
  VNStageIntLLRInputS5xD(172)(3) <= CNStageIntLLROutputS5xD(229)(2);
  VNStageIntLLRInputS5xD(223)(4) <= CNStageIntLLROutputS5xD(229)(3);
  VNStageIntLLRInputS5xD(278)(3) <= CNStageIntLLROutputS5xD(229)(4);
  VNStageIntLLRInputS5xD(372)(3) <= CNStageIntLLROutputS5xD(229)(5);
  VNStageIntLLRInputS5xD(13)(3) <= CNStageIntLLROutputS5xD(230)(0);
  VNStageIntLLRInputS5xD(107)(3) <= CNStageIntLLROutputS5xD(230)(1);
  VNStageIntLLRInputS5xD(158)(4) <= CNStageIntLLROutputS5xD(230)(2);
  VNStageIntLLRInputS5xD(213)(3) <= CNStageIntLLROutputS5xD(230)(3);
  VNStageIntLLRInputS5xD(307)(4) <= CNStageIntLLROutputS5xD(230)(4);
  VNStageIntLLRInputS5xD(355)(4) <= CNStageIntLLROutputS5xD(230)(5);
  VNStageIntLLRInputS5xD(12)(4) <= CNStageIntLLROutputS5xD(231)(0);
  VNStageIntLLRInputS5xD(93)(4) <= CNStageIntLLROutputS5xD(231)(1);
  VNStageIntLLRInputS5xD(148)(4) <= CNStageIntLLROutputS5xD(231)(2);
  VNStageIntLLRInputS5xD(242)(4) <= CNStageIntLLROutputS5xD(231)(3);
  VNStageIntLLRInputS5xD(290)(4) <= CNStageIntLLROutputS5xD(231)(4);
  VNStageIntLLRInputS5xD(322)(3) <= CNStageIntLLROutputS5xD(231)(5);
  VNStageIntLLRInputS5xD(11)(4) <= CNStageIntLLROutputS5xD(232)(0);
  VNStageIntLLRInputS5xD(83)(4) <= CNStageIntLLROutputS5xD(232)(1);
  VNStageIntLLRInputS5xD(177)(4) <= CNStageIntLLROutputS5xD(232)(2);
  VNStageIntLLRInputS5xD(225)(4) <= CNStageIntLLROutputS5xD(232)(3);
  VNStageIntLLRInputS5xD(257)(4) <= CNStageIntLLROutputS5xD(232)(4);
  VNStageIntLLRInputS5xD(345)(3) <= CNStageIntLLROutputS5xD(232)(5);
  VNStageIntLLRInputS5xD(10)(3) <= CNStageIntLLROutputS5xD(233)(0);
  VNStageIntLLRInputS5xD(112)(4) <= CNStageIntLLROutputS5xD(233)(1);
  VNStageIntLLRInputS5xD(160)(4) <= CNStageIntLLROutputS5xD(233)(2);
  VNStageIntLLRInputS5xD(255)(4) <= CNStageIntLLROutputS5xD(233)(3);
  VNStageIntLLRInputS5xD(280)(4) <= CNStageIntLLROutputS5xD(233)(4);
  VNStageIntLLRInputS5xD(381)(3) <= CNStageIntLLROutputS5xD(233)(5);
  VNStageIntLLRInputS5xD(9)(4) <= CNStageIntLLROutputS5xD(234)(0);
  VNStageIntLLRInputS5xD(95)(4) <= CNStageIntLLROutputS5xD(234)(1);
  VNStageIntLLRInputS5xD(190)(2) <= CNStageIntLLROutputS5xD(234)(2);
  VNStageIntLLRInputS5xD(215)(4) <= CNStageIntLLROutputS5xD(234)(3);
  VNStageIntLLRInputS5xD(316)(2) <= CNStageIntLLROutputS5xD(234)(4);
  VNStageIntLLRInputS5xD(365)(4) <= CNStageIntLLROutputS5xD(234)(5);
  VNStageIntLLRInputS5xD(7)(4) <= CNStageIntLLROutputS5xD(235)(0);
  VNStageIntLLRInputS5xD(85)(3) <= CNStageIntLLROutputS5xD(235)(1);
  VNStageIntLLRInputS5xD(186)(3) <= CNStageIntLLROutputS5xD(235)(2);
  VNStageIntLLRInputS5xD(235)(3) <= CNStageIntLLROutputS5xD(235)(3);
  VNStageIntLLRInputS5xD(303)(4) <= CNStageIntLLROutputS5xD(235)(4);
  VNStageIntLLRInputS5xD(346)(4) <= CNStageIntLLROutputS5xD(235)(5);
  VNStageIntLLRInputS5xD(6)(4) <= CNStageIntLLROutputS5xD(236)(0);
  VNStageIntLLRInputS5xD(121)(3) <= CNStageIntLLROutputS5xD(236)(1);
  VNStageIntLLRInputS5xD(170)(3) <= CNStageIntLLROutputS5xD(236)(2);
  VNStageIntLLRInputS5xD(238)(4) <= CNStageIntLLROutputS5xD(236)(3);
  VNStageIntLLRInputS5xD(281)(4) <= CNStageIntLLROutputS5xD(236)(4);
  VNStageIntLLRInputS5xD(321)(4) <= CNStageIntLLROutputS5xD(236)(5);
  VNStageIntLLRInputS5xD(5)(4) <= CNStageIntLLROutputS5xD(237)(0);
  VNStageIntLLRInputS5xD(105)(3) <= CNStageIntLLROutputS5xD(237)(1);
  VNStageIntLLRInputS5xD(173)(4) <= CNStageIntLLROutputS5xD(237)(2);
  VNStageIntLLRInputS5xD(216)(4) <= CNStageIntLLROutputS5xD(237)(3);
  VNStageIntLLRInputS5xD(319)(4) <= CNStageIntLLROutputS5xD(237)(4);
  VNStageIntLLRInputS5xD(382)(3) <= CNStageIntLLROutputS5xD(237)(5);
  VNStageIntLLRInputS5xD(4)(3) <= CNStageIntLLROutputS5xD(238)(0);
  VNStageIntLLRInputS5xD(108)(4) <= CNStageIntLLROutputS5xD(238)(1);
  VNStageIntLLRInputS5xD(151)(4) <= CNStageIntLLROutputS5xD(238)(2);
  VNStageIntLLRInputS5xD(254)(2) <= CNStageIntLLROutputS5xD(238)(3);
  VNStageIntLLRInputS5xD(317)(1) <= CNStageIntLLROutputS5xD(238)(4);
  VNStageIntLLRInputS5xD(344)(4) <= CNStageIntLLROutputS5xD(238)(5);
  VNStageIntLLRInputS5xD(3)(3) <= CNStageIntLLROutputS5xD(239)(0);
  VNStageIntLLRInputS5xD(86)(2) <= CNStageIntLLROutputS5xD(239)(1);
  VNStageIntLLRInputS5xD(189)(3) <= CNStageIntLLROutputS5xD(239)(2);
  VNStageIntLLRInputS5xD(252)(3) <= CNStageIntLLROutputS5xD(239)(3);
  VNStageIntLLRInputS5xD(279)(4) <= CNStageIntLLROutputS5xD(239)(4);
  VNStageIntLLRInputS5xD(352)(4) <= CNStageIntLLROutputS5xD(239)(5);
  VNStageIntLLRInputS5xD(2)(4) <= CNStageIntLLROutputS5xD(240)(0);
  VNStageIntLLRInputS5xD(124)(2) <= CNStageIntLLROutputS5xD(240)(1);
  VNStageIntLLRInputS5xD(187)(3) <= CNStageIntLLROutputS5xD(240)(2);
  VNStageIntLLRInputS5xD(214)(4) <= CNStageIntLLROutputS5xD(240)(3);
  VNStageIntLLRInputS5xD(287)(4) <= CNStageIntLLROutputS5xD(240)(4);
  VNStageIntLLRInputS5xD(332)(4) <= CNStageIntLLROutputS5xD(240)(5);
  VNStageIntLLRInputS5xD(1)(3) <= CNStageIntLLROutputS5xD(241)(0);
  VNStageIntLLRInputS5xD(122)(3) <= CNStageIntLLROutputS5xD(241)(1);
  VNStageIntLLRInputS5xD(149)(4) <= CNStageIntLLROutputS5xD(241)(2);
  VNStageIntLLRInputS5xD(222)(2) <= CNStageIntLLROutputS5xD(241)(3);
  VNStageIntLLRInputS5xD(267)(4) <= CNStageIntLLROutputS5xD(241)(4);
  VNStageIntLLRInputS5xD(326)(3) <= CNStageIntLLROutputS5xD(241)(5);
  VNStageIntLLRInputS5xD(62)(3) <= CNStageIntLLROutputS5xD(242)(0);
  VNStageIntLLRInputS5xD(92)(4) <= CNStageIntLLROutputS5xD(242)(1);
  VNStageIntLLRInputS5xD(137)(4) <= CNStageIntLLROutputS5xD(242)(2);
  VNStageIntLLRInputS5xD(196)(4) <= CNStageIntLLROutputS5xD(242)(3);
  VNStageIntLLRInputS5xD(256)(3) <= CNStageIntLLROutputS5xD(242)(4);
  VNStageIntLLRInputS5xD(325)(4) <= CNStageIntLLROutputS5xD(242)(5);
  VNStageIntLLRInputS5xD(61)(3) <= CNStageIntLLROutputS5xD(243)(0);
  VNStageIntLLRInputS5xD(72)(4) <= CNStageIntLLROutputS5xD(243)(1);
  VNStageIntLLRInputS5xD(131)(3) <= CNStageIntLLROutputS5xD(243)(2);
  VNStageIntLLRInputS5xD(192)(4) <= CNStageIntLLROutputS5xD(243)(3);
  VNStageIntLLRInputS5xD(260)(4) <= CNStageIntLLROutputS5xD(243)(4);
  VNStageIntLLRInputS5xD(330)(4) <= CNStageIntLLROutputS5xD(243)(5);
  VNStageIntLLRInputS5xD(60)(3) <= CNStageIntLLROutputS5xD(244)(0);
  VNStageIntLLRInputS5xD(66)(3) <= CNStageIntLLROutputS5xD(244)(1);
  VNStageIntLLRInputS5xD(128)(4) <= CNStageIntLLROutputS5xD(244)(2);
  VNStageIntLLRInputS5xD(195)(3) <= CNStageIntLLROutputS5xD(244)(3);
  VNStageIntLLRInputS5xD(265)(3) <= CNStageIntLLROutputS5xD(244)(4);
  VNStageIntLLRInputS5xD(349)(3) <= CNStageIntLLROutputS5xD(244)(5);
  VNStageIntLLRInputS5xD(59)(2) <= CNStageIntLLROutputS5xD(245)(0);
  VNStageIntLLRInputS5xD(64)(3) <= CNStageIntLLROutputS5xD(245)(1);
  VNStageIntLLRInputS5xD(130)(4) <= CNStageIntLLROutputS5xD(245)(2);
  VNStageIntLLRInputS5xD(200)(4) <= CNStageIntLLROutputS5xD(245)(3);
  VNStageIntLLRInputS5xD(284)(4) <= CNStageIntLLROutputS5xD(245)(4);
  VNStageIntLLRInputS5xD(340)(4) <= CNStageIntLLROutputS5xD(245)(5);
  VNStageIntLLRInputS5xD(57)(3) <= CNStageIntLLROutputS5xD(246)(0);
  VNStageIntLLRInputS5xD(70)(4) <= CNStageIntLLROutputS5xD(246)(1);
  VNStageIntLLRInputS5xD(154)(3) <= CNStageIntLLROutputS5xD(246)(2);
  VNStageIntLLRInputS5xD(210)(4) <= CNStageIntLLROutputS5xD(246)(3);
  VNStageIntLLRInputS5xD(312)(3) <= CNStageIntLLROutputS5xD(246)(4);
  VNStageIntLLRInputS5xD(378)(3) <= CNStageIntLLROutputS5xD(246)(5);
  VNStageIntLLRInputS5xD(56)(4) <= CNStageIntLLROutputS5xD(247)(0);
  VNStageIntLLRInputS5xD(89)(4) <= CNStageIntLLROutputS5xD(247)(1);
  VNStageIntLLRInputS5xD(145)(4) <= CNStageIntLLROutputS5xD(247)(2);
  VNStageIntLLRInputS5xD(247)(4) <= CNStageIntLLROutputS5xD(247)(3);
  VNStageIntLLRInputS5xD(313)(2) <= CNStageIntLLROutputS5xD(247)(4);
  VNStageIntLLRInputS5xD(339)(4) <= CNStageIntLLROutputS5xD(247)(5);
  VNStageIntLLRInputS5xD(55)(4) <= CNStageIntLLROutputS5xD(248)(0);
  VNStageIntLLRInputS5xD(80)(4) <= CNStageIntLLROutputS5xD(248)(1);
  VNStageIntLLRInputS5xD(182)(4) <= CNStageIntLLROutputS5xD(248)(2);
  VNStageIntLLRInputS5xD(248)(4) <= CNStageIntLLROutputS5xD(248)(3);
  VNStageIntLLRInputS5xD(274)(3) <= CNStageIntLLROutputS5xD(248)(4);
  VNStageIntLLRInputS5xD(360)(4) <= CNStageIntLLROutputS5xD(248)(5);
  VNStageIntLLRInputS5xD(53)(3) <= CNStageIntLLROutputS5xD(249)(0);
  VNStageIntLLRInputS5xD(118)(3) <= CNStageIntLLROutputS5xD(249)(1);
  VNStageIntLLRInputS5xD(144)(4) <= CNStageIntLLROutputS5xD(249)(2);
  VNStageIntLLRInputS5xD(230)(3) <= CNStageIntLLROutputS5xD(249)(3);
  VNStageIntLLRInputS5xD(291)(4) <= CNStageIntLLROutputS5xD(249)(4);
  VNStageIntLLRInputS5xD(371)(3) <= CNStageIntLLROutputS5xD(249)(5);
  VNStageIntLLRInputS5xD(51)(3) <= CNStageIntLLROutputS5xD(250)(0);
  VNStageIntLLRInputS5xD(100)(4) <= CNStageIntLLROutputS5xD(250)(1);
  VNStageIntLLRInputS5xD(161)(4) <= CNStageIntLLROutputS5xD(250)(2);
  VNStageIntLLRInputS5xD(241)(3) <= CNStageIntLLROutputS5xD(250)(3);
  VNStageIntLLRInputS5xD(269)(3) <= CNStageIntLLROutputS5xD(250)(4);
  VNStageIntLLRInputS5xD(373)(2) <= CNStageIntLLROutputS5xD(250)(5);
  VNStageIntLLRInputS5xD(50)(4) <= CNStageIntLLROutputS5xD(251)(0);
  VNStageIntLLRInputS5xD(96)(4) <= CNStageIntLLROutputS5xD(251)(1);
  VNStageIntLLRInputS5xD(176)(4) <= CNStageIntLLROutputS5xD(251)(2);
  VNStageIntLLRInputS5xD(204)(4) <= CNStageIntLLROutputS5xD(251)(3);
  VNStageIntLLRInputS5xD(308)(2) <= CNStageIntLLROutputS5xD(251)(4);
  VNStageIntLLRInputS5xD(342)(3) <= CNStageIntLLROutputS5xD(251)(5);
  VNStageIntLLRInputS5xD(49)(4) <= CNStageIntLLROutputS5xD(252)(0);
  VNStageIntLLRInputS5xD(111)(4) <= CNStageIntLLROutputS5xD(252)(1);
  VNStageIntLLRInputS5xD(139)(4) <= CNStageIntLLROutputS5xD(252)(2);
  VNStageIntLLRInputS5xD(243)(4) <= CNStageIntLLROutputS5xD(252)(3);
  VNStageIntLLRInputS5xD(277)(4) <= CNStageIntLLROutputS5xD(252)(4);
  VNStageIntLLRInputS5xD(358)(3) <= CNStageIntLLROutputS5xD(252)(5);
  VNStageIntLLRInputS5xD(47)(2) <= CNStageIntLLROutputS5xD(253)(0);
  VNStageIntLLRInputS5xD(113)(4) <= CNStageIntLLROutputS5xD(253)(1);
  VNStageIntLLRInputS5xD(147)(4) <= CNStageIntLLROutputS5xD(253)(2);
  VNStageIntLLRInputS5xD(228)(4) <= CNStageIntLLROutputS5xD(253)(3);
  VNStageIntLLRInputS5xD(263)(4) <= CNStageIntLLROutputS5xD(253)(4);
  VNStageIntLLRInputS5xD(337)(4) <= CNStageIntLLROutputS5xD(253)(5);
  VNStageIntLLRInputS5xD(46)(4) <= CNStageIntLLROutputS5xD(254)(0);
  VNStageIntLLRInputS5xD(82)(4) <= CNStageIntLLROutputS5xD(254)(1);
  VNStageIntLLRInputS5xD(163)(3) <= CNStageIntLLROutputS5xD(254)(2);
  VNStageIntLLRInputS5xD(198)(4) <= CNStageIntLLROutputS5xD(254)(3);
  VNStageIntLLRInputS5xD(272)(4) <= CNStageIntLLROutputS5xD(254)(4);
  VNStageIntLLRInputS5xD(350)(4) <= CNStageIntLLROutputS5xD(254)(5);
  VNStageIntLLRInputS5xD(45)(4) <= CNStageIntLLROutputS5xD(255)(0);
  VNStageIntLLRInputS5xD(98)(3) <= CNStageIntLLROutputS5xD(255)(1);
  VNStageIntLLRInputS5xD(133)(2) <= CNStageIntLLROutputS5xD(255)(2);
  VNStageIntLLRInputS5xD(207)(3) <= CNStageIntLLROutputS5xD(255)(3);
  VNStageIntLLRInputS5xD(285)(4) <= CNStageIntLLROutputS5xD(255)(4);
  VNStageIntLLRInputS5xD(329)(4) <= CNStageIntLLROutputS5xD(255)(5);
  VNStageIntLLRInputS5xD(44)(4) <= CNStageIntLLROutputS5xD(256)(0);
  VNStageIntLLRInputS5xD(68)(3) <= CNStageIntLLROutputS5xD(256)(1);
  VNStageIntLLRInputS5xD(142)(3) <= CNStageIntLLROutputS5xD(256)(2);
  VNStageIntLLRInputS5xD(220)(4) <= CNStageIntLLROutputS5xD(256)(3);
  VNStageIntLLRInputS5xD(264)(4) <= CNStageIntLLROutputS5xD(256)(4);
  VNStageIntLLRInputS5xD(357)(4) <= CNStageIntLLROutputS5xD(256)(5);
  VNStageIntLLRInputS5xD(43)(3) <= CNStageIntLLROutputS5xD(257)(0);
  VNStageIntLLRInputS5xD(77)(2) <= CNStageIntLLROutputS5xD(257)(1);
  VNStageIntLLRInputS5xD(155)(4) <= CNStageIntLLROutputS5xD(257)(2);
  VNStageIntLLRInputS5xD(199)(4) <= CNStageIntLLROutputS5xD(257)(3);
  VNStageIntLLRInputS5xD(292)(4) <= CNStageIntLLROutputS5xD(257)(4);
  VNStageIntLLRInputS5xD(359)(4) <= CNStageIntLLROutputS5xD(257)(5);
  VNStageIntLLRInputS5xD(42)(4) <= CNStageIntLLROutputS5xD(258)(0);
  VNStageIntLLRInputS5xD(90)(4) <= CNStageIntLLROutputS5xD(258)(1);
  VNStageIntLLRInputS5xD(134)(3) <= CNStageIntLLROutputS5xD(258)(2);
  VNStageIntLLRInputS5xD(227)(4) <= CNStageIntLLROutputS5xD(258)(3);
  VNStageIntLLRInputS5xD(294)(4) <= CNStageIntLLROutputS5xD(258)(4);
  VNStageIntLLRInputS5xD(341)(4) <= CNStageIntLLROutputS5xD(258)(5);
  VNStageIntLLRInputS5xD(41)(4) <= CNStageIntLLROutputS5xD(259)(0);
  VNStageIntLLRInputS5xD(69)(4) <= CNStageIntLLROutputS5xD(259)(1);
  VNStageIntLLRInputS5xD(162)(4) <= CNStageIntLLROutputS5xD(259)(2);
  VNStageIntLLRInputS5xD(229)(3) <= CNStageIntLLROutputS5xD(259)(3);
  VNStageIntLLRInputS5xD(276)(4) <= CNStageIntLLROutputS5xD(259)(4);
  VNStageIntLLRInputS5xD(348)(4) <= CNStageIntLLROutputS5xD(259)(5);
  VNStageIntLLRInputS5xD(40)(3) <= CNStageIntLLROutputS5xD(260)(0);
  VNStageIntLLRInputS5xD(97)(4) <= CNStageIntLLROutputS5xD(260)(1);
  VNStageIntLLRInputS5xD(164)(4) <= CNStageIntLLROutputS5xD(260)(2);
  VNStageIntLLRInputS5xD(211)(4) <= CNStageIntLLROutputS5xD(260)(3);
  VNStageIntLLRInputS5xD(283)(4) <= CNStageIntLLROutputS5xD(260)(4);
  VNStageIntLLRInputS5xD(375)(3) <= CNStageIntLLROutputS5xD(260)(5);
  VNStageIntLLRInputS5xD(39)(4) <= CNStageIntLLROutputS5xD(261)(0);
  VNStageIntLLRInputS5xD(99)(4) <= CNStageIntLLROutputS5xD(261)(1);
  VNStageIntLLRInputS5xD(146)(3) <= CNStageIntLLROutputS5xD(261)(2);
  VNStageIntLLRInputS5xD(218)(4) <= CNStageIntLLROutputS5xD(261)(3);
  VNStageIntLLRInputS5xD(310)(3) <= CNStageIntLLROutputS5xD(261)(4);
  VNStageIntLLRInputS5xD(363)(3) <= CNStageIntLLROutputS5xD(261)(5);
  VNStageIntLLRInputS5xD(38)(4) <= CNStageIntLLROutputS5xD(262)(0);
  VNStageIntLLRInputS5xD(81)(3) <= CNStageIntLLROutputS5xD(262)(1);
  VNStageIntLLRInputS5xD(153)(4) <= CNStageIntLLROutputS5xD(262)(2);
  VNStageIntLLRInputS5xD(245)(4) <= CNStageIntLLROutputS5xD(262)(3);
  VNStageIntLLRInputS5xD(298)(4) <= CNStageIntLLROutputS5xD(262)(4);
  VNStageIntLLRInputS5xD(369)(3) <= CNStageIntLLROutputS5xD(262)(5);
  VNStageIntLLRInputS5xD(37)(4) <= CNStageIntLLROutputS5xD(263)(0);
  VNStageIntLLRInputS5xD(88)(4) <= CNStageIntLLROutputS5xD(263)(1);
  VNStageIntLLRInputS5xD(180)(2) <= CNStageIntLLROutputS5xD(263)(2);
  VNStageIntLLRInputS5xD(233)(3) <= CNStageIntLLROutputS5xD(263)(3);
  VNStageIntLLRInputS5xD(304)(4) <= CNStageIntLLROutputS5xD(263)(4);
  VNStageIntLLRInputS5xD(364)(4) <= CNStageIntLLROutputS5xD(263)(5);
  VNStageIntLLRInputS5xD(36)(3) <= CNStageIntLLROutputS5xD(264)(0);
  VNStageIntLLRInputS5xD(115)(4) <= CNStageIntLLROutputS5xD(264)(1);
  VNStageIntLLRInputS5xD(168)(3) <= CNStageIntLLROutputS5xD(264)(2);
  VNStageIntLLRInputS5xD(239)(4) <= CNStageIntLLROutputS5xD(264)(3);
  VNStageIntLLRInputS5xD(299)(3) <= CNStageIntLLROutputS5xD(264)(4);
  VNStageIntLLRInputS5xD(374)(4) <= CNStageIntLLROutputS5xD(264)(5);
  VNStageIntLLRInputS5xD(35)(4) <= CNStageIntLLROutputS5xD(265)(0);
  VNStageIntLLRInputS5xD(103)(4) <= CNStageIntLLROutputS5xD(265)(1);
  VNStageIntLLRInputS5xD(174)(3) <= CNStageIntLLROutputS5xD(265)(2);
  VNStageIntLLRInputS5xD(234)(4) <= CNStageIntLLROutputS5xD(265)(3);
  VNStageIntLLRInputS5xD(309)(4) <= CNStageIntLLROutputS5xD(265)(4);
  VNStageIntLLRInputS5xD(333)(3) <= CNStageIntLLROutputS5xD(265)(5);
  VNStageIntLLRInputS5xD(34)(4) <= CNStageIntLLROutputS5xD(266)(0);
  VNStageIntLLRInputS5xD(109)(4) <= CNStageIntLLROutputS5xD(266)(1);
  VNStageIntLLRInputS5xD(169)(4) <= CNStageIntLLROutputS5xD(266)(2);
  VNStageIntLLRInputS5xD(244)(1) <= CNStageIntLLROutputS5xD(266)(3);
  VNStageIntLLRInputS5xD(268)(4) <= CNStageIntLLROutputS5xD(266)(4);
  VNStageIntLLRInputS5xD(351)(3) <= CNStageIntLLROutputS5xD(266)(5);
  VNStageIntLLRInputS5xD(33)(4) <= CNStageIntLLROutputS5xD(267)(0);
  VNStageIntLLRInputS5xD(104)(4) <= CNStageIntLLROutputS5xD(267)(1);
  VNStageIntLLRInputS5xD(179)(4) <= CNStageIntLLROutputS5xD(267)(2);
  VNStageIntLLRInputS5xD(203)(4) <= CNStageIntLLROutputS5xD(267)(3);
  VNStageIntLLRInputS5xD(286)(4) <= CNStageIntLLROutputS5xD(267)(4);
  VNStageIntLLRInputS5xD(336)(3) <= CNStageIntLLROutputS5xD(267)(5);
  VNStageIntLLRInputS5xD(32)(3) <= CNStageIntLLROutputS5xD(268)(0);
  VNStageIntLLRInputS5xD(114)(4) <= CNStageIntLLROutputS5xD(268)(1);
  VNStageIntLLRInputS5xD(138)(4) <= CNStageIntLLROutputS5xD(268)(2);
  VNStageIntLLRInputS5xD(221)(4) <= CNStageIntLLROutputS5xD(268)(3);
  VNStageIntLLRInputS5xD(271)(3) <= CNStageIntLLROutputS5xD(268)(4);
  VNStageIntLLRInputS5xD(323)(3) <= CNStageIntLLROutputS5xD(268)(5);
  VNStageIntLLRInputS5xD(30)(4) <= CNStageIntLLROutputS5xD(269)(0);
  VNStageIntLLRInputS5xD(91)(4) <= CNStageIntLLROutputS5xD(269)(1);
  VNStageIntLLRInputS5xD(141)(2) <= CNStageIntLLROutputS5xD(269)(2);
  VNStageIntLLRInputS5xD(193)(3) <= CNStageIntLLROutputS5xD(269)(3);
  VNStageIntLLRInputS5xD(289)(4) <= CNStageIntLLROutputS5xD(269)(4);
  VNStageIntLLRInputS5xD(366)(4) <= CNStageIntLLROutputS5xD(269)(5);
  VNStageIntLLRInputS5xD(29)(3) <= CNStageIntLLROutputS5xD(270)(0);
  VNStageIntLLRInputS5xD(76)(4) <= CNStageIntLLROutputS5xD(270)(1);
  VNStageIntLLRInputS5xD(191)(4) <= CNStageIntLLROutputS5xD(270)(2);
  VNStageIntLLRInputS5xD(224)(4) <= CNStageIntLLROutputS5xD(270)(3);
  VNStageIntLLRInputS5xD(301)(4) <= CNStageIntLLROutputS5xD(270)(4);
  VNStageIntLLRInputS5xD(380)(3) <= CNStageIntLLROutputS5xD(270)(5);
  VNStageIntLLRInputS5xD(28)(4) <= CNStageIntLLROutputS5xD(271)(0);
  VNStageIntLLRInputS5xD(126)(3) <= CNStageIntLLROutputS5xD(271)(1);
  VNStageIntLLRInputS5xD(159)(3) <= CNStageIntLLROutputS5xD(271)(2);
  VNStageIntLLRInputS5xD(236)(4) <= CNStageIntLLROutputS5xD(271)(3);
  VNStageIntLLRInputS5xD(315)(3) <= CNStageIntLLROutputS5xD(271)(4);
  VNStageIntLLRInputS5xD(361)(4) <= CNStageIntLLROutputS5xD(271)(5);
  VNStageIntLLRInputS5xD(26)(4) <= CNStageIntLLROutputS5xD(272)(0);
  VNStageIntLLRInputS5xD(106)(3) <= CNStageIntLLROutputS5xD(272)(1);
  VNStageIntLLRInputS5xD(185)(1) <= CNStageIntLLROutputS5xD(272)(2);
  VNStageIntLLRInputS5xD(231)(3) <= CNStageIntLLROutputS5xD(272)(3);
  VNStageIntLLRInputS5xD(273)(3) <= CNStageIntLLROutputS5xD(272)(4);
  VNStageIntLLRInputS5xD(327)(4) <= CNStageIntLLROutputS5xD(272)(5);
  VNStageIntLLRInputS5xD(24)(4) <= CNStageIntLLROutputS5xD(273)(0);
  VNStageIntLLRInputS5xD(101)(4) <= CNStageIntLLROutputS5xD(273)(1);
  VNStageIntLLRInputS5xD(143)(4) <= CNStageIntLLROutputS5xD(273)(2);
  VNStageIntLLRInputS5xD(197)(4) <= CNStageIntLLROutputS5xD(273)(3);
  VNStageIntLLRInputS5xD(266)(3) <= CNStageIntLLROutputS5xD(273)(4);
  VNStageIntLLRInputS5xD(324)(4) <= CNStageIntLLROutputS5xD(273)(5);
  VNStageIntLLRInputS5xD(23)(4) <= CNStageIntLLROutputS5xD(274)(0);
  VNStageIntLLRInputS5xD(78)(4) <= CNStageIntLLROutputS5xD(274)(1);
  VNStageIntLLRInputS5xD(132)(3) <= CNStageIntLLROutputS5xD(274)(2);
  VNStageIntLLRInputS5xD(201)(4) <= CNStageIntLLROutputS5xD(274)(3);
  VNStageIntLLRInputS5xD(259)(2) <= CNStageIntLLROutputS5xD(274)(4);
  VNStageIntLLRInputS5xD(335)(4) <= CNStageIntLLROutputS5xD(274)(5);
  VNStageIntLLRInputS5xD(22)(4) <= CNStageIntLLROutputS5xD(275)(0);
  VNStageIntLLRInputS5xD(67)(1) <= CNStageIntLLROutputS5xD(275)(1);
  VNStageIntLLRInputS5xD(136)(4) <= CNStageIntLLROutputS5xD(275)(2);
  VNStageIntLLRInputS5xD(194)(4) <= CNStageIntLLROutputS5xD(275)(3);
  VNStageIntLLRInputS5xD(270)(4) <= CNStageIntLLROutputS5xD(275)(4);
  VNStageIntLLRInputS5xD(370)(3) <= CNStageIntLLROutputS5xD(275)(5);
  VNStageIntLLRInputS5xD(21)(4) <= CNStageIntLLROutputS5xD(276)(0);
  VNStageIntLLRInputS5xD(71)(3) <= CNStageIntLLROutputS5xD(276)(1);
  VNStageIntLLRInputS5xD(129)(4) <= CNStageIntLLROutputS5xD(276)(2);
  VNStageIntLLRInputS5xD(205)(1) <= CNStageIntLLROutputS5xD(276)(3);
  VNStageIntLLRInputS5xD(305)(4) <= CNStageIntLLROutputS5xD(276)(4);
  VNStageIntLLRInputS5xD(362)(4) <= CNStageIntLLROutputS5xD(276)(5);
  VNStageIntLLRInputS5xD(20)(2) <= CNStageIntLLROutputS5xD(277)(0);
  VNStageIntLLRInputS5xD(127)(4) <= CNStageIntLLROutputS5xD(277)(1);
  VNStageIntLLRInputS5xD(140)(4) <= CNStageIntLLROutputS5xD(277)(2);
  VNStageIntLLRInputS5xD(240)(4) <= CNStageIntLLROutputS5xD(277)(3);
  VNStageIntLLRInputS5xD(297)(4) <= CNStageIntLLROutputS5xD(277)(4);
  VNStageIntLLRInputS5xD(379)(2) <= CNStageIntLLROutputS5xD(277)(5);
  VNStageIntLLRInputS5xD(19)(3) <= CNStageIntLLROutputS5xD(278)(0);
  VNStageIntLLRInputS5xD(75)(4) <= CNStageIntLLROutputS5xD(278)(1);
  VNStageIntLLRInputS5xD(175)(4) <= CNStageIntLLROutputS5xD(278)(2);
  VNStageIntLLRInputS5xD(232)(3) <= CNStageIntLLROutputS5xD(278)(3);
  VNStageIntLLRInputS5xD(314)(1) <= CNStageIntLLROutputS5xD(278)(4);
  VNStageIntLLRInputS5xD(376)(3) <= CNStageIntLLROutputS5xD(278)(5);
  VNStageIntLLRInputS5xD(0)(4) <= CNStageIntLLROutputS5xD(279)(0);
  VNStageIntLLRInputS5xD(123)(3) <= CNStageIntLLROutputS5xD(279)(1);
  VNStageIntLLRInputS5xD(188)(2) <= CNStageIntLLROutputS5xD(279)(2);
  VNStageIntLLRInputS5xD(253)(3) <= CNStageIntLLROutputS5xD(279)(3);
  VNStageIntLLRInputS5xD(318)(2) <= CNStageIntLLROutputS5xD(279)(4);
  VNStageIntLLRInputS5xD(383)(4) <= CNStageIntLLROutputS5xD(279)(5);
  VNStageIntLLRInputS5xD(35)(5) <= CNStageIntLLROutputS5xD(280)(0);
  VNStageIntLLRInputS5xD(91)(5) <= CNStageIntLLROutputS5xD(280)(1);
  VNStageIntLLRInputS5xD(191)(5) <= CNStageIntLLROutputS5xD(280)(2);
  VNStageIntLLRInputS5xD(248)(5) <= CNStageIntLLROutputS5xD(280)(3);
  VNStageIntLLRInputS5xD(267)(5) <= CNStageIntLLROutputS5xD(280)(4);
  VNStageIntLLRInputS5xD(329)(5) <= CNStageIntLLROutputS5xD(280)(5);
  VNStageIntLLRInputS5xD(34)(5) <= CNStageIntLLROutputS5xD(281)(0);
  VNStageIntLLRInputS5xD(126)(4) <= CNStageIntLLROutputS5xD(281)(1);
  VNStageIntLLRInputS5xD(183)(3) <= CNStageIntLLROutputS5xD(281)(2);
  VNStageIntLLRInputS5xD(202)(4) <= CNStageIntLLROutputS5xD(281)(3);
  VNStageIntLLRInputS5xD(264)(5) <= CNStageIntLLROutputS5xD(281)(4);
  VNStageIntLLRInputS5xD(363)(4) <= CNStageIntLLROutputS5xD(281)(5);
  VNStageIntLLRInputS5xD(33)(5) <= CNStageIntLLROutputS5xD(282)(0);
  VNStageIntLLRInputS5xD(118)(4) <= CNStageIntLLROutputS5xD(282)(1);
  VNStageIntLLRInputS5xD(137)(5) <= CNStageIntLLROutputS5xD(282)(2);
  VNStageIntLLRInputS5xD(199)(5) <= CNStageIntLLROutputS5xD(282)(3);
  VNStageIntLLRInputS5xD(298)(5) <= CNStageIntLLROutputS5xD(282)(4);
  VNStageIntLLRInputS5xD(383)(5) <= CNStageIntLLROutputS5xD(282)(5);
  VNStageIntLLRInputS5xD(31)(3) <= CNStageIntLLROutputS5xD(283)(0);
  VNStageIntLLRInputS5xD(69)(5) <= CNStageIntLLROutputS5xD(283)(1);
  VNStageIntLLRInputS5xD(168)(4) <= CNStageIntLLROutputS5xD(283)(2);
  VNStageIntLLRInputS5xD(253)(4) <= CNStageIntLLROutputS5xD(283)(3);
  VNStageIntLLRInputS5xD(304)(5) <= CNStageIntLLROutputS5xD(283)(4);
  VNStageIntLLRInputS5xD(359)(5) <= CNStageIntLLROutputS5xD(283)(5);
  VNStageIntLLRInputS5xD(30)(5) <= CNStageIntLLROutputS5xD(284)(0);
  VNStageIntLLRInputS5xD(103)(5) <= CNStageIntLLROutputS5xD(284)(1);
  VNStageIntLLRInputS5xD(188)(3) <= CNStageIntLLROutputS5xD(284)(2);
  VNStageIntLLRInputS5xD(239)(5) <= CNStageIntLLROutputS5xD(284)(3);
  VNStageIntLLRInputS5xD(294)(5) <= CNStageIntLLROutputS5xD(284)(4);
  VNStageIntLLRInputS5xD(325)(5) <= CNStageIntLLROutputS5xD(284)(5);
  VNStageIntLLRInputS5xD(27)(4) <= CNStageIntLLROutputS5xD(285)(0);
  VNStageIntLLRInputS5xD(99)(5) <= CNStageIntLLROutputS5xD(285)(1);
  VNStageIntLLRInputS5xD(130)(5) <= CNStageIntLLROutputS5xD(285)(2);
  VNStageIntLLRInputS5xD(241)(4) <= CNStageIntLLROutputS5xD(285)(3);
  VNStageIntLLRInputS5xD(273)(4) <= CNStageIntLLROutputS5xD(285)(4);
  VNStageIntLLRInputS5xD(361)(5) <= CNStageIntLLROutputS5xD(285)(5);
  VNStageIntLLRInputS5xD(26)(5) <= CNStageIntLLROutputS5xD(286)(0);
  VNStageIntLLRInputS5xD(65)(4) <= CNStageIntLLROutputS5xD(286)(1);
  VNStageIntLLRInputS5xD(176)(5) <= CNStageIntLLROutputS5xD(286)(2);
  VNStageIntLLRInputS5xD(208)(4) <= CNStageIntLLROutputS5xD(286)(3);
  VNStageIntLLRInputS5xD(296)(4) <= CNStageIntLLROutputS5xD(286)(4);
  VNStageIntLLRInputS5xD(334)(3) <= CNStageIntLLROutputS5xD(286)(5);
  VNStageIntLLRInputS5xD(25)(4) <= CNStageIntLLROutputS5xD(287)(0);
  VNStageIntLLRInputS5xD(111)(5) <= CNStageIntLLROutputS5xD(287)(1);
  VNStageIntLLRInputS5xD(143)(5) <= CNStageIntLLROutputS5xD(287)(2);
  VNStageIntLLRInputS5xD(231)(4) <= CNStageIntLLROutputS5xD(287)(3);
  VNStageIntLLRInputS5xD(269)(4) <= CNStageIntLLROutputS5xD(287)(4);
  VNStageIntLLRInputS5xD(381)(4) <= CNStageIntLLROutputS5xD(287)(5);
  VNStageIntLLRInputS5xD(24)(5) <= CNStageIntLLROutputS5xD(288)(0);
  VNStageIntLLRInputS5xD(78)(5) <= CNStageIntLLROutputS5xD(288)(1);
  VNStageIntLLRInputS5xD(166)(4) <= CNStageIntLLROutputS5xD(288)(2);
  VNStageIntLLRInputS5xD(204)(5) <= CNStageIntLLROutputS5xD(288)(3);
  VNStageIntLLRInputS5xD(316)(3) <= CNStageIntLLROutputS5xD(288)(4);
  VNStageIntLLRInputS5xD(321)(5) <= CNStageIntLLROutputS5xD(288)(5);
  VNStageIntLLRInputS5xD(23)(5) <= CNStageIntLLROutputS5xD(289)(0);
  VNStageIntLLRInputS5xD(101)(5) <= CNStageIntLLROutputS5xD(289)(1);
  VNStageIntLLRInputS5xD(139)(5) <= CNStageIntLLROutputS5xD(289)(2);
  VNStageIntLLRInputS5xD(251)(3) <= CNStageIntLLROutputS5xD(289)(3);
  VNStageIntLLRInputS5xD(319)(5) <= CNStageIntLLROutputS5xD(289)(4);
  VNStageIntLLRInputS5xD(362)(5) <= CNStageIntLLROutputS5xD(289)(5);
  VNStageIntLLRInputS5xD(22)(5) <= CNStageIntLLROutputS5xD(290)(0);
  VNStageIntLLRInputS5xD(74)(4) <= CNStageIntLLROutputS5xD(290)(1);
  VNStageIntLLRInputS5xD(186)(4) <= CNStageIntLLROutputS5xD(290)(2);
  VNStageIntLLRInputS5xD(254)(3) <= CNStageIntLLROutputS5xD(290)(3);
  VNStageIntLLRInputS5xD(297)(5) <= CNStageIntLLROutputS5xD(290)(4);
  VNStageIntLLRInputS5xD(337)(5) <= CNStageIntLLROutputS5xD(290)(5);
  VNStageIntLLRInputS5xD(21)(5) <= CNStageIntLLROutputS5xD(291)(0);
  VNStageIntLLRInputS5xD(121)(4) <= CNStageIntLLROutputS5xD(291)(1);
  VNStageIntLLRInputS5xD(189)(4) <= CNStageIntLLROutputS5xD(291)(2);
  VNStageIntLLRInputS5xD(232)(4) <= CNStageIntLLROutputS5xD(291)(3);
  VNStageIntLLRInputS5xD(272)(5) <= CNStageIntLLROutputS5xD(291)(4);
  VNStageIntLLRInputS5xD(335)(5) <= CNStageIntLLROutputS5xD(291)(5);
  VNStageIntLLRInputS5xD(20)(3) <= CNStageIntLLROutputS5xD(292)(0);
  VNStageIntLLRInputS5xD(124)(3) <= CNStageIntLLROutputS5xD(292)(1);
  VNStageIntLLRInputS5xD(167)(5) <= CNStageIntLLROutputS5xD(292)(2);
  VNStageIntLLRInputS5xD(207)(4) <= CNStageIntLLROutputS5xD(292)(3);
  VNStageIntLLRInputS5xD(270)(5) <= CNStageIntLLROutputS5xD(292)(4);
  VNStageIntLLRInputS5xD(360)(5) <= CNStageIntLLROutputS5xD(292)(5);
  VNStageIntLLRInputS5xD(18)(5) <= CNStageIntLLROutputS5xD(293)(0);
  VNStageIntLLRInputS5xD(77)(3) <= CNStageIntLLROutputS5xD(293)(1);
  VNStageIntLLRInputS5xD(140)(5) <= CNStageIntLLROutputS5xD(293)(2);
  VNStageIntLLRInputS5xD(230)(4) <= CNStageIntLLROutputS5xD(293)(3);
  VNStageIntLLRInputS5xD(303)(5) <= CNStageIntLLROutputS5xD(293)(4);
  VNStageIntLLRInputS5xD(348)(5) <= CNStageIntLLROutputS5xD(293)(5);
  VNStageIntLLRInputS5xD(17)(5) <= CNStageIntLLROutputS5xD(294)(0);
  VNStageIntLLRInputS5xD(75)(5) <= CNStageIntLLROutputS5xD(294)(1);
  VNStageIntLLRInputS5xD(165)(4) <= CNStageIntLLROutputS5xD(294)(2);
  VNStageIntLLRInputS5xD(238)(5) <= CNStageIntLLROutputS5xD(294)(3);
  VNStageIntLLRInputS5xD(283)(5) <= CNStageIntLLROutputS5xD(294)(4);
  VNStageIntLLRInputS5xD(342)(4) <= CNStageIntLLROutputS5xD(294)(5);
  VNStageIntLLRInputS5xD(16)(4) <= CNStageIntLLROutputS5xD(295)(0);
  VNStageIntLLRInputS5xD(100)(5) <= CNStageIntLLROutputS5xD(295)(1);
  VNStageIntLLRInputS5xD(173)(5) <= CNStageIntLLROutputS5xD(295)(2);
  VNStageIntLLRInputS5xD(218)(5) <= CNStageIntLLROutputS5xD(295)(3);
  VNStageIntLLRInputS5xD(277)(5) <= CNStageIntLLROutputS5xD(295)(4);
  VNStageIntLLRInputS5xD(320)(3) <= CNStageIntLLROutputS5xD(295)(5);
  VNStageIntLLRInputS5xD(15)(5) <= CNStageIntLLROutputS5xD(296)(0);
  VNStageIntLLRInputS5xD(108)(5) <= CNStageIntLLROutputS5xD(296)(1);
  VNStageIntLLRInputS5xD(153)(5) <= CNStageIntLLROutputS5xD(296)(2);
  VNStageIntLLRInputS5xD(212)(4) <= CNStageIntLLROutputS5xD(296)(3);
  VNStageIntLLRInputS5xD(256)(4) <= CNStageIntLLROutputS5xD(296)(4);
  VNStageIntLLRInputS5xD(341)(5) <= CNStageIntLLROutputS5xD(296)(5);
  VNStageIntLLRInputS5xD(14)(5) <= CNStageIntLLROutputS5xD(297)(0);
  VNStageIntLLRInputS5xD(88)(5) <= CNStageIntLLROutputS5xD(297)(1);
  VNStageIntLLRInputS5xD(147)(5) <= CNStageIntLLROutputS5xD(297)(2);
  VNStageIntLLRInputS5xD(192)(5) <= CNStageIntLLROutputS5xD(297)(3);
  VNStageIntLLRInputS5xD(276)(5) <= CNStageIntLLROutputS5xD(297)(4);
  VNStageIntLLRInputS5xD(346)(5) <= CNStageIntLLROutputS5xD(297)(5);
  VNStageIntLLRInputS5xD(13)(4) <= CNStageIntLLROutputS5xD(298)(0);
  VNStageIntLLRInputS5xD(82)(5) <= CNStageIntLLROutputS5xD(298)(1);
  VNStageIntLLRInputS5xD(128)(5) <= CNStageIntLLROutputS5xD(298)(2);
  VNStageIntLLRInputS5xD(211)(5) <= CNStageIntLLROutputS5xD(298)(3);
  VNStageIntLLRInputS5xD(281)(5) <= CNStageIntLLROutputS5xD(298)(4);
  VNStageIntLLRInputS5xD(365)(5) <= CNStageIntLLROutputS5xD(298)(5);
  VNStageIntLLRInputS5xD(12)(5) <= CNStageIntLLROutputS5xD(299)(0);
  VNStageIntLLRInputS5xD(64)(4) <= CNStageIntLLROutputS5xD(299)(1);
  VNStageIntLLRInputS5xD(146)(4) <= CNStageIntLLROutputS5xD(299)(2);
  VNStageIntLLRInputS5xD(216)(5) <= CNStageIntLLROutputS5xD(299)(3);
  VNStageIntLLRInputS5xD(300)(4) <= CNStageIntLLROutputS5xD(299)(4);
  VNStageIntLLRInputS5xD(356)(4) <= CNStageIntLLROutputS5xD(299)(5);
  VNStageIntLLRInputS5xD(9)(5) <= CNStageIntLLROutputS5xD(300)(0);
  VNStageIntLLRInputS5xD(105)(4) <= CNStageIntLLROutputS5xD(300)(1);
  VNStageIntLLRInputS5xD(161)(5) <= CNStageIntLLROutputS5xD(300)(2);
  VNStageIntLLRInputS5xD(200)(5) <= CNStageIntLLROutputS5xD(300)(3);
  VNStageIntLLRInputS5xD(266)(4) <= CNStageIntLLROutputS5xD(300)(4);
  VNStageIntLLRInputS5xD(355)(5) <= CNStageIntLLROutputS5xD(300)(5);
  VNStageIntLLRInputS5xD(7)(5) <= CNStageIntLLROutputS5xD(301)(0);
  VNStageIntLLRInputS5xD(70)(5) <= CNStageIntLLROutputS5xD(301)(1);
  VNStageIntLLRInputS5xD(136)(5) <= CNStageIntLLROutputS5xD(301)(2);
  VNStageIntLLRInputS5xD(225)(5) <= CNStageIntLLROutputS5xD(301)(3);
  VNStageIntLLRInputS5xD(311)(4) <= CNStageIntLLROutputS5xD(301)(4);
  VNStageIntLLRInputS5xD(372)(4) <= CNStageIntLLROutputS5xD(301)(5);
  VNStageIntLLRInputS5xD(6)(5) <= CNStageIntLLROutputS5xD(302)(0);
  VNStageIntLLRInputS5xD(71)(4) <= CNStageIntLLROutputS5xD(302)(1);
  VNStageIntLLRInputS5xD(160)(5) <= CNStageIntLLROutputS5xD(302)(2);
  VNStageIntLLRInputS5xD(246)(5) <= CNStageIntLLROutputS5xD(302)(3);
  VNStageIntLLRInputS5xD(307)(5) <= CNStageIntLLROutputS5xD(302)(4);
  VNStageIntLLRInputS5xD(324)(5) <= CNStageIntLLROutputS5xD(302)(5);
  VNStageIntLLRInputS5xD(5)(5) <= CNStageIntLLROutputS5xD(303)(0);
  VNStageIntLLRInputS5xD(95)(5) <= CNStageIntLLROutputS5xD(303)(1);
  VNStageIntLLRInputS5xD(181)(5) <= CNStageIntLLROutputS5xD(303)(2);
  VNStageIntLLRInputS5xD(242)(5) <= CNStageIntLLROutputS5xD(303)(3);
  VNStageIntLLRInputS5xD(259)(3) <= CNStageIntLLROutputS5xD(303)(4);
  VNStageIntLLRInputS5xD(350)(5) <= CNStageIntLLROutputS5xD(303)(5);
  VNStageIntLLRInputS5xD(4)(4) <= CNStageIntLLROutputS5xD(304)(0);
  VNStageIntLLRInputS5xD(116)(4) <= CNStageIntLLROutputS5xD(304)(1);
  VNStageIntLLRInputS5xD(177)(5) <= CNStageIntLLROutputS5xD(304)(2);
  VNStageIntLLRInputS5xD(194)(5) <= CNStageIntLLROutputS5xD(304)(3);
  VNStageIntLLRInputS5xD(285)(5) <= CNStageIntLLROutputS5xD(304)(4);
  VNStageIntLLRInputS5xD(326)(4) <= CNStageIntLLROutputS5xD(304)(5);
  VNStageIntLLRInputS5xD(3)(4) <= CNStageIntLLROutputS5xD(305)(0);
  VNStageIntLLRInputS5xD(112)(5) <= CNStageIntLLROutputS5xD(305)(1);
  VNStageIntLLRInputS5xD(129)(5) <= CNStageIntLLROutputS5xD(305)(2);
  VNStageIntLLRInputS5xD(220)(5) <= CNStageIntLLROutputS5xD(305)(3);
  VNStageIntLLRInputS5xD(261)(4) <= CNStageIntLLROutputS5xD(305)(4);
  VNStageIntLLRInputS5xD(358)(4) <= CNStageIntLLROutputS5xD(305)(5);
  VNStageIntLLRInputS5xD(2)(5) <= CNStageIntLLROutputS5xD(306)(0);
  VNStageIntLLRInputS5xD(127)(5) <= CNStageIntLLROutputS5xD(306)(1);
  VNStageIntLLRInputS5xD(155)(5) <= CNStageIntLLROutputS5xD(306)(2);
  VNStageIntLLRInputS5xD(196)(5) <= CNStageIntLLROutputS5xD(306)(3);
  VNStageIntLLRInputS5xD(293)(4) <= CNStageIntLLROutputS5xD(306)(4);
  VNStageIntLLRInputS5xD(374)(5) <= CNStageIntLLROutputS5xD(306)(5);
  VNStageIntLLRInputS5xD(1)(4) <= CNStageIntLLROutputS5xD(307)(0);
  VNStageIntLLRInputS5xD(90)(5) <= CNStageIntLLROutputS5xD(307)(1);
  VNStageIntLLRInputS5xD(131)(4) <= CNStageIntLLROutputS5xD(307)(2);
  VNStageIntLLRInputS5xD(228)(5) <= CNStageIntLLROutputS5xD(307)(3);
  VNStageIntLLRInputS5xD(309)(5) <= CNStageIntLLROutputS5xD(307)(4);
  VNStageIntLLRInputS5xD(344)(5) <= CNStageIntLLROutputS5xD(307)(5);
  VNStageIntLLRInputS5xD(62)(4) <= CNStageIntLLROutputS5xD(308)(0);
  VNStageIntLLRInputS5xD(98)(4) <= CNStageIntLLROutputS5xD(308)(1);
  VNStageIntLLRInputS5xD(179)(5) <= CNStageIntLLROutputS5xD(308)(2);
  VNStageIntLLRInputS5xD(214)(5) <= CNStageIntLLROutputS5xD(308)(3);
  VNStageIntLLRInputS5xD(288)(5) <= CNStageIntLLROutputS5xD(308)(4);
  VNStageIntLLRInputS5xD(366)(5) <= CNStageIntLLROutputS5xD(308)(5);
  VNStageIntLLRInputS5xD(61)(4) <= CNStageIntLLROutputS5xD(309)(0);
  VNStageIntLLRInputS5xD(114)(5) <= CNStageIntLLROutputS5xD(309)(1);
  VNStageIntLLRInputS5xD(149)(5) <= CNStageIntLLROutputS5xD(309)(2);
  VNStageIntLLRInputS5xD(223)(5) <= CNStageIntLLROutputS5xD(309)(3);
  VNStageIntLLRInputS5xD(301)(5) <= CNStageIntLLROutputS5xD(309)(4);
  VNStageIntLLRInputS5xD(345)(4) <= CNStageIntLLROutputS5xD(309)(5);
  VNStageIntLLRInputS5xD(60)(4) <= CNStageIntLLROutputS5xD(310)(0);
  VNStageIntLLRInputS5xD(84)(4) <= CNStageIntLLROutputS5xD(310)(1);
  VNStageIntLLRInputS5xD(158)(5) <= CNStageIntLLROutputS5xD(310)(2);
  VNStageIntLLRInputS5xD(236)(5) <= CNStageIntLLROutputS5xD(310)(3);
  VNStageIntLLRInputS5xD(280)(5) <= CNStageIntLLROutputS5xD(310)(4);
  VNStageIntLLRInputS5xD(373)(3) <= CNStageIntLLROutputS5xD(310)(5);
  VNStageIntLLRInputS5xD(59)(3) <= CNStageIntLLROutputS5xD(311)(0);
  VNStageIntLLRInputS5xD(93)(5) <= CNStageIntLLROutputS5xD(311)(1);
  VNStageIntLLRInputS5xD(171)(3) <= CNStageIntLLROutputS5xD(311)(2);
  VNStageIntLLRInputS5xD(215)(5) <= CNStageIntLLROutputS5xD(311)(3);
  VNStageIntLLRInputS5xD(308)(3) <= CNStageIntLLROutputS5xD(311)(4);
  VNStageIntLLRInputS5xD(375)(4) <= CNStageIntLLROutputS5xD(311)(5);
  VNStageIntLLRInputS5xD(58)(3) <= CNStageIntLLROutputS5xD(312)(0);
  VNStageIntLLRInputS5xD(106)(4) <= CNStageIntLLROutputS5xD(312)(1);
  VNStageIntLLRInputS5xD(150)(4) <= CNStageIntLLROutputS5xD(312)(2);
  VNStageIntLLRInputS5xD(243)(5) <= CNStageIntLLROutputS5xD(312)(3);
  VNStageIntLLRInputS5xD(310)(4) <= CNStageIntLLROutputS5xD(312)(4);
  VNStageIntLLRInputS5xD(357)(5) <= CNStageIntLLROutputS5xD(312)(5);
  VNStageIntLLRInputS5xD(57)(4) <= CNStageIntLLROutputS5xD(313)(0);
  VNStageIntLLRInputS5xD(85)(4) <= CNStageIntLLROutputS5xD(313)(1);
  VNStageIntLLRInputS5xD(178)(4) <= CNStageIntLLROutputS5xD(313)(2);
  VNStageIntLLRInputS5xD(245)(5) <= CNStageIntLLROutputS5xD(313)(3);
  VNStageIntLLRInputS5xD(292)(5) <= CNStageIntLLROutputS5xD(313)(4);
  VNStageIntLLRInputS5xD(364)(5) <= CNStageIntLLROutputS5xD(313)(5);
  VNStageIntLLRInputS5xD(56)(5) <= CNStageIntLLROutputS5xD(314)(0);
  VNStageIntLLRInputS5xD(113)(5) <= CNStageIntLLROutputS5xD(314)(1);
  VNStageIntLLRInputS5xD(180)(3) <= CNStageIntLLROutputS5xD(314)(2);
  VNStageIntLLRInputS5xD(227)(5) <= CNStageIntLLROutputS5xD(314)(3);
  VNStageIntLLRInputS5xD(299)(4) <= CNStageIntLLROutputS5xD(314)(4);
  VNStageIntLLRInputS5xD(328)(3) <= CNStageIntLLROutputS5xD(314)(5);
  VNStageIntLLRInputS5xD(55)(5) <= CNStageIntLLROutputS5xD(315)(0);
  VNStageIntLLRInputS5xD(115)(5) <= CNStageIntLLROutputS5xD(315)(1);
  VNStageIntLLRInputS5xD(162)(5) <= CNStageIntLLROutputS5xD(315)(2);
  VNStageIntLLRInputS5xD(234)(5) <= CNStageIntLLROutputS5xD(315)(3);
  VNStageIntLLRInputS5xD(263)(5) <= CNStageIntLLROutputS5xD(315)(4);
  VNStageIntLLRInputS5xD(379)(3) <= CNStageIntLLROutputS5xD(315)(5);
  VNStageIntLLRInputS5xD(54)(4) <= CNStageIntLLROutputS5xD(316)(0);
  VNStageIntLLRInputS5xD(97)(5) <= CNStageIntLLROutputS5xD(316)(1);
  VNStageIntLLRInputS5xD(169)(5) <= CNStageIntLLROutputS5xD(316)(2);
  VNStageIntLLRInputS5xD(198)(5) <= CNStageIntLLROutputS5xD(316)(3);
  VNStageIntLLRInputS5xD(314)(2) <= CNStageIntLLROutputS5xD(316)(4);
  VNStageIntLLRInputS5xD(322)(4) <= CNStageIntLLROutputS5xD(316)(5);
  VNStageIntLLRInputS5xD(53)(4) <= CNStageIntLLROutputS5xD(317)(0);
  VNStageIntLLRInputS5xD(104)(5) <= CNStageIntLLROutputS5xD(317)(1);
  VNStageIntLLRInputS5xD(133)(3) <= CNStageIntLLROutputS5xD(317)(2);
  VNStageIntLLRInputS5xD(249)(3) <= CNStageIntLLROutputS5xD(317)(3);
  VNStageIntLLRInputS5xD(257)(5) <= CNStageIntLLROutputS5xD(317)(4);
  VNStageIntLLRInputS5xD(380)(4) <= CNStageIntLLROutputS5xD(317)(5);
  VNStageIntLLRInputS5xD(52)(3) <= CNStageIntLLROutputS5xD(318)(0);
  VNStageIntLLRInputS5xD(68)(4) <= CNStageIntLLROutputS5xD(318)(1);
  VNStageIntLLRInputS5xD(184)(5) <= CNStageIntLLROutputS5xD(318)(2);
  VNStageIntLLRInputS5xD(255)(5) <= CNStageIntLLROutputS5xD(318)(3);
  VNStageIntLLRInputS5xD(315)(4) <= CNStageIntLLROutputS5xD(318)(4);
  VNStageIntLLRInputS5xD(327)(5) <= CNStageIntLLROutputS5xD(318)(5);
  VNStageIntLLRInputS5xD(51)(4) <= CNStageIntLLROutputS5xD(319)(0);
  VNStageIntLLRInputS5xD(119)(4) <= CNStageIntLLROutputS5xD(319)(1);
  VNStageIntLLRInputS5xD(190)(3) <= CNStageIntLLROutputS5xD(319)(2);
  VNStageIntLLRInputS5xD(250)(3) <= CNStageIntLLROutputS5xD(319)(3);
  VNStageIntLLRInputS5xD(262)(4) <= CNStageIntLLROutputS5xD(319)(4);
  VNStageIntLLRInputS5xD(349)(4) <= CNStageIntLLROutputS5xD(319)(5);
  VNStageIntLLRInputS5xD(50)(5) <= CNStageIntLLROutputS5xD(320)(0);
  VNStageIntLLRInputS5xD(125)(2) <= CNStageIntLLROutputS5xD(320)(1);
  VNStageIntLLRInputS5xD(185)(2) <= CNStageIntLLROutputS5xD(320)(2);
  VNStageIntLLRInputS5xD(197)(5) <= CNStageIntLLROutputS5xD(320)(3);
  VNStageIntLLRInputS5xD(284)(5) <= CNStageIntLLROutputS5xD(320)(4);
  VNStageIntLLRInputS5xD(367)(5) <= CNStageIntLLROutputS5xD(320)(5);
  VNStageIntLLRInputS5xD(49)(5) <= CNStageIntLLROutputS5xD(321)(0);
  VNStageIntLLRInputS5xD(120)(2) <= CNStageIntLLROutputS5xD(321)(1);
  VNStageIntLLRInputS5xD(132)(4) <= CNStageIntLLROutputS5xD(321)(2);
  VNStageIntLLRInputS5xD(219)(4) <= CNStageIntLLROutputS5xD(321)(3);
  VNStageIntLLRInputS5xD(302)(5) <= CNStageIntLLROutputS5xD(321)(4);
  VNStageIntLLRInputS5xD(352)(5) <= CNStageIntLLROutputS5xD(321)(5);
  VNStageIntLLRInputS5xD(48)(2) <= CNStageIntLLROutputS5xD(322)(0);
  VNStageIntLLRInputS5xD(67)(2) <= CNStageIntLLROutputS5xD(322)(1);
  VNStageIntLLRInputS5xD(154)(4) <= CNStageIntLLROutputS5xD(322)(2);
  VNStageIntLLRInputS5xD(237)(4) <= CNStageIntLLROutputS5xD(322)(3);
  VNStageIntLLRInputS5xD(287)(5) <= CNStageIntLLROutputS5xD(322)(4);
  VNStageIntLLRInputS5xD(339)(5) <= CNStageIntLLROutputS5xD(322)(5);
  VNStageIntLLRInputS5xD(46)(5) <= CNStageIntLLROutputS5xD(323)(0);
  VNStageIntLLRInputS5xD(107)(4) <= CNStageIntLLROutputS5xD(323)(1);
  VNStageIntLLRInputS5xD(157)(4) <= CNStageIntLLROutputS5xD(323)(2);
  VNStageIntLLRInputS5xD(209)(4) <= CNStageIntLLROutputS5xD(323)(3);
  VNStageIntLLRInputS5xD(305)(5) <= CNStageIntLLROutputS5xD(323)(4);
  VNStageIntLLRInputS5xD(382)(4) <= CNStageIntLLROutputS5xD(323)(5);
  VNStageIntLLRInputS5xD(45)(5) <= CNStageIntLLROutputS5xD(324)(0);
  VNStageIntLLRInputS5xD(92)(5) <= CNStageIntLLROutputS5xD(324)(1);
  VNStageIntLLRInputS5xD(144)(5) <= CNStageIntLLROutputS5xD(324)(2);
  VNStageIntLLRInputS5xD(240)(5) <= CNStageIntLLROutputS5xD(324)(3);
  VNStageIntLLRInputS5xD(317)(2) <= CNStageIntLLROutputS5xD(324)(4);
  VNStageIntLLRInputS5xD(333)(4) <= CNStageIntLLROutputS5xD(324)(5);
  VNStageIntLLRInputS5xD(44)(5) <= CNStageIntLLROutputS5xD(325)(0);
  VNStageIntLLRInputS5xD(79)(4) <= CNStageIntLLROutputS5xD(325)(1);
  VNStageIntLLRInputS5xD(175)(5) <= CNStageIntLLROutputS5xD(325)(2);
  VNStageIntLLRInputS5xD(252)(4) <= CNStageIntLLROutputS5xD(325)(3);
  VNStageIntLLRInputS5xD(268)(5) <= CNStageIntLLROutputS5xD(325)(4);
  VNStageIntLLRInputS5xD(377)(3) <= CNStageIntLLROutputS5xD(325)(5);
  VNStageIntLLRInputS5xD(43)(4) <= CNStageIntLLROutputS5xD(326)(0);
  VNStageIntLLRInputS5xD(110)(5) <= CNStageIntLLROutputS5xD(326)(1);
  VNStageIntLLRInputS5xD(187)(4) <= CNStageIntLLROutputS5xD(326)(2);
  VNStageIntLLRInputS5xD(203)(5) <= CNStageIntLLROutputS5xD(326)(3);
  VNStageIntLLRInputS5xD(312)(4) <= CNStageIntLLROutputS5xD(326)(4);
  VNStageIntLLRInputS5xD(354)(4) <= CNStageIntLLROutputS5xD(326)(5);
  VNStageIntLLRInputS5xD(42)(5) <= CNStageIntLLROutputS5xD(327)(0);
  VNStageIntLLRInputS5xD(122)(4) <= CNStageIntLLROutputS5xD(327)(1);
  VNStageIntLLRInputS5xD(138)(5) <= CNStageIntLLROutputS5xD(327)(2);
  VNStageIntLLRInputS5xD(247)(5) <= CNStageIntLLROutputS5xD(327)(3);
  VNStageIntLLRInputS5xD(289)(5) <= CNStageIntLLROutputS5xD(327)(4);
  VNStageIntLLRInputS5xD(343)(5) <= CNStageIntLLROutputS5xD(327)(5);
  VNStageIntLLRInputS5xD(41)(5) <= CNStageIntLLROutputS5xD(328)(0);
  VNStageIntLLRInputS5xD(73)(4) <= CNStageIntLLROutputS5xD(328)(1);
  VNStageIntLLRInputS5xD(182)(5) <= CNStageIntLLROutputS5xD(328)(2);
  VNStageIntLLRInputS5xD(224)(5) <= CNStageIntLLROutputS5xD(328)(3);
  VNStageIntLLRInputS5xD(278)(4) <= CNStageIntLLROutputS5xD(328)(4);
  VNStageIntLLRInputS5xD(347)(5) <= CNStageIntLLROutputS5xD(328)(5);
  VNStageIntLLRInputS5xD(39)(5) <= CNStageIntLLROutputS5xD(329)(0);
  VNStageIntLLRInputS5xD(94)(3) <= CNStageIntLLROutputS5xD(329)(1);
  VNStageIntLLRInputS5xD(148)(5) <= CNStageIntLLROutputS5xD(329)(2);
  VNStageIntLLRInputS5xD(217)(5) <= CNStageIntLLROutputS5xD(329)(3);
  VNStageIntLLRInputS5xD(275)(4) <= CNStageIntLLROutputS5xD(329)(4);
  VNStageIntLLRInputS5xD(351)(4) <= CNStageIntLLROutputS5xD(329)(5);
  VNStageIntLLRInputS5xD(38)(5) <= CNStageIntLLROutputS5xD(330)(0);
  VNStageIntLLRInputS5xD(83)(5) <= CNStageIntLLROutputS5xD(330)(1);
  VNStageIntLLRInputS5xD(152)(5) <= CNStageIntLLROutputS5xD(330)(2);
  VNStageIntLLRInputS5xD(210)(5) <= CNStageIntLLROutputS5xD(330)(3);
  VNStageIntLLRInputS5xD(286)(5) <= CNStageIntLLROutputS5xD(330)(4);
  VNStageIntLLRInputS5xD(323)(4) <= CNStageIntLLROutputS5xD(330)(5);
  VNStageIntLLRInputS5xD(37)(5) <= CNStageIntLLROutputS5xD(331)(0);
  VNStageIntLLRInputS5xD(87)(5) <= CNStageIntLLROutputS5xD(331)(1);
  VNStageIntLLRInputS5xD(145)(5) <= CNStageIntLLROutputS5xD(331)(2);
  VNStageIntLLRInputS5xD(221)(5) <= CNStageIntLLROutputS5xD(331)(3);
  VNStageIntLLRInputS5xD(258)(2) <= CNStageIntLLROutputS5xD(331)(4);
  VNStageIntLLRInputS5xD(378)(4) <= CNStageIntLLROutputS5xD(331)(5);
  VNStageIntLLRInputS5xD(0)(5) <= CNStageIntLLROutputS5xD(332)(0);
  VNStageIntLLRInputS5xD(76)(5) <= CNStageIntLLROutputS5xD(332)(1);
  VNStageIntLLRInputS5xD(141)(3) <= CNStageIntLLROutputS5xD(332)(2);
  VNStageIntLLRInputS5xD(206)(3) <= CNStageIntLLROutputS5xD(332)(3);
  VNStageIntLLRInputS5xD(271)(4) <= CNStageIntLLROutputS5xD(332)(4);
  VNStageIntLLRInputS5xD(336)(4) <= CNStageIntLLROutputS5xD(332)(5);
  VNStageIntLLRInputS5xD(28)(5) <= CNStageIntLLROutputS5xD(333)(0);
  VNStageIntLLRInputS5xD(106)(5) <= CNStageIntLLROutputS5xD(333)(1);
  VNStageIntLLRInputS5xD(144)(6) <= CNStageIntLLROutputS5xD(333)(2);
  VNStageIntLLRInputS5xD(193)(4) <= CNStageIntLLROutputS5xD(333)(3);
  VNStageIntLLRInputS5xD(261)(5) <= CNStageIntLLROutputS5xD(333)(4);
  VNStageIntLLRInputS5xD(367)(6) <= CNStageIntLLROutputS5xD(333)(5);
  VNStageIntLLRInputS5xD(26)(6) <= CNStageIntLLROutputS5xD(334)(0);
  VNStageIntLLRInputS5xD(126)(5) <= CNStageIntLLROutputS5xD(334)(1);
  VNStageIntLLRInputS5xD(131)(5) <= CNStageIntLLROutputS5xD(334)(2);
  VNStageIntLLRInputS5xD(237)(5) <= CNStageIntLLROutputS5xD(334)(3);
  VNStageIntLLRInputS5xD(277)(6) <= CNStageIntLLROutputS5xD(334)(4);
  VNStageIntLLRInputS5xD(340)(5) <= CNStageIntLLROutputS5xD(334)(5);
  VNStageIntLLRInputS5xD(24)(6) <= CNStageIntLLROutputS5xD(335)(0);
  VNStageIntLLRInputS5xD(107)(5) <= CNStageIntLLROutputS5xD(335)(1);
  VNStageIntLLRInputS5xD(147)(6) <= CNStageIntLLROutputS5xD(335)(2);
  VNStageIntLLRInputS5xD(210)(6) <= CNStageIntLLROutputS5xD(335)(3);
  VNStageIntLLRInputS5xD(300)(5) <= CNStageIntLLROutputS5xD(335)(4);
  VNStageIntLLRInputS5xD(373)(4) <= CNStageIntLLROutputS5xD(335)(5);
  VNStageIntLLRInputS5xD(23)(6) <= CNStageIntLLROutputS5xD(336)(0);
  VNStageIntLLRInputS5xD(82)(6) <= CNStageIntLLROutputS5xD(336)(1);
  VNStageIntLLRInputS5xD(145)(6) <= CNStageIntLLROutputS5xD(336)(2);
  VNStageIntLLRInputS5xD(235)(4) <= CNStageIntLLROutputS5xD(336)(3);
  VNStageIntLLRInputS5xD(308)(4) <= CNStageIntLLROutputS5xD(336)(4);
  VNStageIntLLRInputS5xD(353)(5) <= CNStageIntLLROutputS5xD(336)(5);
  VNStageIntLLRInputS5xD(22)(6) <= CNStageIntLLROutputS5xD(337)(0);
  VNStageIntLLRInputS5xD(80)(5) <= CNStageIntLLROutputS5xD(337)(1);
  VNStageIntLLRInputS5xD(170)(4) <= CNStageIntLLROutputS5xD(337)(2);
  VNStageIntLLRInputS5xD(243)(6) <= CNStageIntLLROutputS5xD(337)(3);
  VNStageIntLLRInputS5xD(288)(6) <= CNStageIntLLROutputS5xD(337)(4);
  VNStageIntLLRInputS5xD(347)(6) <= CNStageIntLLROutputS5xD(337)(5);
  VNStageIntLLRInputS5xD(21)(6) <= CNStageIntLLROutputS5xD(338)(0);
  VNStageIntLLRInputS5xD(105)(5) <= CNStageIntLLROutputS5xD(338)(1);
  VNStageIntLLRInputS5xD(178)(5) <= CNStageIntLLROutputS5xD(338)(2);
  VNStageIntLLRInputS5xD(223)(6) <= CNStageIntLLROutputS5xD(338)(3);
  VNStageIntLLRInputS5xD(282)(5) <= CNStageIntLLROutputS5xD(338)(4);
  VNStageIntLLRInputS5xD(320)(4) <= CNStageIntLLROutputS5xD(338)(5);
  VNStageIntLLRInputS5xD(20)(4) <= CNStageIntLLROutputS5xD(339)(0);
  VNStageIntLLRInputS5xD(113)(6) <= CNStageIntLLROutputS5xD(339)(1);
  VNStageIntLLRInputS5xD(158)(6) <= CNStageIntLLROutputS5xD(339)(2);
  VNStageIntLLRInputS5xD(217)(6) <= CNStageIntLLROutputS5xD(339)(3);
  VNStageIntLLRInputS5xD(256)(5) <= CNStageIntLLROutputS5xD(339)(4);
  VNStageIntLLRInputS5xD(346)(6) <= CNStageIntLLROutputS5xD(339)(5);
  VNStageIntLLRInputS5xD(19)(4) <= CNStageIntLLROutputS5xD(340)(0);
  VNStageIntLLRInputS5xD(93)(6) <= CNStageIntLLROutputS5xD(340)(1);
  VNStageIntLLRInputS5xD(152)(6) <= CNStageIntLLROutputS5xD(340)(2);
  VNStageIntLLRInputS5xD(192)(6) <= CNStageIntLLROutputS5xD(340)(3);
  VNStageIntLLRInputS5xD(281)(6) <= CNStageIntLLROutputS5xD(340)(4);
  VNStageIntLLRInputS5xD(351)(5) <= CNStageIntLLROutputS5xD(340)(5);
  VNStageIntLLRInputS5xD(18)(6) <= CNStageIntLLROutputS5xD(341)(0);
  VNStageIntLLRInputS5xD(87)(6) <= CNStageIntLLROutputS5xD(341)(1);
  VNStageIntLLRInputS5xD(128)(6) <= CNStageIntLLROutputS5xD(341)(2);
  VNStageIntLLRInputS5xD(216)(6) <= CNStageIntLLROutputS5xD(341)(3);
  VNStageIntLLRInputS5xD(286)(6) <= CNStageIntLLROutputS5xD(341)(4);
  VNStageIntLLRInputS5xD(370)(4) <= CNStageIntLLROutputS5xD(341)(5);
  VNStageIntLLRInputS5xD(17)(6) <= CNStageIntLLROutputS5xD(342)(0);
  VNStageIntLLRInputS5xD(64)(5) <= CNStageIntLLROutputS5xD(342)(1);
  VNStageIntLLRInputS5xD(151)(5) <= CNStageIntLLROutputS5xD(342)(2);
  VNStageIntLLRInputS5xD(221)(6) <= CNStageIntLLROutputS5xD(342)(3);
  VNStageIntLLRInputS5xD(305)(6) <= CNStageIntLLROutputS5xD(342)(4);
  VNStageIntLLRInputS5xD(361)(6) <= CNStageIntLLROutputS5xD(342)(5);
  VNStageIntLLRInputS5xD(16)(5) <= CNStageIntLLROutputS5xD(343)(0);
  VNStageIntLLRInputS5xD(86)(3) <= CNStageIntLLROutputS5xD(343)(1);
  VNStageIntLLRInputS5xD(156)(3) <= CNStageIntLLROutputS5xD(343)(2);
  VNStageIntLLRInputS5xD(240)(6) <= CNStageIntLLROutputS5xD(343)(3);
  VNStageIntLLRInputS5xD(296)(5) <= CNStageIntLLROutputS5xD(343)(4);
  VNStageIntLLRInputS5xD(335)(6) <= CNStageIntLLROutputS5xD(343)(5);
  VNStageIntLLRInputS5xD(15)(6) <= CNStageIntLLROutputS5xD(344)(0);
  VNStageIntLLRInputS5xD(91)(6) <= CNStageIntLLROutputS5xD(344)(1);
  VNStageIntLLRInputS5xD(175)(6) <= CNStageIntLLROutputS5xD(344)(2);
  VNStageIntLLRInputS5xD(231)(5) <= CNStageIntLLROutputS5xD(344)(3);
  VNStageIntLLRInputS5xD(270)(6) <= CNStageIntLLROutputS5xD(344)(4);
  VNStageIntLLRInputS5xD(336)(5) <= CNStageIntLLROutputS5xD(344)(5);
  VNStageIntLLRInputS5xD(14)(6) <= CNStageIntLLROutputS5xD(345)(0);
  VNStageIntLLRInputS5xD(110)(6) <= CNStageIntLLROutputS5xD(345)(1);
  VNStageIntLLRInputS5xD(166)(5) <= CNStageIntLLROutputS5xD(345)(2);
  VNStageIntLLRInputS5xD(205)(2) <= CNStageIntLLROutputS5xD(345)(3);
  VNStageIntLLRInputS5xD(271)(5) <= CNStageIntLLROutputS5xD(345)(4);
  VNStageIntLLRInputS5xD(360)(6) <= CNStageIntLLROutputS5xD(345)(5);
  VNStageIntLLRInputS5xD(13)(5) <= CNStageIntLLROutputS5xD(346)(0);
  VNStageIntLLRInputS5xD(101)(6) <= CNStageIntLLROutputS5xD(346)(1);
  VNStageIntLLRInputS5xD(140)(6) <= CNStageIntLLROutputS5xD(346)(2);
  VNStageIntLLRInputS5xD(206)(4) <= CNStageIntLLROutputS5xD(346)(3);
  VNStageIntLLRInputS5xD(295)(4) <= CNStageIntLLROutputS5xD(346)(4);
  VNStageIntLLRInputS5xD(381)(5) <= CNStageIntLLROutputS5xD(346)(5);
  VNStageIntLLRInputS5xD(12)(6) <= CNStageIntLLROutputS5xD(347)(0);
  VNStageIntLLRInputS5xD(75)(6) <= CNStageIntLLROutputS5xD(347)(1);
  VNStageIntLLRInputS5xD(141)(4) <= CNStageIntLLROutputS5xD(347)(2);
  VNStageIntLLRInputS5xD(230)(5) <= CNStageIntLLROutputS5xD(347)(3);
  VNStageIntLLRInputS5xD(316)(4) <= CNStageIntLLROutputS5xD(347)(4);
  VNStageIntLLRInputS5xD(377)(4) <= CNStageIntLLROutputS5xD(347)(5);
  VNStageIntLLRInputS5xD(11)(5) <= CNStageIntLLROutputS5xD(348)(0);
  VNStageIntLLRInputS5xD(76)(6) <= CNStageIntLLROutputS5xD(348)(1);
  VNStageIntLLRInputS5xD(165)(5) <= CNStageIntLLROutputS5xD(348)(2);
  VNStageIntLLRInputS5xD(251)(4) <= CNStageIntLLROutputS5xD(348)(3);
  VNStageIntLLRInputS5xD(312)(5) <= CNStageIntLLROutputS5xD(348)(4);
  VNStageIntLLRInputS5xD(329)(6) <= CNStageIntLLROutputS5xD(348)(5);
  VNStageIntLLRInputS5xD(10)(4) <= CNStageIntLLROutputS5xD(349)(0);
  VNStageIntLLRInputS5xD(100)(6) <= CNStageIntLLROutputS5xD(349)(1);
  VNStageIntLLRInputS5xD(186)(5) <= CNStageIntLLROutputS5xD(349)(2);
  VNStageIntLLRInputS5xD(247)(6) <= CNStageIntLLROutputS5xD(349)(3);
  VNStageIntLLRInputS5xD(264)(6) <= CNStageIntLLROutputS5xD(349)(4);
  VNStageIntLLRInputS5xD(355)(6) <= CNStageIntLLROutputS5xD(349)(5);
  VNStageIntLLRInputS5xD(9)(6) <= CNStageIntLLROutputS5xD(350)(0);
  VNStageIntLLRInputS5xD(121)(5) <= CNStageIntLLROutputS5xD(350)(1);
  VNStageIntLLRInputS5xD(182)(6) <= CNStageIntLLROutputS5xD(350)(2);
  VNStageIntLLRInputS5xD(199)(6) <= CNStageIntLLROutputS5xD(350)(3);
  VNStageIntLLRInputS5xD(290)(5) <= CNStageIntLLROutputS5xD(350)(4);
  VNStageIntLLRInputS5xD(331)(4) <= CNStageIntLLROutputS5xD(350)(5);
  VNStageIntLLRInputS5xD(7)(6) <= CNStageIntLLROutputS5xD(351)(0);
  VNStageIntLLRInputS5xD(69)(6) <= CNStageIntLLROutputS5xD(351)(1);
  VNStageIntLLRInputS5xD(160)(6) <= CNStageIntLLROutputS5xD(351)(2);
  VNStageIntLLRInputS5xD(201)(5) <= CNStageIntLLROutputS5xD(351)(3);
  VNStageIntLLRInputS5xD(298)(6) <= CNStageIntLLROutputS5xD(351)(4);
  VNStageIntLLRInputS5xD(379)(4) <= CNStageIntLLROutputS5xD(351)(5);
  VNStageIntLLRInputS5xD(6)(6) <= CNStageIntLLROutputS5xD(352)(0);
  VNStageIntLLRInputS5xD(95)(6) <= CNStageIntLLROutputS5xD(352)(1);
  VNStageIntLLRInputS5xD(136)(6) <= CNStageIntLLROutputS5xD(352)(2);
  VNStageIntLLRInputS5xD(233)(4) <= CNStageIntLLROutputS5xD(352)(3);
  VNStageIntLLRInputS5xD(314)(3) <= CNStageIntLLROutputS5xD(352)(4);
  VNStageIntLLRInputS5xD(349)(5) <= CNStageIntLLROutputS5xD(352)(5);
  VNStageIntLLRInputS5xD(5)(6) <= CNStageIntLLROutputS5xD(353)(0);
  VNStageIntLLRInputS5xD(71)(5) <= CNStageIntLLROutputS5xD(353)(1);
  VNStageIntLLRInputS5xD(168)(5) <= CNStageIntLLROutputS5xD(353)(2);
  VNStageIntLLRInputS5xD(249)(4) <= CNStageIntLLROutputS5xD(353)(3);
  VNStageIntLLRInputS5xD(284)(6) <= CNStageIntLLROutputS5xD(353)(4);
  VNStageIntLLRInputS5xD(358)(5) <= CNStageIntLLROutputS5xD(353)(5);
  VNStageIntLLRInputS5xD(4)(5) <= CNStageIntLLROutputS5xD(354)(0);
  VNStageIntLLRInputS5xD(103)(6) <= CNStageIntLLROutputS5xD(354)(1);
  VNStageIntLLRInputS5xD(184)(6) <= CNStageIntLLROutputS5xD(354)(2);
  VNStageIntLLRInputS5xD(219)(5) <= CNStageIntLLROutputS5xD(354)(3);
  VNStageIntLLRInputS5xD(293)(5) <= CNStageIntLLROutputS5xD(354)(4);
  VNStageIntLLRInputS5xD(371)(4) <= CNStageIntLLROutputS5xD(354)(5);
  VNStageIntLLRInputS5xD(2)(6) <= CNStageIntLLROutputS5xD(355)(0);
  VNStageIntLLRInputS5xD(89)(5) <= CNStageIntLLROutputS5xD(355)(1);
  VNStageIntLLRInputS5xD(163)(4) <= CNStageIntLLROutputS5xD(355)(2);
  VNStageIntLLRInputS5xD(241)(5) <= CNStageIntLLROutputS5xD(355)(3);
  VNStageIntLLRInputS5xD(285)(6) <= CNStageIntLLROutputS5xD(355)(4);
  VNStageIntLLRInputS5xD(378)(5) <= CNStageIntLLROutputS5xD(355)(5);
  VNStageIntLLRInputS5xD(1)(5) <= CNStageIntLLROutputS5xD(356)(0);
  VNStageIntLLRInputS5xD(98)(5) <= CNStageIntLLROutputS5xD(356)(1);
  VNStageIntLLRInputS5xD(176)(6) <= CNStageIntLLROutputS5xD(356)(2);
  VNStageIntLLRInputS5xD(220)(6) <= CNStageIntLLROutputS5xD(356)(3);
  VNStageIntLLRInputS5xD(313)(3) <= CNStageIntLLROutputS5xD(356)(4);
  VNStageIntLLRInputS5xD(380)(5) <= CNStageIntLLROutputS5xD(356)(5);
  VNStageIntLLRInputS5xD(63)(3) <= CNStageIntLLROutputS5xD(357)(0);
  VNStageIntLLRInputS5xD(111)(6) <= CNStageIntLLROutputS5xD(357)(1);
  VNStageIntLLRInputS5xD(155)(6) <= CNStageIntLLROutputS5xD(357)(2);
  VNStageIntLLRInputS5xD(248)(6) <= CNStageIntLLROutputS5xD(357)(3);
  VNStageIntLLRInputS5xD(315)(5) <= CNStageIntLLROutputS5xD(357)(4);
  VNStageIntLLRInputS5xD(362)(6) <= CNStageIntLLROutputS5xD(357)(5);
  VNStageIntLLRInputS5xD(62)(5) <= CNStageIntLLROutputS5xD(358)(0);
  VNStageIntLLRInputS5xD(90)(6) <= CNStageIntLLROutputS5xD(358)(1);
  VNStageIntLLRInputS5xD(183)(4) <= CNStageIntLLROutputS5xD(358)(2);
  VNStageIntLLRInputS5xD(250)(4) <= CNStageIntLLROutputS5xD(358)(3);
  VNStageIntLLRInputS5xD(297)(6) <= CNStageIntLLROutputS5xD(358)(4);
  VNStageIntLLRInputS5xD(369)(4) <= CNStageIntLLROutputS5xD(358)(5);
  VNStageIntLLRInputS5xD(61)(5) <= CNStageIntLLROutputS5xD(359)(0);
  VNStageIntLLRInputS5xD(118)(5) <= CNStageIntLLROutputS5xD(359)(1);
  VNStageIntLLRInputS5xD(185)(3) <= CNStageIntLLROutputS5xD(359)(2);
  VNStageIntLLRInputS5xD(232)(5) <= CNStageIntLLROutputS5xD(359)(3);
  VNStageIntLLRInputS5xD(304)(6) <= CNStageIntLLROutputS5xD(359)(4);
  VNStageIntLLRInputS5xD(333)(5) <= CNStageIntLLROutputS5xD(359)(5);
  VNStageIntLLRInputS5xD(60)(5) <= CNStageIntLLROutputS5xD(360)(0);
  VNStageIntLLRInputS5xD(120)(3) <= CNStageIntLLROutputS5xD(360)(1);
  VNStageIntLLRInputS5xD(167)(6) <= CNStageIntLLROutputS5xD(360)(2);
  VNStageIntLLRInputS5xD(239)(6) <= CNStageIntLLROutputS5xD(360)(3);
  VNStageIntLLRInputS5xD(268)(6) <= CNStageIntLLROutputS5xD(360)(4);
  VNStageIntLLRInputS5xD(321)(6) <= CNStageIntLLROutputS5xD(360)(5);
  VNStageIntLLRInputS5xD(59)(4) <= CNStageIntLLROutputS5xD(361)(0);
  VNStageIntLLRInputS5xD(102)(5) <= CNStageIntLLROutputS5xD(361)(1);
  VNStageIntLLRInputS5xD(174)(4) <= CNStageIntLLROutputS5xD(361)(2);
  VNStageIntLLRInputS5xD(203)(6) <= CNStageIntLLROutputS5xD(361)(3);
  VNStageIntLLRInputS5xD(319)(6) <= CNStageIntLLROutputS5xD(361)(4);
  VNStageIntLLRInputS5xD(327)(6) <= CNStageIntLLROutputS5xD(361)(5);
  VNStageIntLLRInputS5xD(58)(4) <= CNStageIntLLROutputS5xD(362)(0);
  VNStageIntLLRInputS5xD(109)(5) <= CNStageIntLLROutputS5xD(362)(1);
  VNStageIntLLRInputS5xD(138)(6) <= CNStageIntLLROutputS5xD(362)(2);
  VNStageIntLLRInputS5xD(254)(4) <= CNStageIntLLROutputS5xD(362)(3);
  VNStageIntLLRInputS5xD(262)(5) <= CNStageIntLLROutputS5xD(362)(4);
  VNStageIntLLRInputS5xD(322)(5) <= CNStageIntLLROutputS5xD(362)(5);
  VNStageIntLLRInputS5xD(57)(5) <= CNStageIntLLROutputS5xD(363)(0);
  VNStageIntLLRInputS5xD(73)(5) <= CNStageIntLLROutputS5xD(363)(1);
  VNStageIntLLRInputS5xD(189)(5) <= CNStageIntLLROutputS5xD(363)(2);
  VNStageIntLLRInputS5xD(197)(6) <= CNStageIntLLROutputS5xD(363)(3);
  VNStageIntLLRInputS5xD(257)(6) <= CNStageIntLLROutputS5xD(363)(4);
  VNStageIntLLRInputS5xD(332)(5) <= CNStageIntLLROutputS5xD(363)(5);
  VNStageIntLLRInputS5xD(56)(6) <= CNStageIntLLROutputS5xD(364)(0);
  VNStageIntLLRInputS5xD(124)(4) <= CNStageIntLLROutputS5xD(364)(1);
  VNStageIntLLRInputS5xD(132)(5) <= CNStageIntLLROutputS5xD(364)(2);
  VNStageIntLLRInputS5xD(255)(6) <= CNStageIntLLROutputS5xD(364)(3);
  VNStageIntLLRInputS5xD(267)(6) <= CNStageIntLLROutputS5xD(364)(4);
  VNStageIntLLRInputS5xD(354)(5) <= CNStageIntLLROutputS5xD(364)(5);
  VNStageIntLLRInputS5xD(55)(6) <= CNStageIntLLROutputS5xD(365)(0);
  VNStageIntLLRInputS5xD(67)(3) <= CNStageIntLLROutputS5xD(365)(1);
  VNStageIntLLRInputS5xD(190)(4) <= CNStageIntLLROutputS5xD(365)(2);
  VNStageIntLLRInputS5xD(202)(5) <= CNStageIntLLROutputS5xD(365)(3);
  VNStageIntLLRInputS5xD(289)(6) <= CNStageIntLLROutputS5xD(365)(4);
  VNStageIntLLRInputS5xD(372)(5) <= CNStageIntLLROutputS5xD(365)(5);
  VNStageIntLLRInputS5xD(54)(5) <= CNStageIntLLROutputS5xD(366)(0);
  VNStageIntLLRInputS5xD(125)(3) <= CNStageIntLLROutputS5xD(366)(1);
  VNStageIntLLRInputS5xD(137)(6) <= CNStageIntLLROutputS5xD(366)(2);
  VNStageIntLLRInputS5xD(224)(6) <= CNStageIntLLROutputS5xD(366)(3);
  VNStageIntLLRInputS5xD(307)(6) <= CNStageIntLLROutputS5xD(366)(4);
  VNStageIntLLRInputS5xD(357)(6) <= CNStageIntLLROutputS5xD(366)(5);
  VNStageIntLLRInputS5xD(53)(5) <= CNStageIntLLROutputS5xD(367)(0);
  VNStageIntLLRInputS5xD(72)(5) <= CNStageIntLLROutputS5xD(367)(1);
  VNStageIntLLRInputS5xD(159)(4) <= CNStageIntLLROutputS5xD(367)(2);
  VNStageIntLLRInputS5xD(242)(6) <= CNStageIntLLROutputS5xD(367)(3);
  VNStageIntLLRInputS5xD(292)(6) <= CNStageIntLLROutputS5xD(367)(4);
  VNStageIntLLRInputS5xD(344)(6) <= CNStageIntLLROutputS5xD(367)(5);
  VNStageIntLLRInputS5xD(52)(4) <= CNStageIntLLROutputS5xD(368)(0);
  VNStageIntLLRInputS5xD(94)(4) <= CNStageIntLLROutputS5xD(368)(1);
  VNStageIntLLRInputS5xD(177)(6) <= CNStageIntLLROutputS5xD(368)(2);
  VNStageIntLLRInputS5xD(227)(6) <= CNStageIntLLROutputS5xD(368)(3);
  VNStageIntLLRInputS5xD(279)(5) <= CNStageIntLLROutputS5xD(368)(4);
  VNStageIntLLRInputS5xD(375)(5) <= CNStageIntLLROutputS5xD(368)(5);
  VNStageIntLLRInputS5xD(51)(5) <= CNStageIntLLROutputS5xD(369)(0);
  VNStageIntLLRInputS5xD(112)(6) <= CNStageIntLLROutputS5xD(369)(1);
  VNStageIntLLRInputS5xD(162)(6) <= CNStageIntLLROutputS5xD(369)(2);
  VNStageIntLLRInputS5xD(214)(6) <= CNStageIntLLROutputS5xD(369)(3);
  VNStageIntLLRInputS5xD(310)(5) <= CNStageIntLLROutputS5xD(369)(4);
  VNStageIntLLRInputS5xD(324)(6) <= CNStageIntLLROutputS5xD(369)(5);
  VNStageIntLLRInputS5xD(50)(6) <= CNStageIntLLROutputS5xD(370)(0);
  VNStageIntLLRInputS5xD(97)(6) <= CNStageIntLLROutputS5xD(370)(1);
  VNStageIntLLRInputS5xD(149)(6) <= CNStageIntLLROutputS5xD(370)(2);
  VNStageIntLLRInputS5xD(245)(6) <= CNStageIntLLROutputS5xD(370)(3);
  VNStageIntLLRInputS5xD(259)(4) <= CNStageIntLLROutputS5xD(370)(4);
  VNStageIntLLRInputS5xD(338)(4) <= CNStageIntLLROutputS5xD(370)(5);
  VNStageIntLLRInputS5xD(49)(6) <= CNStageIntLLROutputS5xD(371)(0);
  VNStageIntLLRInputS5xD(84)(5) <= CNStageIntLLROutputS5xD(371)(1);
  VNStageIntLLRInputS5xD(180)(4) <= CNStageIntLLROutputS5xD(371)(2);
  VNStageIntLLRInputS5xD(194)(6) <= CNStageIntLLROutputS5xD(371)(3);
  VNStageIntLLRInputS5xD(273)(5) <= CNStageIntLLROutputS5xD(371)(4);
  VNStageIntLLRInputS5xD(382)(5) <= CNStageIntLLROutputS5xD(371)(5);
  VNStageIntLLRInputS5xD(48)(3) <= CNStageIntLLROutputS5xD(372)(0);
  VNStageIntLLRInputS5xD(115)(6) <= CNStageIntLLROutputS5xD(372)(1);
  VNStageIntLLRInputS5xD(129)(6) <= CNStageIntLLROutputS5xD(372)(2);
  VNStageIntLLRInputS5xD(208)(5) <= CNStageIntLLROutputS5xD(372)(3);
  VNStageIntLLRInputS5xD(317)(3) <= CNStageIntLLROutputS5xD(372)(4);
  VNStageIntLLRInputS5xD(359)(6) <= CNStageIntLLROutputS5xD(372)(5);
  VNStageIntLLRInputS5xD(47)(3) <= CNStageIntLLROutputS5xD(373)(0);
  VNStageIntLLRInputS5xD(127)(6) <= CNStageIntLLROutputS5xD(373)(1);
  VNStageIntLLRInputS5xD(143)(6) <= CNStageIntLLROutputS5xD(373)(2);
  VNStageIntLLRInputS5xD(252)(5) <= CNStageIntLLROutputS5xD(373)(3);
  VNStageIntLLRInputS5xD(294)(6) <= CNStageIntLLROutputS5xD(373)(4);
  VNStageIntLLRInputS5xD(348)(6) <= CNStageIntLLROutputS5xD(373)(5);
  VNStageIntLLRInputS5xD(46)(6) <= CNStageIntLLROutputS5xD(374)(0);
  VNStageIntLLRInputS5xD(78)(6) <= CNStageIntLLROutputS5xD(374)(1);
  VNStageIntLLRInputS5xD(187)(5) <= CNStageIntLLROutputS5xD(374)(2);
  VNStageIntLLRInputS5xD(229)(4) <= CNStageIntLLROutputS5xD(374)(3);
  VNStageIntLLRInputS5xD(283)(6) <= CNStageIntLLROutputS5xD(374)(4);
  VNStageIntLLRInputS5xD(352)(6) <= CNStageIntLLROutputS5xD(374)(5);
  VNStageIntLLRInputS5xD(45)(6) <= CNStageIntLLROutputS5xD(375)(0);
  VNStageIntLLRInputS5xD(122)(5) <= CNStageIntLLROutputS5xD(375)(1);
  VNStageIntLLRInputS5xD(164)(5) <= CNStageIntLLROutputS5xD(375)(2);
  VNStageIntLLRInputS5xD(218)(6) <= CNStageIntLLROutputS5xD(375)(3);
  VNStageIntLLRInputS5xD(287)(6) <= CNStageIntLLROutputS5xD(375)(4);
  VNStageIntLLRInputS5xD(345)(5) <= CNStageIntLLROutputS5xD(375)(5);
  VNStageIntLLRInputS5xD(44)(6) <= CNStageIntLLROutputS5xD(376)(0);
  VNStageIntLLRInputS5xD(99)(6) <= CNStageIntLLROutputS5xD(376)(1);
  VNStageIntLLRInputS5xD(153)(6) <= CNStageIntLLROutputS5xD(376)(2);
  VNStageIntLLRInputS5xD(222)(3) <= CNStageIntLLROutputS5xD(376)(3);
  VNStageIntLLRInputS5xD(280)(6) <= CNStageIntLLROutputS5xD(376)(4);
  VNStageIntLLRInputS5xD(356)(5) <= CNStageIntLLROutputS5xD(376)(5);
  VNStageIntLLRInputS5xD(43)(5) <= CNStageIntLLROutputS5xD(377)(0);
  VNStageIntLLRInputS5xD(88)(6) <= CNStageIntLLROutputS5xD(377)(1);
  VNStageIntLLRInputS5xD(157)(5) <= CNStageIntLLROutputS5xD(377)(2);
  VNStageIntLLRInputS5xD(215)(6) <= CNStageIntLLROutputS5xD(377)(3);
  VNStageIntLLRInputS5xD(291)(5) <= CNStageIntLLROutputS5xD(377)(4);
  VNStageIntLLRInputS5xD(328)(4) <= CNStageIntLLROutputS5xD(377)(5);
  VNStageIntLLRInputS5xD(42)(6) <= CNStageIntLLROutputS5xD(378)(0);
  VNStageIntLLRInputS5xD(92)(6) <= CNStageIntLLROutputS5xD(378)(1);
  VNStageIntLLRInputS5xD(150)(5) <= CNStageIntLLROutputS5xD(378)(2);
  VNStageIntLLRInputS5xD(226)(2) <= CNStageIntLLROutputS5xD(378)(3);
  VNStageIntLLRInputS5xD(263)(6) <= CNStageIntLLROutputS5xD(378)(4);
  VNStageIntLLRInputS5xD(383)(6) <= CNStageIntLLROutputS5xD(378)(5);
  VNStageIntLLRInputS5xD(41)(6) <= CNStageIntLLROutputS5xD(379)(0);
  VNStageIntLLRInputS5xD(85)(5) <= CNStageIntLLROutputS5xD(379)(1);
  VNStageIntLLRInputS5xD(161)(6) <= CNStageIntLLROutputS5xD(379)(2);
  VNStageIntLLRInputS5xD(198)(6) <= CNStageIntLLROutputS5xD(379)(3);
  VNStageIntLLRInputS5xD(318)(3) <= CNStageIntLLROutputS5xD(379)(4);
  VNStageIntLLRInputS5xD(337)(6) <= CNStageIntLLROutputS5xD(379)(5);
  VNStageIntLLRInputS5xD(40)(4) <= CNStageIntLLROutputS5xD(380)(0);
  VNStageIntLLRInputS5xD(96)(5) <= CNStageIntLLROutputS5xD(380)(1);
  VNStageIntLLRInputS5xD(133)(4) <= CNStageIntLLROutputS5xD(380)(2);
  VNStageIntLLRInputS5xD(253)(5) <= CNStageIntLLROutputS5xD(380)(3);
  VNStageIntLLRInputS5xD(272)(6) <= CNStageIntLLROutputS5xD(380)(4);
  VNStageIntLLRInputS5xD(334)(4) <= CNStageIntLLROutputS5xD(380)(5);
  VNStageIntLLRInputS5xD(39)(6) <= CNStageIntLLROutputS5xD(381)(0);
  VNStageIntLLRInputS5xD(68)(5) <= CNStageIntLLROutputS5xD(381)(1);
  VNStageIntLLRInputS5xD(188)(4) <= CNStageIntLLROutputS5xD(381)(2);
  VNStageIntLLRInputS5xD(207)(5) <= CNStageIntLLROutputS5xD(381)(3);
  VNStageIntLLRInputS5xD(269)(5) <= CNStageIntLLROutputS5xD(381)(4);
  VNStageIntLLRInputS5xD(368)(2) <= CNStageIntLLROutputS5xD(381)(5);
  VNStageIntLLRInputS5xD(38)(6) <= CNStageIntLLROutputS5xD(382)(0);
  VNStageIntLLRInputS5xD(123)(4) <= CNStageIntLLROutputS5xD(382)(1);
  VNStageIntLLRInputS5xD(142)(4) <= CNStageIntLLROutputS5xD(382)(2);
  VNStageIntLLRInputS5xD(204)(6) <= CNStageIntLLROutputS5xD(382)(3);
  VNStageIntLLRInputS5xD(303)(6) <= CNStageIntLLROutputS5xD(382)(4);
  VNStageIntLLRInputS5xD(325)(6) <= CNStageIntLLROutputS5xD(382)(5);
  VNStageIntLLRInputS5xD(37)(6) <= CNStageIntLLROutputS5xD(383)(0);
  VNStageIntLLRInputS5xD(77)(4) <= CNStageIntLLROutputS5xD(383)(1);
  VNStageIntLLRInputS5xD(139)(6) <= CNStageIntLLROutputS5xD(383)(2);
  VNStageIntLLRInputS5xD(238)(6) <= CNStageIntLLROutputS5xD(383)(3);
  VNStageIntLLRInputS5xD(260)(5) <= CNStageIntLLROutputS5xD(383)(4);
  VNStageIntLLRInputS5xD(374)(6) <= CNStageIntLLROutputS5xD(383)(5);

  -- Check Nodes (Iteration 6)
  CNStageIntLLRInputS6xD(53)(0) <= VNStageIntLLROutputS5xD(0)(0);
  CNStageIntLLRInputS6xD(110)(0) <= VNStageIntLLROutputS5xD(0)(1);
  CNStageIntLLRInputS6xD(170)(0) <= VNStageIntLLROutputS5xD(0)(2);
  CNStageIntLLRInputS6xD(224)(0) <= VNStageIntLLROutputS5xD(0)(3);
  CNStageIntLLRInputS6xD(279)(0) <= VNStageIntLLROutputS5xD(0)(4);
  CNStageIntLLRInputS6xD(332)(0) <= VNStageIntLLROutputS5xD(0)(5);
  CNStageIntLLRInputS6xD(51)(0) <= VNStageIntLLROutputS5xD(1)(0);
  CNStageIntLLRInputS6xD(139)(0) <= VNStageIntLLROutputS5xD(1)(1);
  CNStageIntLLRInputS6xD(223)(0) <= VNStageIntLLROutputS5xD(1)(2);
  CNStageIntLLRInputS6xD(241)(0) <= VNStageIntLLROutputS5xD(1)(3);
  CNStageIntLLRInputS6xD(307)(0) <= VNStageIntLLROutputS5xD(1)(4);
  CNStageIntLLRInputS6xD(356)(0) <= VNStageIntLLROutputS5xD(1)(5);
  CNStageIntLLRInputS6xD(50)(0) <= VNStageIntLLROutputS5xD(2)(0);
  CNStageIntLLRInputS6xD(92)(0) <= VNStageIntLLROutputS5xD(2)(1);
  CNStageIntLLRInputS6xD(138)(0) <= VNStageIntLLROutputS5xD(2)(2);
  CNStageIntLLRInputS6xD(222)(0) <= VNStageIntLLROutputS5xD(2)(3);
  CNStageIntLLRInputS6xD(240)(0) <= VNStageIntLLROutputS5xD(2)(4);
  CNStageIntLLRInputS6xD(306)(0) <= VNStageIntLLROutputS5xD(2)(5);
  CNStageIntLLRInputS6xD(355)(0) <= VNStageIntLLROutputS5xD(2)(6);
  CNStageIntLLRInputS6xD(91)(0) <= VNStageIntLLROutputS5xD(3)(0);
  CNStageIntLLRInputS6xD(137)(0) <= VNStageIntLLROutputS5xD(3)(1);
  CNStageIntLLRInputS6xD(221)(0) <= VNStageIntLLROutputS5xD(3)(2);
  CNStageIntLLRInputS6xD(239)(0) <= VNStageIntLLROutputS5xD(3)(3);
  CNStageIntLLRInputS6xD(305)(0) <= VNStageIntLLROutputS5xD(3)(4);
  CNStageIntLLRInputS6xD(49)(0) <= VNStageIntLLROutputS5xD(4)(0);
  CNStageIntLLRInputS6xD(90)(0) <= VNStageIntLLROutputS5xD(4)(1);
  CNStageIntLLRInputS6xD(220)(0) <= VNStageIntLLROutputS5xD(4)(2);
  CNStageIntLLRInputS6xD(238)(0) <= VNStageIntLLROutputS5xD(4)(3);
  CNStageIntLLRInputS6xD(304)(0) <= VNStageIntLLROutputS5xD(4)(4);
  CNStageIntLLRInputS6xD(354)(0) <= VNStageIntLLROutputS5xD(4)(5);
  CNStageIntLLRInputS6xD(48)(0) <= VNStageIntLLROutputS5xD(5)(0);
  CNStageIntLLRInputS6xD(89)(0) <= VNStageIntLLROutputS5xD(5)(1);
  CNStageIntLLRInputS6xD(136)(0) <= VNStageIntLLROutputS5xD(5)(2);
  CNStageIntLLRInputS6xD(219)(0) <= VNStageIntLLROutputS5xD(5)(3);
  CNStageIntLLRInputS6xD(237)(0) <= VNStageIntLLROutputS5xD(5)(4);
  CNStageIntLLRInputS6xD(303)(0) <= VNStageIntLLROutputS5xD(5)(5);
  CNStageIntLLRInputS6xD(353)(0) <= VNStageIntLLROutputS5xD(5)(6);
  CNStageIntLLRInputS6xD(47)(0) <= VNStageIntLLROutputS5xD(6)(0);
  CNStageIntLLRInputS6xD(88)(0) <= VNStageIntLLROutputS5xD(6)(1);
  CNStageIntLLRInputS6xD(135)(0) <= VNStageIntLLROutputS5xD(6)(2);
  CNStageIntLLRInputS6xD(218)(0) <= VNStageIntLLROutputS5xD(6)(3);
  CNStageIntLLRInputS6xD(236)(0) <= VNStageIntLLROutputS5xD(6)(4);
  CNStageIntLLRInputS6xD(302)(0) <= VNStageIntLLROutputS5xD(6)(5);
  CNStageIntLLRInputS6xD(352)(0) <= VNStageIntLLROutputS5xD(6)(6);
  CNStageIntLLRInputS6xD(46)(0) <= VNStageIntLLROutputS5xD(7)(0);
  CNStageIntLLRInputS6xD(87)(0) <= VNStageIntLLROutputS5xD(7)(1);
  CNStageIntLLRInputS6xD(134)(0) <= VNStageIntLLROutputS5xD(7)(2);
  CNStageIntLLRInputS6xD(217)(0) <= VNStageIntLLROutputS5xD(7)(3);
  CNStageIntLLRInputS6xD(235)(0) <= VNStageIntLLROutputS5xD(7)(4);
  CNStageIntLLRInputS6xD(301)(0) <= VNStageIntLLROutputS5xD(7)(5);
  CNStageIntLLRInputS6xD(351)(0) <= VNStageIntLLROutputS5xD(7)(6);
  CNStageIntLLRInputS6xD(45)(0) <= VNStageIntLLROutputS5xD(8)(0);
  CNStageIntLLRInputS6xD(133)(0) <= VNStageIntLLROutputS5xD(8)(1);
  CNStageIntLLRInputS6xD(216)(0) <= VNStageIntLLROutputS5xD(8)(2);
  CNStageIntLLRInputS6xD(44)(0) <= VNStageIntLLROutputS5xD(9)(0);
  CNStageIntLLRInputS6xD(86)(0) <= VNStageIntLLROutputS5xD(9)(1);
  CNStageIntLLRInputS6xD(132)(0) <= VNStageIntLLROutputS5xD(9)(2);
  CNStageIntLLRInputS6xD(215)(0) <= VNStageIntLLROutputS5xD(9)(3);
  CNStageIntLLRInputS6xD(234)(0) <= VNStageIntLLROutputS5xD(9)(4);
  CNStageIntLLRInputS6xD(300)(0) <= VNStageIntLLROutputS5xD(9)(5);
  CNStageIntLLRInputS6xD(350)(0) <= VNStageIntLLROutputS5xD(9)(6);
  CNStageIntLLRInputS6xD(43)(0) <= VNStageIntLLROutputS5xD(10)(0);
  CNStageIntLLRInputS6xD(85)(0) <= VNStageIntLLROutputS5xD(10)(1);
  CNStageIntLLRInputS6xD(131)(0) <= VNStageIntLLROutputS5xD(10)(2);
  CNStageIntLLRInputS6xD(233)(0) <= VNStageIntLLROutputS5xD(10)(3);
  CNStageIntLLRInputS6xD(349)(0) <= VNStageIntLLROutputS5xD(10)(4);
  CNStageIntLLRInputS6xD(42)(0) <= VNStageIntLLROutputS5xD(11)(0);
  CNStageIntLLRInputS6xD(84)(0) <= VNStageIntLLROutputS5xD(11)(1);
  CNStageIntLLRInputS6xD(130)(0) <= VNStageIntLLROutputS5xD(11)(2);
  CNStageIntLLRInputS6xD(214)(0) <= VNStageIntLLROutputS5xD(11)(3);
  CNStageIntLLRInputS6xD(232)(0) <= VNStageIntLLROutputS5xD(11)(4);
  CNStageIntLLRInputS6xD(348)(0) <= VNStageIntLLROutputS5xD(11)(5);
  CNStageIntLLRInputS6xD(41)(0) <= VNStageIntLLROutputS5xD(12)(0);
  CNStageIntLLRInputS6xD(83)(0) <= VNStageIntLLROutputS5xD(12)(1);
  CNStageIntLLRInputS6xD(129)(0) <= VNStageIntLLROutputS5xD(12)(2);
  CNStageIntLLRInputS6xD(213)(0) <= VNStageIntLLROutputS5xD(12)(3);
  CNStageIntLLRInputS6xD(231)(0) <= VNStageIntLLROutputS5xD(12)(4);
  CNStageIntLLRInputS6xD(299)(0) <= VNStageIntLLROutputS5xD(12)(5);
  CNStageIntLLRInputS6xD(347)(0) <= VNStageIntLLROutputS5xD(12)(6);
  CNStageIntLLRInputS6xD(82)(0) <= VNStageIntLLROutputS5xD(13)(0);
  CNStageIntLLRInputS6xD(128)(0) <= VNStageIntLLROutputS5xD(13)(1);
  CNStageIntLLRInputS6xD(212)(0) <= VNStageIntLLROutputS5xD(13)(2);
  CNStageIntLLRInputS6xD(230)(0) <= VNStageIntLLROutputS5xD(13)(3);
  CNStageIntLLRInputS6xD(298)(0) <= VNStageIntLLROutputS5xD(13)(4);
  CNStageIntLLRInputS6xD(346)(0) <= VNStageIntLLROutputS5xD(13)(5);
  CNStageIntLLRInputS6xD(40)(0) <= VNStageIntLLROutputS5xD(14)(0);
  CNStageIntLLRInputS6xD(81)(0) <= VNStageIntLLROutputS5xD(14)(1);
  CNStageIntLLRInputS6xD(127)(0) <= VNStageIntLLROutputS5xD(14)(2);
  CNStageIntLLRInputS6xD(211)(0) <= VNStageIntLLROutputS5xD(14)(3);
  CNStageIntLLRInputS6xD(229)(0) <= VNStageIntLLROutputS5xD(14)(4);
  CNStageIntLLRInputS6xD(297)(0) <= VNStageIntLLROutputS5xD(14)(5);
  CNStageIntLLRInputS6xD(345)(0) <= VNStageIntLLROutputS5xD(14)(6);
  CNStageIntLLRInputS6xD(39)(0) <= VNStageIntLLROutputS5xD(15)(0);
  CNStageIntLLRInputS6xD(80)(0) <= VNStageIntLLROutputS5xD(15)(1);
  CNStageIntLLRInputS6xD(126)(0) <= VNStageIntLLROutputS5xD(15)(2);
  CNStageIntLLRInputS6xD(210)(0) <= VNStageIntLLROutputS5xD(15)(3);
  CNStageIntLLRInputS6xD(228)(0) <= VNStageIntLLROutputS5xD(15)(4);
  CNStageIntLLRInputS6xD(296)(0) <= VNStageIntLLROutputS5xD(15)(5);
  CNStageIntLLRInputS6xD(344)(0) <= VNStageIntLLROutputS5xD(15)(6);
  CNStageIntLLRInputS6xD(38)(0) <= VNStageIntLLROutputS5xD(16)(0);
  CNStageIntLLRInputS6xD(125)(0) <= VNStageIntLLROutputS5xD(16)(1);
  CNStageIntLLRInputS6xD(209)(0) <= VNStageIntLLROutputS5xD(16)(2);
  CNStageIntLLRInputS6xD(227)(0) <= VNStageIntLLROutputS5xD(16)(3);
  CNStageIntLLRInputS6xD(295)(0) <= VNStageIntLLROutputS5xD(16)(4);
  CNStageIntLLRInputS6xD(343)(0) <= VNStageIntLLROutputS5xD(16)(5);
  CNStageIntLLRInputS6xD(37)(0) <= VNStageIntLLROutputS5xD(17)(0);
  CNStageIntLLRInputS6xD(79)(0) <= VNStageIntLLROutputS5xD(17)(1);
  CNStageIntLLRInputS6xD(124)(0) <= VNStageIntLLROutputS5xD(17)(2);
  CNStageIntLLRInputS6xD(208)(0) <= VNStageIntLLROutputS5xD(17)(3);
  CNStageIntLLRInputS6xD(226)(0) <= VNStageIntLLROutputS5xD(17)(4);
  CNStageIntLLRInputS6xD(294)(0) <= VNStageIntLLROutputS5xD(17)(5);
  CNStageIntLLRInputS6xD(342)(0) <= VNStageIntLLROutputS5xD(17)(6);
  CNStageIntLLRInputS6xD(36)(0) <= VNStageIntLLROutputS5xD(18)(0);
  CNStageIntLLRInputS6xD(78)(0) <= VNStageIntLLROutputS5xD(18)(1);
  CNStageIntLLRInputS6xD(123)(0) <= VNStageIntLLROutputS5xD(18)(2);
  CNStageIntLLRInputS6xD(207)(0) <= VNStageIntLLROutputS5xD(18)(3);
  CNStageIntLLRInputS6xD(225)(0) <= VNStageIntLLROutputS5xD(18)(4);
  CNStageIntLLRInputS6xD(293)(0) <= VNStageIntLLROutputS5xD(18)(5);
  CNStageIntLLRInputS6xD(341)(0) <= VNStageIntLLROutputS5xD(18)(6);
  CNStageIntLLRInputS6xD(35)(0) <= VNStageIntLLROutputS5xD(19)(0);
  CNStageIntLLRInputS6xD(77)(0) <= VNStageIntLLROutputS5xD(19)(1);
  CNStageIntLLRInputS6xD(122)(0) <= VNStageIntLLROutputS5xD(19)(2);
  CNStageIntLLRInputS6xD(278)(0) <= VNStageIntLLROutputS5xD(19)(3);
  CNStageIntLLRInputS6xD(340)(0) <= VNStageIntLLROutputS5xD(19)(4);
  CNStageIntLLRInputS6xD(34)(0) <= VNStageIntLLROutputS5xD(20)(0);
  CNStageIntLLRInputS6xD(76)(0) <= VNStageIntLLROutputS5xD(20)(1);
  CNStageIntLLRInputS6xD(277)(0) <= VNStageIntLLROutputS5xD(20)(2);
  CNStageIntLLRInputS6xD(292)(0) <= VNStageIntLLROutputS5xD(20)(3);
  CNStageIntLLRInputS6xD(339)(0) <= VNStageIntLLROutputS5xD(20)(4);
  CNStageIntLLRInputS6xD(33)(0) <= VNStageIntLLROutputS5xD(21)(0);
  CNStageIntLLRInputS6xD(75)(0) <= VNStageIntLLROutputS5xD(21)(1);
  CNStageIntLLRInputS6xD(121)(0) <= VNStageIntLLROutputS5xD(21)(2);
  CNStageIntLLRInputS6xD(206)(0) <= VNStageIntLLROutputS5xD(21)(3);
  CNStageIntLLRInputS6xD(276)(0) <= VNStageIntLLROutputS5xD(21)(4);
  CNStageIntLLRInputS6xD(291)(0) <= VNStageIntLLROutputS5xD(21)(5);
  CNStageIntLLRInputS6xD(338)(0) <= VNStageIntLLROutputS5xD(21)(6);
  CNStageIntLLRInputS6xD(32)(0) <= VNStageIntLLROutputS5xD(22)(0);
  CNStageIntLLRInputS6xD(74)(0) <= VNStageIntLLROutputS5xD(22)(1);
  CNStageIntLLRInputS6xD(120)(0) <= VNStageIntLLROutputS5xD(22)(2);
  CNStageIntLLRInputS6xD(205)(0) <= VNStageIntLLROutputS5xD(22)(3);
  CNStageIntLLRInputS6xD(275)(0) <= VNStageIntLLROutputS5xD(22)(4);
  CNStageIntLLRInputS6xD(290)(0) <= VNStageIntLLROutputS5xD(22)(5);
  CNStageIntLLRInputS6xD(337)(0) <= VNStageIntLLROutputS5xD(22)(6);
  CNStageIntLLRInputS6xD(31)(0) <= VNStageIntLLROutputS5xD(23)(0);
  CNStageIntLLRInputS6xD(73)(0) <= VNStageIntLLROutputS5xD(23)(1);
  CNStageIntLLRInputS6xD(119)(0) <= VNStageIntLLROutputS5xD(23)(2);
  CNStageIntLLRInputS6xD(204)(0) <= VNStageIntLLROutputS5xD(23)(3);
  CNStageIntLLRInputS6xD(274)(0) <= VNStageIntLLROutputS5xD(23)(4);
  CNStageIntLLRInputS6xD(289)(0) <= VNStageIntLLROutputS5xD(23)(5);
  CNStageIntLLRInputS6xD(336)(0) <= VNStageIntLLROutputS5xD(23)(6);
  CNStageIntLLRInputS6xD(30)(0) <= VNStageIntLLROutputS5xD(24)(0);
  CNStageIntLLRInputS6xD(72)(0) <= VNStageIntLLROutputS5xD(24)(1);
  CNStageIntLLRInputS6xD(118)(0) <= VNStageIntLLROutputS5xD(24)(2);
  CNStageIntLLRInputS6xD(203)(0) <= VNStageIntLLROutputS5xD(24)(3);
  CNStageIntLLRInputS6xD(273)(0) <= VNStageIntLLROutputS5xD(24)(4);
  CNStageIntLLRInputS6xD(288)(0) <= VNStageIntLLROutputS5xD(24)(5);
  CNStageIntLLRInputS6xD(335)(0) <= VNStageIntLLROutputS5xD(24)(6);
  CNStageIntLLRInputS6xD(29)(0) <= VNStageIntLLROutputS5xD(25)(0);
  CNStageIntLLRInputS6xD(71)(0) <= VNStageIntLLROutputS5xD(25)(1);
  CNStageIntLLRInputS6xD(117)(0) <= VNStageIntLLROutputS5xD(25)(2);
  CNStageIntLLRInputS6xD(202)(0) <= VNStageIntLLROutputS5xD(25)(3);
  CNStageIntLLRInputS6xD(287)(0) <= VNStageIntLLROutputS5xD(25)(4);
  CNStageIntLLRInputS6xD(28)(0) <= VNStageIntLLROutputS5xD(26)(0);
  CNStageIntLLRInputS6xD(70)(0) <= VNStageIntLLROutputS5xD(26)(1);
  CNStageIntLLRInputS6xD(116)(0) <= VNStageIntLLROutputS5xD(26)(2);
  CNStageIntLLRInputS6xD(201)(0) <= VNStageIntLLROutputS5xD(26)(3);
  CNStageIntLLRInputS6xD(272)(0) <= VNStageIntLLROutputS5xD(26)(4);
  CNStageIntLLRInputS6xD(286)(0) <= VNStageIntLLROutputS5xD(26)(5);
  CNStageIntLLRInputS6xD(334)(0) <= VNStageIntLLROutputS5xD(26)(6);
  CNStageIntLLRInputS6xD(27)(0) <= VNStageIntLLROutputS5xD(27)(0);
  CNStageIntLLRInputS6xD(69)(0) <= VNStageIntLLROutputS5xD(27)(1);
  CNStageIntLLRInputS6xD(115)(0) <= VNStageIntLLROutputS5xD(27)(2);
  CNStageIntLLRInputS6xD(200)(0) <= VNStageIntLLROutputS5xD(27)(3);
  CNStageIntLLRInputS6xD(285)(0) <= VNStageIntLLROutputS5xD(27)(4);
  CNStageIntLLRInputS6xD(26)(0) <= VNStageIntLLROutputS5xD(28)(0);
  CNStageIntLLRInputS6xD(68)(0) <= VNStageIntLLROutputS5xD(28)(1);
  CNStageIntLLRInputS6xD(114)(0) <= VNStageIntLLROutputS5xD(28)(2);
  CNStageIntLLRInputS6xD(199)(0) <= VNStageIntLLROutputS5xD(28)(3);
  CNStageIntLLRInputS6xD(271)(0) <= VNStageIntLLROutputS5xD(28)(4);
  CNStageIntLLRInputS6xD(333)(0) <= VNStageIntLLROutputS5xD(28)(5);
  CNStageIntLLRInputS6xD(25)(0) <= VNStageIntLLROutputS5xD(29)(0);
  CNStageIntLLRInputS6xD(67)(0) <= VNStageIntLLROutputS5xD(29)(1);
  CNStageIntLLRInputS6xD(113)(0) <= VNStageIntLLROutputS5xD(29)(2);
  CNStageIntLLRInputS6xD(270)(0) <= VNStageIntLLROutputS5xD(29)(3);
  CNStageIntLLRInputS6xD(24)(0) <= VNStageIntLLROutputS5xD(30)(0);
  CNStageIntLLRInputS6xD(66)(0) <= VNStageIntLLROutputS5xD(30)(1);
  CNStageIntLLRInputS6xD(112)(0) <= VNStageIntLLROutputS5xD(30)(2);
  CNStageIntLLRInputS6xD(198)(0) <= VNStageIntLLROutputS5xD(30)(3);
  CNStageIntLLRInputS6xD(269)(0) <= VNStageIntLLROutputS5xD(30)(4);
  CNStageIntLLRInputS6xD(284)(0) <= VNStageIntLLROutputS5xD(30)(5);
  CNStageIntLLRInputS6xD(23)(0) <= VNStageIntLLROutputS5xD(31)(0);
  CNStageIntLLRInputS6xD(65)(0) <= VNStageIntLLROutputS5xD(31)(1);
  CNStageIntLLRInputS6xD(197)(0) <= VNStageIntLLROutputS5xD(31)(2);
  CNStageIntLLRInputS6xD(283)(0) <= VNStageIntLLROutputS5xD(31)(3);
  CNStageIntLLRInputS6xD(22)(0) <= VNStageIntLLROutputS5xD(32)(0);
  CNStageIntLLRInputS6xD(64)(0) <= VNStageIntLLROutputS5xD(32)(1);
  CNStageIntLLRInputS6xD(111)(0) <= VNStageIntLLROutputS5xD(32)(2);
  CNStageIntLLRInputS6xD(268)(0) <= VNStageIntLLROutputS5xD(32)(3);
  CNStageIntLLRInputS6xD(21)(0) <= VNStageIntLLROutputS5xD(33)(0);
  CNStageIntLLRInputS6xD(63)(0) <= VNStageIntLLROutputS5xD(33)(1);
  CNStageIntLLRInputS6xD(169)(0) <= VNStageIntLLROutputS5xD(33)(2);
  CNStageIntLLRInputS6xD(196)(0) <= VNStageIntLLROutputS5xD(33)(3);
  CNStageIntLLRInputS6xD(267)(0) <= VNStageIntLLROutputS5xD(33)(4);
  CNStageIntLLRInputS6xD(282)(0) <= VNStageIntLLROutputS5xD(33)(5);
  CNStageIntLLRInputS6xD(20)(0) <= VNStageIntLLROutputS5xD(34)(0);
  CNStageIntLLRInputS6xD(62)(0) <= VNStageIntLLROutputS5xD(34)(1);
  CNStageIntLLRInputS6xD(168)(0) <= VNStageIntLLROutputS5xD(34)(2);
  CNStageIntLLRInputS6xD(195)(0) <= VNStageIntLLROutputS5xD(34)(3);
  CNStageIntLLRInputS6xD(266)(0) <= VNStageIntLLROutputS5xD(34)(4);
  CNStageIntLLRInputS6xD(281)(0) <= VNStageIntLLROutputS5xD(34)(5);
  CNStageIntLLRInputS6xD(19)(0) <= VNStageIntLLROutputS5xD(35)(0);
  CNStageIntLLRInputS6xD(61)(0) <= VNStageIntLLROutputS5xD(35)(1);
  CNStageIntLLRInputS6xD(167)(0) <= VNStageIntLLROutputS5xD(35)(2);
  CNStageIntLLRInputS6xD(194)(0) <= VNStageIntLLROutputS5xD(35)(3);
  CNStageIntLLRInputS6xD(265)(0) <= VNStageIntLLROutputS5xD(35)(4);
  CNStageIntLLRInputS6xD(280)(0) <= VNStageIntLLROutputS5xD(35)(5);
  CNStageIntLLRInputS6xD(18)(0) <= VNStageIntLLROutputS5xD(36)(0);
  CNStageIntLLRInputS6xD(60)(0) <= VNStageIntLLROutputS5xD(36)(1);
  CNStageIntLLRInputS6xD(166)(0) <= VNStageIntLLROutputS5xD(36)(2);
  CNStageIntLLRInputS6xD(264)(0) <= VNStageIntLLROutputS5xD(36)(3);
  CNStageIntLLRInputS6xD(17)(0) <= VNStageIntLLROutputS5xD(37)(0);
  CNStageIntLLRInputS6xD(59)(0) <= VNStageIntLLROutputS5xD(37)(1);
  CNStageIntLLRInputS6xD(165)(0) <= VNStageIntLLROutputS5xD(37)(2);
  CNStageIntLLRInputS6xD(193)(0) <= VNStageIntLLROutputS5xD(37)(3);
  CNStageIntLLRInputS6xD(263)(0) <= VNStageIntLLROutputS5xD(37)(4);
  CNStageIntLLRInputS6xD(331)(0) <= VNStageIntLLROutputS5xD(37)(5);
  CNStageIntLLRInputS6xD(383)(0) <= VNStageIntLLROutputS5xD(37)(6);
  CNStageIntLLRInputS6xD(16)(0) <= VNStageIntLLROutputS5xD(38)(0);
  CNStageIntLLRInputS6xD(58)(0) <= VNStageIntLLROutputS5xD(38)(1);
  CNStageIntLLRInputS6xD(164)(0) <= VNStageIntLLROutputS5xD(38)(2);
  CNStageIntLLRInputS6xD(192)(0) <= VNStageIntLLROutputS5xD(38)(3);
  CNStageIntLLRInputS6xD(262)(0) <= VNStageIntLLROutputS5xD(38)(4);
  CNStageIntLLRInputS6xD(330)(0) <= VNStageIntLLROutputS5xD(38)(5);
  CNStageIntLLRInputS6xD(382)(0) <= VNStageIntLLROutputS5xD(38)(6);
  CNStageIntLLRInputS6xD(15)(0) <= VNStageIntLLROutputS5xD(39)(0);
  CNStageIntLLRInputS6xD(57)(0) <= VNStageIntLLROutputS5xD(39)(1);
  CNStageIntLLRInputS6xD(163)(0) <= VNStageIntLLROutputS5xD(39)(2);
  CNStageIntLLRInputS6xD(191)(0) <= VNStageIntLLROutputS5xD(39)(3);
  CNStageIntLLRInputS6xD(261)(0) <= VNStageIntLLROutputS5xD(39)(4);
  CNStageIntLLRInputS6xD(329)(0) <= VNStageIntLLROutputS5xD(39)(5);
  CNStageIntLLRInputS6xD(381)(0) <= VNStageIntLLROutputS5xD(39)(6);
  CNStageIntLLRInputS6xD(14)(0) <= VNStageIntLLROutputS5xD(40)(0);
  CNStageIntLLRInputS6xD(56)(0) <= VNStageIntLLROutputS5xD(40)(1);
  CNStageIntLLRInputS6xD(162)(0) <= VNStageIntLLROutputS5xD(40)(2);
  CNStageIntLLRInputS6xD(260)(0) <= VNStageIntLLROutputS5xD(40)(3);
  CNStageIntLLRInputS6xD(380)(0) <= VNStageIntLLROutputS5xD(40)(4);
  CNStageIntLLRInputS6xD(13)(0) <= VNStageIntLLROutputS5xD(41)(0);
  CNStageIntLLRInputS6xD(55)(0) <= VNStageIntLLROutputS5xD(41)(1);
  CNStageIntLLRInputS6xD(161)(0) <= VNStageIntLLROutputS5xD(41)(2);
  CNStageIntLLRInputS6xD(190)(0) <= VNStageIntLLROutputS5xD(41)(3);
  CNStageIntLLRInputS6xD(259)(0) <= VNStageIntLLROutputS5xD(41)(4);
  CNStageIntLLRInputS6xD(328)(0) <= VNStageIntLLROutputS5xD(41)(5);
  CNStageIntLLRInputS6xD(379)(0) <= VNStageIntLLROutputS5xD(41)(6);
  CNStageIntLLRInputS6xD(12)(0) <= VNStageIntLLROutputS5xD(42)(0);
  CNStageIntLLRInputS6xD(54)(0) <= VNStageIntLLROutputS5xD(42)(1);
  CNStageIntLLRInputS6xD(160)(0) <= VNStageIntLLROutputS5xD(42)(2);
  CNStageIntLLRInputS6xD(189)(0) <= VNStageIntLLROutputS5xD(42)(3);
  CNStageIntLLRInputS6xD(258)(0) <= VNStageIntLLROutputS5xD(42)(4);
  CNStageIntLLRInputS6xD(327)(0) <= VNStageIntLLROutputS5xD(42)(5);
  CNStageIntLLRInputS6xD(378)(0) <= VNStageIntLLROutputS5xD(42)(6);
  CNStageIntLLRInputS6xD(109)(0) <= VNStageIntLLROutputS5xD(43)(0);
  CNStageIntLLRInputS6xD(159)(0) <= VNStageIntLLROutputS5xD(43)(1);
  CNStageIntLLRInputS6xD(188)(0) <= VNStageIntLLROutputS5xD(43)(2);
  CNStageIntLLRInputS6xD(257)(0) <= VNStageIntLLROutputS5xD(43)(3);
  CNStageIntLLRInputS6xD(326)(0) <= VNStageIntLLROutputS5xD(43)(4);
  CNStageIntLLRInputS6xD(377)(0) <= VNStageIntLLROutputS5xD(43)(5);
  CNStageIntLLRInputS6xD(11)(0) <= VNStageIntLLROutputS5xD(44)(0);
  CNStageIntLLRInputS6xD(108)(0) <= VNStageIntLLROutputS5xD(44)(1);
  CNStageIntLLRInputS6xD(158)(0) <= VNStageIntLLROutputS5xD(44)(2);
  CNStageIntLLRInputS6xD(187)(0) <= VNStageIntLLROutputS5xD(44)(3);
  CNStageIntLLRInputS6xD(256)(0) <= VNStageIntLLROutputS5xD(44)(4);
  CNStageIntLLRInputS6xD(325)(0) <= VNStageIntLLROutputS5xD(44)(5);
  CNStageIntLLRInputS6xD(376)(0) <= VNStageIntLLROutputS5xD(44)(6);
  CNStageIntLLRInputS6xD(10)(0) <= VNStageIntLLROutputS5xD(45)(0);
  CNStageIntLLRInputS6xD(107)(0) <= VNStageIntLLROutputS5xD(45)(1);
  CNStageIntLLRInputS6xD(157)(0) <= VNStageIntLLROutputS5xD(45)(2);
  CNStageIntLLRInputS6xD(186)(0) <= VNStageIntLLROutputS5xD(45)(3);
  CNStageIntLLRInputS6xD(255)(0) <= VNStageIntLLROutputS5xD(45)(4);
  CNStageIntLLRInputS6xD(324)(0) <= VNStageIntLLROutputS5xD(45)(5);
  CNStageIntLLRInputS6xD(375)(0) <= VNStageIntLLROutputS5xD(45)(6);
  CNStageIntLLRInputS6xD(9)(0) <= VNStageIntLLROutputS5xD(46)(0);
  CNStageIntLLRInputS6xD(106)(0) <= VNStageIntLLROutputS5xD(46)(1);
  CNStageIntLLRInputS6xD(156)(0) <= VNStageIntLLROutputS5xD(46)(2);
  CNStageIntLLRInputS6xD(185)(0) <= VNStageIntLLROutputS5xD(46)(3);
  CNStageIntLLRInputS6xD(254)(0) <= VNStageIntLLROutputS5xD(46)(4);
  CNStageIntLLRInputS6xD(323)(0) <= VNStageIntLLROutputS5xD(46)(5);
  CNStageIntLLRInputS6xD(374)(0) <= VNStageIntLLROutputS5xD(46)(6);
  CNStageIntLLRInputS6xD(8)(0) <= VNStageIntLLROutputS5xD(47)(0);
  CNStageIntLLRInputS6xD(155)(0) <= VNStageIntLLROutputS5xD(47)(1);
  CNStageIntLLRInputS6xD(253)(0) <= VNStageIntLLROutputS5xD(47)(2);
  CNStageIntLLRInputS6xD(373)(0) <= VNStageIntLLROutputS5xD(47)(3);
  CNStageIntLLRInputS6xD(7)(0) <= VNStageIntLLROutputS5xD(48)(0);
  CNStageIntLLRInputS6xD(154)(0) <= VNStageIntLLROutputS5xD(48)(1);
  CNStageIntLLRInputS6xD(322)(0) <= VNStageIntLLROutputS5xD(48)(2);
  CNStageIntLLRInputS6xD(372)(0) <= VNStageIntLLROutputS5xD(48)(3);
  CNStageIntLLRInputS6xD(6)(0) <= VNStageIntLLROutputS5xD(49)(0);
  CNStageIntLLRInputS6xD(105)(0) <= VNStageIntLLROutputS5xD(49)(1);
  CNStageIntLLRInputS6xD(153)(0) <= VNStageIntLLROutputS5xD(49)(2);
  CNStageIntLLRInputS6xD(184)(0) <= VNStageIntLLROutputS5xD(49)(3);
  CNStageIntLLRInputS6xD(252)(0) <= VNStageIntLLROutputS5xD(49)(4);
  CNStageIntLLRInputS6xD(321)(0) <= VNStageIntLLROutputS5xD(49)(5);
  CNStageIntLLRInputS6xD(371)(0) <= VNStageIntLLROutputS5xD(49)(6);
  CNStageIntLLRInputS6xD(5)(0) <= VNStageIntLLROutputS5xD(50)(0);
  CNStageIntLLRInputS6xD(104)(0) <= VNStageIntLLROutputS5xD(50)(1);
  CNStageIntLLRInputS6xD(152)(0) <= VNStageIntLLROutputS5xD(50)(2);
  CNStageIntLLRInputS6xD(183)(0) <= VNStageIntLLROutputS5xD(50)(3);
  CNStageIntLLRInputS6xD(251)(0) <= VNStageIntLLROutputS5xD(50)(4);
  CNStageIntLLRInputS6xD(320)(0) <= VNStageIntLLROutputS5xD(50)(5);
  CNStageIntLLRInputS6xD(370)(0) <= VNStageIntLLROutputS5xD(50)(6);
  CNStageIntLLRInputS6xD(4)(0) <= VNStageIntLLROutputS5xD(51)(0);
  CNStageIntLLRInputS6xD(103)(0) <= VNStageIntLLROutputS5xD(51)(1);
  CNStageIntLLRInputS6xD(182)(0) <= VNStageIntLLROutputS5xD(51)(2);
  CNStageIntLLRInputS6xD(250)(0) <= VNStageIntLLROutputS5xD(51)(3);
  CNStageIntLLRInputS6xD(319)(0) <= VNStageIntLLROutputS5xD(51)(4);
  CNStageIntLLRInputS6xD(369)(0) <= VNStageIntLLROutputS5xD(51)(5);
  CNStageIntLLRInputS6xD(102)(0) <= VNStageIntLLROutputS5xD(52)(0);
  CNStageIntLLRInputS6xD(151)(0) <= VNStageIntLLROutputS5xD(52)(1);
  CNStageIntLLRInputS6xD(181)(0) <= VNStageIntLLROutputS5xD(52)(2);
  CNStageIntLLRInputS6xD(318)(0) <= VNStageIntLLROutputS5xD(52)(3);
  CNStageIntLLRInputS6xD(368)(0) <= VNStageIntLLROutputS5xD(52)(4);
  CNStageIntLLRInputS6xD(3)(0) <= VNStageIntLLROutputS5xD(53)(0);
  CNStageIntLLRInputS6xD(150)(0) <= VNStageIntLLROutputS5xD(53)(1);
  CNStageIntLLRInputS6xD(180)(0) <= VNStageIntLLROutputS5xD(53)(2);
  CNStageIntLLRInputS6xD(249)(0) <= VNStageIntLLROutputS5xD(53)(3);
  CNStageIntLLRInputS6xD(317)(0) <= VNStageIntLLROutputS5xD(53)(4);
  CNStageIntLLRInputS6xD(367)(0) <= VNStageIntLLROutputS5xD(53)(5);
  CNStageIntLLRInputS6xD(2)(0) <= VNStageIntLLROutputS5xD(54)(0);
  CNStageIntLLRInputS6xD(101)(0) <= VNStageIntLLROutputS5xD(54)(1);
  CNStageIntLLRInputS6xD(149)(0) <= VNStageIntLLROutputS5xD(54)(2);
  CNStageIntLLRInputS6xD(179)(0) <= VNStageIntLLROutputS5xD(54)(3);
  CNStageIntLLRInputS6xD(316)(0) <= VNStageIntLLROutputS5xD(54)(4);
  CNStageIntLLRInputS6xD(366)(0) <= VNStageIntLLROutputS5xD(54)(5);
  CNStageIntLLRInputS6xD(1)(0) <= VNStageIntLLROutputS5xD(55)(0);
  CNStageIntLLRInputS6xD(100)(0) <= VNStageIntLLROutputS5xD(55)(1);
  CNStageIntLLRInputS6xD(148)(0) <= VNStageIntLLROutputS5xD(55)(2);
  CNStageIntLLRInputS6xD(178)(0) <= VNStageIntLLROutputS5xD(55)(3);
  CNStageIntLLRInputS6xD(248)(0) <= VNStageIntLLROutputS5xD(55)(4);
  CNStageIntLLRInputS6xD(315)(0) <= VNStageIntLLROutputS5xD(55)(5);
  CNStageIntLLRInputS6xD(365)(0) <= VNStageIntLLROutputS5xD(55)(6);
  CNStageIntLLRInputS6xD(0)(0) <= VNStageIntLLROutputS5xD(56)(0);
  CNStageIntLLRInputS6xD(99)(0) <= VNStageIntLLROutputS5xD(56)(1);
  CNStageIntLLRInputS6xD(147)(0) <= VNStageIntLLROutputS5xD(56)(2);
  CNStageIntLLRInputS6xD(177)(0) <= VNStageIntLLROutputS5xD(56)(3);
  CNStageIntLLRInputS6xD(247)(0) <= VNStageIntLLROutputS5xD(56)(4);
  CNStageIntLLRInputS6xD(314)(0) <= VNStageIntLLROutputS5xD(56)(5);
  CNStageIntLLRInputS6xD(364)(0) <= VNStageIntLLROutputS5xD(56)(6);
  CNStageIntLLRInputS6xD(98)(0) <= VNStageIntLLROutputS5xD(57)(0);
  CNStageIntLLRInputS6xD(146)(0) <= VNStageIntLLROutputS5xD(57)(1);
  CNStageIntLLRInputS6xD(176)(0) <= VNStageIntLLROutputS5xD(57)(2);
  CNStageIntLLRInputS6xD(246)(0) <= VNStageIntLLROutputS5xD(57)(3);
  CNStageIntLLRInputS6xD(313)(0) <= VNStageIntLLROutputS5xD(57)(4);
  CNStageIntLLRInputS6xD(363)(0) <= VNStageIntLLROutputS5xD(57)(5);
  CNStageIntLLRInputS6xD(97)(0) <= VNStageIntLLROutputS5xD(58)(0);
  CNStageIntLLRInputS6xD(145)(0) <= VNStageIntLLROutputS5xD(58)(1);
  CNStageIntLLRInputS6xD(175)(0) <= VNStageIntLLROutputS5xD(58)(2);
  CNStageIntLLRInputS6xD(312)(0) <= VNStageIntLLROutputS5xD(58)(3);
  CNStageIntLLRInputS6xD(362)(0) <= VNStageIntLLROutputS5xD(58)(4);
  CNStageIntLLRInputS6xD(144)(0) <= VNStageIntLLROutputS5xD(59)(0);
  CNStageIntLLRInputS6xD(174)(0) <= VNStageIntLLROutputS5xD(59)(1);
  CNStageIntLLRInputS6xD(245)(0) <= VNStageIntLLROutputS5xD(59)(2);
  CNStageIntLLRInputS6xD(311)(0) <= VNStageIntLLROutputS5xD(59)(3);
  CNStageIntLLRInputS6xD(361)(0) <= VNStageIntLLROutputS5xD(59)(4);
  CNStageIntLLRInputS6xD(96)(0) <= VNStageIntLLROutputS5xD(60)(0);
  CNStageIntLLRInputS6xD(143)(0) <= VNStageIntLLROutputS5xD(60)(1);
  CNStageIntLLRInputS6xD(173)(0) <= VNStageIntLLROutputS5xD(60)(2);
  CNStageIntLLRInputS6xD(244)(0) <= VNStageIntLLROutputS5xD(60)(3);
  CNStageIntLLRInputS6xD(310)(0) <= VNStageIntLLROutputS5xD(60)(4);
  CNStageIntLLRInputS6xD(360)(0) <= VNStageIntLLROutputS5xD(60)(5);
  CNStageIntLLRInputS6xD(95)(0) <= VNStageIntLLROutputS5xD(61)(0);
  CNStageIntLLRInputS6xD(142)(0) <= VNStageIntLLROutputS5xD(61)(1);
  CNStageIntLLRInputS6xD(172)(0) <= VNStageIntLLROutputS5xD(61)(2);
  CNStageIntLLRInputS6xD(243)(0) <= VNStageIntLLROutputS5xD(61)(3);
  CNStageIntLLRInputS6xD(309)(0) <= VNStageIntLLROutputS5xD(61)(4);
  CNStageIntLLRInputS6xD(359)(0) <= VNStageIntLLROutputS5xD(61)(5);
  CNStageIntLLRInputS6xD(94)(0) <= VNStageIntLLROutputS5xD(62)(0);
  CNStageIntLLRInputS6xD(141)(0) <= VNStageIntLLROutputS5xD(62)(1);
  CNStageIntLLRInputS6xD(171)(0) <= VNStageIntLLROutputS5xD(62)(2);
  CNStageIntLLRInputS6xD(242)(0) <= VNStageIntLLROutputS5xD(62)(3);
  CNStageIntLLRInputS6xD(308)(0) <= VNStageIntLLROutputS5xD(62)(4);
  CNStageIntLLRInputS6xD(358)(0) <= VNStageIntLLROutputS5xD(62)(5);
  CNStageIntLLRInputS6xD(52)(0) <= VNStageIntLLROutputS5xD(63)(0);
  CNStageIntLLRInputS6xD(93)(0) <= VNStageIntLLROutputS5xD(63)(1);
  CNStageIntLLRInputS6xD(140)(0) <= VNStageIntLLROutputS5xD(63)(2);
  CNStageIntLLRInputS6xD(357)(0) <= VNStageIntLLROutputS5xD(63)(3);
  CNStageIntLLRInputS6xD(53)(1) <= VNStageIntLLROutputS5xD(64)(0);
  CNStageIntLLRInputS6xD(109)(1) <= VNStageIntLLROutputS5xD(64)(1);
  CNStageIntLLRInputS6xD(130)(1) <= VNStageIntLLROutputS5xD(64)(2);
  CNStageIntLLRInputS6xD(245)(1) <= VNStageIntLLROutputS5xD(64)(3);
  CNStageIntLLRInputS6xD(299)(1) <= VNStageIntLLROutputS5xD(64)(4);
  CNStageIntLLRInputS6xD(342)(1) <= VNStageIntLLROutputS5xD(64)(5);
  CNStageIntLLRInputS6xD(51)(1) <= VNStageIntLLROutputS5xD(65)(0);
  CNStageIntLLRInputS6xD(74)(1) <= VNStageIntLLROutputS5xD(65)(1);
  CNStageIntLLRInputS6xD(141)(1) <= VNStageIntLLROutputS5xD(65)(2);
  CNStageIntLLRInputS6xD(189)(1) <= VNStageIntLLROutputS5xD(65)(3);
  CNStageIntLLRInputS6xD(286)(1) <= VNStageIntLLROutputS5xD(65)(4);
  CNStageIntLLRInputS6xD(50)(1) <= VNStageIntLLROutputS5xD(66)(0);
  CNStageIntLLRInputS6xD(66)(1) <= VNStageIntLLROutputS5xD(66)(1);
  CNStageIntLLRInputS6xD(155)(1) <= VNStageIntLLROutputS5xD(66)(2);
  CNStageIntLLRInputS6xD(244)(1) <= VNStageIntLLROutputS5xD(66)(3);
  CNStageIntLLRInputS6xD(97)(1) <= VNStageIntLLROutputS5xD(67)(0);
  CNStageIntLLRInputS6xD(275)(1) <= VNStageIntLLROutputS5xD(67)(1);
  CNStageIntLLRInputS6xD(322)(1) <= VNStageIntLLROutputS5xD(67)(2);
  CNStageIntLLRInputS6xD(365)(1) <= VNStageIntLLROutputS5xD(67)(3);
  CNStageIntLLRInputS6xD(49)(1) <= VNStageIntLLROutputS5xD(68)(0);
  CNStageIntLLRInputS6xD(112)(1) <= VNStageIntLLROutputS5xD(68)(1);
  CNStageIntLLRInputS6xD(210)(1) <= VNStageIntLLROutputS5xD(68)(2);
  CNStageIntLLRInputS6xD(256)(1) <= VNStageIntLLROutputS5xD(68)(3);
  CNStageIntLLRInputS6xD(318)(1) <= VNStageIntLLROutputS5xD(68)(4);
  CNStageIntLLRInputS6xD(381)(1) <= VNStageIntLLROutputS5xD(68)(5);
  CNStageIntLLRInputS6xD(48)(1) <= VNStageIntLLROutputS5xD(69)(0);
  CNStageIntLLRInputS6xD(101)(1) <= VNStageIntLLROutputS5xD(69)(1);
  CNStageIntLLRInputS6xD(135)(1) <= VNStageIntLLROutputS5xD(69)(2);
  CNStageIntLLRInputS6xD(215)(1) <= VNStageIntLLROutputS5xD(69)(3);
  CNStageIntLLRInputS6xD(259)(1) <= VNStageIntLLROutputS5xD(69)(4);
  CNStageIntLLRInputS6xD(283)(1) <= VNStageIntLLROutputS5xD(69)(5);
  CNStageIntLLRInputS6xD(351)(1) <= VNStageIntLLROutputS5xD(69)(6);
  CNStageIntLLRInputS6xD(47)(1) <= VNStageIntLLROutputS5xD(70)(0);
  CNStageIntLLRInputS6xD(104)(1) <= VNStageIntLLROutputS5xD(70)(1);
  CNStageIntLLRInputS6xD(136)(1) <= VNStageIntLLROutputS5xD(70)(2);
  CNStageIntLLRInputS6xD(206)(1) <= VNStageIntLLROutputS5xD(70)(3);
  CNStageIntLLRInputS6xD(246)(1) <= VNStageIntLLROutputS5xD(70)(4);
  CNStageIntLLRInputS6xD(301)(1) <= VNStageIntLLROutputS5xD(70)(5);
  CNStageIntLLRInputS6xD(46)(1) <= VNStageIntLLROutputS5xD(71)(0);
  CNStageIntLLRInputS6xD(95)(1) <= VNStageIntLLROutputS5xD(71)(1);
  CNStageIntLLRInputS6xD(176)(1) <= VNStageIntLLROutputS5xD(71)(2);
  CNStageIntLLRInputS6xD(276)(1) <= VNStageIntLLROutputS5xD(71)(3);
  CNStageIntLLRInputS6xD(302)(1) <= VNStageIntLLROutputS5xD(71)(4);
  CNStageIntLLRInputS6xD(353)(1) <= VNStageIntLLROutputS5xD(71)(5);
  CNStageIntLLRInputS6xD(45)(1) <= VNStageIntLLROutputS5xD(72)(0);
  CNStageIntLLRInputS6xD(75)(1) <= VNStageIntLLROutputS5xD(72)(1);
  CNStageIntLLRInputS6xD(162)(1) <= VNStageIntLLROutputS5xD(72)(2);
  CNStageIntLLRInputS6xD(183)(1) <= VNStageIntLLROutputS5xD(72)(3);
  CNStageIntLLRInputS6xD(243)(1) <= VNStageIntLLROutputS5xD(72)(4);
  CNStageIntLLRInputS6xD(367)(1) <= VNStageIntLLROutputS5xD(72)(5);
  CNStageIntLLRInputS6xD(44)(1) <= VNStageIntLLROutputS5xD(73)(0);
  CNStageIntLLRInputS6xD(56)(1) <= VNStageIntLLROutputS5xD(73)(1);
  CNStageIntLLRInputS6xD(121)(1) <= VNStageIntLLROutputS5xD(73)(2);
  CNStageIntLLRInputS6xD(219)(1) <= VNStageIntLLROutputS5xD(73)(3);
  CNStageIntLLRInputS6xD(328)(1) <= VNStageIntLLROutputS5xD(73)(4);
  CNStageIntLLRInputS6xD(363)(1) <= VNStageIntLLROutputS5xD(73)(5);
  CNStageIntLLRInputS6xD(43)(1) <= VNStageIntLLROutputS5xD(74)(0);
  CNStageIntLLRInputS6xD(70)(1) <= VNStageIntLLROutputS5xD(74)(1);
  CNStageIntLLRInputS6xD(125)(1) <= VNStageIntLLROutputS5xD(74)(2);
  CNStageIntLLRInputS6xD(221)(1) <= VNStageIntLLROutputS5xD(74)(3);
  CNStageIntLLRInputS6xD(290)(1) <= VNStageIntLLROutputS5xD(74)(4);
  CNStageIntLLRInputS6xD(42)(1) <= VNStageIntLLROutputS5xD(75)(0);
  CNStageIntLLRInputS6xD(81)(1) <= VNStageIntLLROutputS5xD(75)(1);
  CNStageIntLLRInputS6xD(170)(1) <= VNStageIntLLROutputS5xD(75)(2);
  CNStageIntLLRInputS6xD(192)(1) <= VNStageIntLLROutputS5xD(75)(3);
  CNStageIntLLRInputS6xD(278)(1) <= VNStageIntLLROutputS5xD(75)(4);
  CNStageIntLLRInputS6xD(294)(1) <= VNStageIntLLROutputS5xD(75)(5);
  CNStageIntLLRInputS6xD(347)(1) <= VNStageIntLLROutputS5xD(75)(6);
  CNStageIntLLRInputS6xD(41)(1) <= VNStageIntLLROutputS5xD(76)(0);
  CNStageIntLLRInputS6xD(106)(1) <= VNStageIntLLROutputS5xD(76)(1);
  CNStageIntLLRInputS6xD(124)(1) <= VNStageIntLLROutputS5xD(76)(2);
  CNStageIntLLRInputS6xD(174)(1) <= VNStageIntLLROutputS5xD(76)(3);
  CNStageIntLLRInputS6xD(270)(1) <= VNStageIntLLROutputS5xD(76)(4);
  CNStageIntLLRInputS6xD(332)(1) <= VNStageIntLLROutputS5xD(76)(5);
  CNStageIntLLRInputS6xD(348)(1) <= VNStageIntLLROutputS5xD(76)(6);
  CNStageIntLLRInputS6xD(119)(1) <= VNStageIntLLROutputS5xD(77)(0);
  CNStageIntLLRInputS6xD(185)(1) <= VNStageIntLLROutputS5xD(77)(1);
  CNStageIntLLRInputS6xD(257)(1) <= VNStageIntLLROutputS5xD(77)(2);
  CNStageIntLLRInputS6xD(293)(1) <= VNStageIntLLROutputS5xD(77)(3);
  CNStageIntLLRInputS6xD(383)(1) <= VNStageIntLLROutputS5xD(77)(4);
  CNStageIntLLRInputS6xD(40)(1) <= VNStageIntLLROutputS5xD(78)(0);
  CNStageIntLLRInputS6xD(84)(1) <= VNStageIntLLROutputS5xD(78)(1);
  CNStageIntLLRInputS6xD(159)(1) <= VNStageIntLLROutputS5xD(78)(2);
  CNStageIntLLRInputS6xD(193)(1) <= VNStageIntLLROutputS5xD(78)(3);
  CNStageIntLLRInputS6xD(274)(1) <= VNStageIntLLROutputS5xD(78)(4);
  CNStageIntLLRInputS6xD(288)(1) <= VNStageIntLLROutputS5xD(78)(5);
  CNStageIntLLRInputS6xD(374)(1) <= VNStageIntLLROutputS5xD(78)(6);
  CNStageIntLLRInputS6xD(39)(1) <= VNStageIntLLROutputS5xD(79)(0);
  CNStageIntLLRInputS6xD(99)(1) <= VNStageIntLLROutputS5xD(79)(1);
  CNStageIntLLRInputS6xD(167)(1) <= VNStageIntLLROutputS5xD(79)(2);
  CNStageIntLLRInputS6xD(220)(1) <= VNStageIntLLROutputS5xD(79)(3);
  CNStageIntLLRInputS6xD(325)(1) <= VNStageIntLLROutputS5xD(79)(4);
  CNStageIntLLRInputS6xD(38)(1) <= VNStageIntLLROutputS5xD(80)(0);
  CNStageIntLLRInputS6xD(62)(1) <= VNStageIntLLROutputS5xD(80)(1);
  CNStageIntLLRInputS6xD(131)(1) <= VNStageIntLLROutputS5xD(80)(2);
  CNStageIntLLRInputS6xD(182)(1) <= VNStageIntLLROutputS5xD(80)(3);
  CNStageIntLLRInputS6xD(248)(1) <= VNStageIntLLROutputS5xD(80)(4);
  CNStageIntLLRInputS6xD(337)(1) <= VNStageIntLLROutputS5xD(80)(5);
  CNStageIntLLRInputS6xD(37)(1) <= VNStageIntLLROutputS5xD(81)(0);
  CNStageIntLLRInputS6xD(72)(1) <= VNStageIntLLROutputS5xD(81)(1);
  CNStageIntLLRInputS6xD(129)(1) <= VNStageIntLLROutputS5xD(81)(2);
  CNStageIntLLRInputS6xD(262)(1) <= VNStageIntLLROutputS5xD(81)(3);
  CNStageIntLLRInputS6xD(36)(1) <= VNStageIntLLROutputS5xD(82)(0);
  CNStageIntLLRInputS6xD(67)(1) <= VNStageIntLLROutputS5xD(82)(1);
  CNStageIntLLRInputS6xD(165)(1) <= VNStageIntLLROutputS5xD(82)(2);
  CNStageIntLLRInputS6xD(188)(1) <= VNStageIntLLROutputS5xD(82)(3);
  CNStageIntLLRInputS6xD(254)(1) <= VNStageIntLLROutputS5xD(82)(4);
  CNStageIntLLRInputS6xD(298)(1) <= VNStageIntLLROutputS5xD(82)(5);
  CNStageIntLLRInputS6xD(336)(1) <= VNStageIntLLROutputS5xD(82)(6);
  CNStageIntLLRInputS6xD(35)(1) <= VNStageIntLLROutputS5xD(83)(0);
  CNStageIntLLRInputS6xD(73)(1) <= VNStageIntLLROutputS5xD(83)(1);
  CNStageIntLLRInputS6xD(144)(1) <= VNStageIntLLROutputS5xD(83)(2);
  CNStageIntLLRInputS6xD(208)(1) <= VNStageIntLLROutputS5xD(83)(3);
  CNStageIntLLRInputS6xD(232)(1) <= VNStageIntLLROutputS5xD(83)(4);
  CNStageIntLLRInputS6xD(330)(1) <= VNStageIntLLROutputS5xD(83)(5);
  CNStageIntLLRInputS6xD(34)(1) <= VNStageIntLLROutputS5xD(84)(0);
  CNStageIntLLRInputS6xD(61)(1) <= VNStageIntLLROutputS5xD(84)(1);
  CNStageIntLLRInputS6xD(147)(1) <= VNStageIntLLROutputS5xD(84)(2);
  CNStageIntLLRInputS6xD(222)(1) <= VNStageIntLLROutputS5xD(84)(3);
  CNStageIntLLRInputS6xD(310)(1) <= VNStageIntLLROutputS5xD(84)(4);
  CNStageIntLLRInputS6xD(371)(1) <= VNStageIntLLROutputS5xD(84)(5);
  CNStageIntLLRInputS6xD(33)(1) <= VNStageIntLLROutputS5xD(85)(0);
  CNStageIntLLRInputS6xD(132)(1) <= VNStageIntLLROutputS5xD(85)(1);
  CNStageIntLLRInputS6xD(218)(1) <= VNStageIntLLROutputS5xD(85)(2);
  CNStageIntLLRInputS6xD(235)(1) <= VNStageIntLLROutputS5xD(85)(3);
  CNStageIntLLRInputS6xD(313)(1) <= VNStageIntLLROutputS5xD(85)(4);
  CNStageIntLLRInputS6xD(379)(1) <= VNStageIntLLROutputS5xD(85)(5);
  CNStageIntLLRInputS6xD(32)(1) <= VNStageIntLLROutputS5xD(86)(0);
  CNStageIntLLRInputS6xD(166)(1) <= VNStageIntLLROutputS5xD(86)(1);
  CNStageIntLLRInputS6xD(239)(1) <= VNStageIntLLROutputS5xD(86)(2);
  CNStageIntLLRInputS6xD(343)(1) <= VNStageIntLLROutputS5xD(86)(3);
  CNStageIntLLRInputS6xD(31)(1) <= VNStageIntLLROutputS5xD(87)(0);
  CNStageIntLLRInputS6xD(77)(1) <= VNStageIntLLROutputS5xD(87)(1);
  CNStageIntLLRInputS6xD(128)(1) <= VNStageIntLLROutputS5xD(87)(2);
  CNStageIntLLRInputS6xD(203)(1) <= VNStageIntLLROutputS5xD(87)(3);
  CNStageIntLLRInputS6xD(229)(1) <= VNStageIntLLROutputS5xD(87)(4);
  CNStageIntLLRInputS6xD(331)(1) <= VNStageIntLLROutputS5xD(87)(5);
  CNStageIntLLRInputS6xD(341)(1) <= VNStageIntLLROutputS5xD(87)(6);
  CNStageIntLLRInputS6xD(30)(1) <= VNStageIntLLROutputS5xD(88)(0);
  CNStageIntLLRInputS6xD(79)(1) <= VNStageIntLLROutputS5xD(88)(1);
  CNStageIntLLRInputS6xD(156)(1) <= VNStageIntLLROutputS5xD(88)(2);
  CNStageIntLLRInputS6xD(204)(1) <= VNStageIntLLROutputS5xD(88)(3);
  CNStageIntLLRInputS6xD(263)(1) <= VNStageIntLLROutputS5xD(88)(4);
  CNStageIntLLRInputS6xD(297)(1) <= VNStageIntLLROutputS5xD(88)(5);
  CNStageIntLLRInputS6xD(377)(1) <= VNStageIntLLROutputS5xD(88)(6);
  CNStageIntLLRInputS6xD(29)(1) <= VNStageIntLLROutputS5xD(89)(0);
  CNStageIntLLRInputS6xD(102)(1) <= VNStageIntLLROutputS5xD(89)(1);
  CNStageIntLLRInputS6xD(140)(1) <= VNStageIntLLROutputS5xD(89)(2);
  CNStageIntLLRInputS6xD(184)(1) <= VNStageIntLLROutputS5xD(89)(3);
  CNStageIntLLRInputS6xD(247)(1) <= VNStageIntLLROutputS5xD(89)(4);
  CNStageIntLLRInputS6xD(355)(1) <= VNStageIntLLROutputS5xD(89)(5);
  CNStageIntLLRInputS6xD(28)(1) <= VNStageIntLLROutputS5xD(90)(0);
  CNStageIntLLRInputS6xD(85)(1) <= VNStageIntLLROutputS5xD(90)(1);
  CNStageIntLLRInputS6xD(168)(1) <= VNStageIntLLROutputS5xD(90)(2);
  CNStageIntLLRInputS6xD(175)(1) <= VNStageIntLLROutputS5xD(90)(3);
  CNStageIntLLRInputS6xD(258)(1) <= VNStageIntLLROutputS5xD(90)(4);
  CNStageIntLLRInputS6xD(307)(1) <= VNStageIntLLROutputS5xD(90)(5);
  CNStageIntLLRInputS6xD(358)(1) <= VNStageIntLLROutputS5xD(90)(6);
  CNStageIntLLRInputS6xD(27)(1) <= VNStageIntLLROutputS5xD(91)(0);
  CNStageIntLLRInputS6xD(96)(1) <= VNStageIntLLROutputS5xD(91)(1);
  CNStageIntLLRInputS6xD(158)(1) <= VNStageIntLLROutputS5xD(91)(2);
  CNStageIntLLRInputS6xD(191)(1) <= VNStageIntLLROutputS5xD(91)(3);
  CNStageIntLLRInputS6xD(269)(1) <= VNStageIntLLROutputS5xD(91)(4);
  CNStageIntLLRInputS6xD(280)(1) <= VNStageIntLLROutputS5xD(91)(5);
  CNStageIntLLRInputS6xD(344)(1) <= VNStageIntLLROutputS5xD(91)(6);
  CNStageIntLLRInputS6xD(26)(1) <= VNStageIntLLROutputS5xD(92)(0);
  CNStageIntLLRInputS6xD(103)(1) <= VNStageIntLLROutputS5xD(92)(1);
  CNStageIntLLRInputS6xD(145)(1) <= VNStageIntLLROutputS5xD(92)(2);
  CNStageIntLLRInputS6xD(195)(1) <= VNStageIntLLROutputS5xD(92)(3);
  CNStageIntLLRInputS6xD(242)(1) <= VNStageIntLLROutputS5xD(92)(4);
  CNStageIntLLRInputS6xD(324)(1) <= VNStageIntLLROutputS5xD(92)(5);
  CNStageIntLLRInputS6xD(378)(1) <= VNStageIntLLROutputS5xD(92)(6);
  CNStageIntLLRInputS6xD(25)(1) <= VNStageIntLLROutputS5xD(93)(0);
  CNStageIntLLRInputS6xD(78)(1) <= VNStageIntLLROutputS5xD(93)(1);
  CNStageIntLLRInputS6xD(164)(1) <= VNStageIntLLROutputS5xD(93)(2);
  CNStageIntLLRInputS6xD(224)(1) <= VNStageIntLLROutputS5xD(93)(3);
  CNStageIntLLRInputS6xD(231)(1) <= VNStageIntLLROutputS5xD(93)(4);
  CNStageIntLLRInputS6xD(311)(1) <= VNStageIntLLROutputS5xD(93)(5);
  CNStageIntLLRInputS6xD(340)(1) <= VNStageIntLLROutputS5xD(93)(6);
  CNStageIntLLRInputS6xD(24)(1) <= VNStageIntLLROutputS5xD(94)(0);
  CNStageIntLLRInputS6xD(92)(1) <= VNStageIntLLROutputS5xD(94)(1);
  CNStageIntLLRInputS6xD(194)(1) <= VNStageIntLLROutputS5xD(94)(2);
  CNStageIntLLRInputS6xD(329)(1) <= VNStageIntLLROutputS5xD(94)(3);
  CNStageIntLLRInputS6xD(368)(1) <= VNStageIntLLROutputS5xD(94)(4);
  CNStageIntLLRInputS6xD(23)(1) <= VNStageIntLLROutputS5xD(95)(0);
  CNStageIntLLRInputS6xD(63)(1) <= VNStageIntLLROutputS5xD(95)(1);
  CNStageIntLLRInputS6xD(134)(1) <= VNStageIntLLROutputS5xD(95)(2);
  CNStageIntLLRInputS6xD(190)(1) <= VNStageIntLLROutputS5xD(95)(3);
  CNStageIntLLRInputS6xD(234)(1) <= VNStageIntLLROutputS5xD(95)(4);
  CNStageIntLLRInputS6xD(303)(1) <= VNStageIntLLROutputS5xD(95)(5);
  CNStageIntLLRInputS6xD(352)(1) <= VNStageIntLLROutputS5xD(95)(6);
  CNStageIntLLRInputS6xD(22)(1) <= VNStageIntLLROutputS5xD(96)(0);
  CNStageIntLLRInputS6xD(98)(1) <= VNStageIntLLROutputS5xD(96)(1);
  CNStageIntLLRInputS6xD(150)(1) <= VNStageIntLLROutputS5xD(96)(2);
  CNStageIntLLRInputS6xD(172)(1) <= VNStageIntLLROutputS5xD(96)(3);
  CNStageIntLLRInputS6xD(251)(1) <= VNStageIntLLROutputS5xD(96)(4);
  CNStageIntLLRInputS6xD(380)(1) <= VNStageIntLLROutputS5xD(96)(5);
  CNStageIntLLRInputS6xD(21)(1) <= VNStageIntLLROutputS5xD(97)(0);
  CNStageIntLLRInputS6xD(65)(1) <= VNStageIntLLROutputS5xD(97)(1);
  CNStageIntLLRInputS6xD(142)(1) <= VNStageIntLLROutputS5xD(97)(2);
  CNStageIntLLRInputS6xD(180)(1) <= VNStageIntLLROutputS5xD(97)(3);
  CNStageIntLLRInputS6xD(260)(1) <= VNStageIntLLROutputS5xD(97)(4);
  CNStageIntLLRInputS6xD(316)(1) <= VNStageIntLLROutputS5xD(97)(5);
  CNStageIntLLRInputS6xD(370)(1) <= VNStageIntLLROutputS5xD(97)(6);
  CNStageIntLLRInputS6xD(20)(1) <= VNStageIntLLROutputS5xD(98)(0);
  CNStageIntLLRInputS6xD(116)(1) <= VNStageIntLLROutputS5xD(98)(1);
  CNStageIntLLRInputS6xD(199)(1) <= VNStageIntLLROutputS5xD(98)(2);
  CNStageIntLLRInputS6xD(255)(1) <= VNStageIntLLROutputS5xD(98)(3);
  CNStageIntLLRInputS6xD(308)(1) <= VNStageIntLLROutputS5xD(98)(4);
  CNStageIntLLRInputS6xD(356)(1) <= VNStageIntLLROutputS5xD(98)(5);
  CNStageIntLLRInputS6xD(19)(1) <= VNStageIntLLROutputS5xD(99)(0);
  CNStageIntLLRInputS6xD(76)(1) <= VNStageIntLLROutputS5xD(99)(1);
  CNStageIntLLRInputS6xD(126)(1) <= VNStageIntLLROutputS5xD(99)(2);
  CNStageIntLLRInputS6xD(198)(1) <= VNStageIntLLROutputS5xD(99)(3);
  CNStageIntLLRInputS6xD(261)(1) <= VNStageIntLLROutputS5xD(99)(4);
  CNStageIntLLRInputS6xD(285)(1) <= VNStageIntLLROutputS5xD(99)(5);
  CNStageIntLLRInputS6xD(376)(1) <= VNStageIntLLROutputS5xD(99)(6);
  CNStageIntLLRInputS6xD(18)(1) <= VNStageIntLLROutputS5xD(100)(0);
  CNStageIntLLRInputS6xD(94)(1) <= VNStageIntLLROutputS5xD(100)(1);
  CNStageIntLLRInputS6xD(120)(1) <= VNStageIntLLROutputS5xD(100)(2);
  CNStageIntLLRInputS6xD(178)(1) <= VNStageIntLLROutputS5xD(100)(3);
  CNStageIntLLRInputS6xD(250)(1) <= VNStageIntLLROutputS5xD(100)(4);
  CNStageIntLLRInputS6xD(295)(1) <= VNStageIntLLROutputS5xD(100)(5);
  CNStageIntLLRInputS6xD(349)(1) <= VNStageIntLLROutputS5xD(100)(6);
  CNStageIntLLRInputS6xD(17)(1) <= VNStageIntLLROutputS5xD(101)(0);
  CNStageIntLLRInputS6xD(58)(1) <= VNStageIntLLROutputS5xD(101)(1);
  CNStageIntLLRInputS6xD(123)(1) <= VNStageIntLLROutputS5xD(101)(2);
  CNStageIntLLRInputS6xD(211)(1) <= VNStageIntLLROutputS5xD(101)(3);
  CNStageIntLLRInputS6xD(273)(1) <= VNStageIntLLROutputS5xD(101)(4);
  CNStageIntLLRInputS6xD(289)(1) <= VNStageIntLLROutputS5xD(101)(5);
  CNStageIntLLRInputS6xD(346)(1) <= VNStageIntLLROutputS5xD(101)(6);
  CNStageIntLLRInputS6xD(16)(1) <= VNStageIntLLROutputS5xD(102)(0);
  CNStageIntLLRInputS6xD(59)(1) <= VNStageIntLLROutputS5xD(102)(1);
  CNStageIntLLRInputS6xD(113)(1) <= VNStageIntLLROutputS5xD(102)(2);
  CNStageIntLLRInputS6xD(214)(1) <= VNStageIntLLROutputS5xD(102)(3);
  CNStageIntLLRInputS6xD(226)(1) <= VNStageIntLLROutputS5xD(102)(4);
  CNStageIntLLRInputS6xD(361)(1) <= VNStageIntLLROutputS5xD(102)(5);
  CNStageIntLLRInputS6xD(15)(1) <= VNStageIntLLROutputS5xD(103)(0);
  CNStageIntLLRInputS6xD(93)(1) <= VNStageIntLLROutputS5xD(103)(1);
  CNStageIntLLRInputS6xD(151)(1) <= VNStageIntLLROutputS5xD(103)(2);
  CNStageIntLLRInputS6xD(200)(1) <= VNStageIntLLROutputS5xD(103)(3);
  CNStageIntLLRInputS6xD(265)(1) <= VNStageIntLLROutputS5xD(103)(4);
  CNStageIntLLRInputS6xD(284)(1) <= VNStageIntLLROutputS5xD(103)(5);
  CNStageIntLLRInputS6xD(354)(1) <= VNStageIntLLROutputS5xD(103)(6);
  CNStageIntLLRInputS6xD(14)(1) <= VNStageIntLLROutputS5xD(104)(0);
  CNStageIntLLRInputS6xD(86)(1) <= VNStageIntLLROutputS5xD(104)(1);
  CNStageIntLLRInputS6xD(133)(1) <= VNStageIntLLROutputS5xD(104)(2);
  CNStageIntLLRInputS6xD(179)(1) <= VNStageIntLLROutputS5xD(104)(3);
  CNStageIntLLRInputS6xD(267)(1) <= VNStageIntLLROutputS5xD(104)(4);
  CNStageIntLLRInputS6xD(317)(1) <= VNStageIntLLROutputS5xD(104)(5);
  CNStageIntLLRInputS6xD(13)(1) <= VNStageIntLLROutputS5xD(105)(0);
  CNStageIntLLRInputS6xD(146)(1) <= VNStageIntLLROutputS5xD(105)(1);
  CNStageIntLLRInputS6xD(197)(1) <= VNStageIntLLROutputS5xD(105)(2);
  CNStageIntLLRInputS6xD(237)(1) <= VNStageIntLLROutputS5xD(105)(3);
  CNStageIntLLRInputS6xD(300)(1) <= VNStageIntLLROutputS5xD(105)(4);
  CNStageIntLLRInputS6xD(338)(1) <= VNStageIntLLROutputS5xD(105)(5);
  CNStageIntLLRInputS6xD(12)(1) <= VNStageIntLLROutputS5xD(106)(0);
  CNStageIntLLRInputS6xD(157)(1) <= VNStageIntLLROutputS5xD(106)(1);
  CNStageIntLLRInputS6xD(223)(1) <= VNStageIntLLROutputS5xD(106)(2);
  CNStageIntLLRInputS6xD(272)(1) <= VNStageIntLLROutputS5xD(106)(3);
  CNStageIntLLRInputS6xD(312)(1) <= VNStageIntLLROutputS5xD(106)(4);
  CNStageIntLLRInputS6xD(333)(1) <= VNStageIntLLROutputS5xD(106)(5);
  CNStageIntLLRInputS6xD(110)(1) <= VNStageIntLLROutputS5xD(107)(0);
  CNStageIntLLRInputS6xD(127)(1) <= VNStageIntLLROutputS5xD(107)(1);
  CNStageIntLLRInputS6xD(207)(1) <= VNStageIntLLROutputS5xD(107)(2);
  CNStageIntLLRInputS6xD(230)(1) <= VNStageIntLLROutputS5xD(107)(3);
  CNStageIntLLRInputS6xD(323)(1) <= VNStageIntLLROutputS5xD(107)(4);
  CNStageIntLLRInputS6xD(335)(1) <= VNStageIntLLROutputS5xD(107)(5);
  CNStageIntLLRInputS6xD(11)(1) <= VNStageIntLLROutputS5xD(108)(0);
  CNStageIntLLRInputS6xD(105)(1) <= VNStageIntLLROutputS5xD(108)(1);
  CNStageIntLLRInputS6xD(115)(1) <= VNStageIntLLROutputS5xD(108)(2);
  CNStageIntLLRInputS6xD(181)(1) <= VNStageIntLLROutputS5xD(108)(3);
  CNStageIntLLRInputS6xD(238)(1) <= VNStageIntLLROutputS5xD(108)(4);
  CNStageIntLLRInputS6xD(296)(1) <= VNStageIntLLROutputS5xD(108)(5);
  CNStageIntLLRInputS6xD(10)(1) <= VNStageIntLLROutputS5xD(109)(0);
  CNStageIntLLRInputS6xD(100)(1) <= VNStageIntLLROutputS5xD(109)(1);
  CNStageIntLLRInputS6xD(160)(1) <= VNStageIntLLROutputS5xD(109)(2);
  CNStageIntLLRInputS6xD(171)(1) <= VNStageIntLLROutputS5xD(109)(3);
  CNStageIntLLRInputS6xD(266)(1) <= VNStageIntLLROutputS5xD(109)(4);
  CNStageIntLLRInputS6xD(362)(1) <= VNStageIntLLROutputS5xD(109)(5);
  CNStageIntLLRInputS6xD(9)(1) <= VNStageIntLLROutputS5xD(110)(0);
  CNStageIntLLRInputS6xD(83)(1) <= VNStageIntLLROutputS5xD(110)(1);
  CNStageIntLLRInputS6xD(118)(1) <= VNStageIntLLROutputS5xD(110)(2);
  CNStageIntLLRInputS6xD(212)(1) <= VNStageIntLLROutputS5xD(110)(3);
  CNStageIntLLRInputS6xD(225)(1) <= VNStageIntLLROutputS5xD(110)(4);
  CNStageIntLLRInputS6xD(326)(1) <= VNStageIntLLROutputS5xD(110)(5);
  CNStageIntLLRInputS6xD(345)(1) <= VNStageIntLLROutputS5xD(110)(6);
  CNStageIntLLRInputS6xD(8)(1) <= VNStageIntLLROutputS5xD(111)(0);
  CNStageIntLLRInputS6xD(90)(1) <= VNStageIntLLROutputS5xD(111)(1);
  CNStageIntLLRInputS6xD(138)(1) <= VNStageIntLLROutputS5xD(111)(2);
  CNStageIntLLRInputS6xD(177)(1) <= VNStageIntLLROutputS5xD(111)(3);
  CNStageIntLLRInputS6xD(252)(1) <= VNStageIntLLROutputS5xD(111)(4);
  CNStageIntLLRInputS6xD(287)(1) <= VNStageIntLLROutputS5xD(111)(5);
  CNStageIntLLRInputS6xD(357)(1) <= VNStageIntLLROutputS5xD(111)(6);
  CNStageIntLLRInputS6xD(7)(1) <= VNStageIntLLROutputS5xD(112)(0);
  CNStageIntLLRInputS6xD(54)(1) <= VNStageIntLLROutputS5xD(112)(1);
  CNStageIntLLRInputS6xD(148)(1) <= VNStageIntLLROutputS5xD(112)(2);
  CNStageIntLLRInputS6xD(205)(1) <= VNStageIntLLROutputS5xD(112)(3);
  CNStageIntLLRInputS6xD(233)(1) <= VNStageIntLLROutputS5xD(112)(4);
  CNStageIntLLRInputS6xD(305)(1) <= VNStageIntLLROutputS5xD(112)(5);
  CNStageIntLLRInputS6xD(369)(1) <= VNStageIntLLROutputS5xD(112)(6);
  CNStageIntLLRInputS6xD(6)(1) <= VNStageIntLLROutputS5xD(113)(0);
  CNStageIntLLRInputS6xD(108)(1) <= VNStageIntLLROutputS5xD(113)(1);
  CNStageIntLLRInputS6xD(143)(1) <= VNStageIntLLROutputS5xD(113)(2);
  CNStageIntLLRInputS6xD(202)(1) <= VNStageIntLLROutputS5xD(113)(3);
  CNStageIntLLRInputS6xD(253)(1) <= VNStageIntLLROutputS5xD(113)(4);
  CNStageIntLLRInputS6xD(314)(1) <= VNStageIntLLROutputS5xD(113)(5);
  CNStageIntLLRInputS6xD(339)(1) <= VNStageIntLLROutputS5xD(113)(6);
  CNStageIntLLRInputS6xD(5)(1) <= VNStageIntLLROutputS5xD(114)(0);
  CNStageIntLLRInputS6xD(88)(1) <= VNStageIntLLROutputS5xD(114)(1);
  CNStageIntLLRInputS6xD(149)(1) <= VNStageIntLLROutputS5xD(114)(2);
  CNStageIntLLRInputS6xD(216)(1) <= VNStageIntLLROutputS5xD(114)(3);
  CNStageIntLLRInputS6xD(268)(1) <= VNStageIntLLROutputS5xD(114)(4);
  CNStageIntLLRInputS6xD(309)(1) <= VNStageIntLLROutputS5xD(114)(5);
  CNStageIntLLRInputS6xD(4)(1) <= VNStageIntLLROutputS5xD(115)(0);
  CNStageIntLLRInputS6xD(68)(1) <= VNStageIntLLROutputS5xD(115)(1);
  CNStageIntLLRInputS6xD(137)(1) <= VNStageIntLLROutputS5xD(115)(2);
  CNStageIntLLRInputS6xD(209)(1) <= VNStageIntLLROutputS5xD(115)(3);
  CNStageIntLLRInputS6xD(264)(1) <= VNStageIntLLROutputS5xD(115)(4);
  CNStageIntLLRInputS6xD(315)(1) <= VNStageIntLLROutputS5xD(115)(5);
  CNStageIntLLRInputS6xD(372)(1) <= VNStageIntLLROutputS5xD(115)(6);
  CNStageIntLLRInputS6xD(71)(1) <= VNStageIntLLROutputS5xD(116)(0);
  CNStageIntLLRInputS6xD(163)(1) <= VNStageIntLLROutputS5xD(116)(1);
  CNStageIntLLRInputS6xD(187)(1) <= VNStageIntLLROutputS5xD(116)(2);
  CNStageIntLLRInputS6xD(228)(1) <= VNStageIntLLROutputS5xD(116)(3);
  CNStageIntLLRInputS6xD(304)(1) <= VNStageIntLLROutputS5xD(116)(4);
  CNStageIntLLRInputS6xD(3)(1) <= VNStageIntLLROutputS5xD(117)(0);
  CNStageIntLLRInputS6xD(55)(1) <= VNStageIntLLROutputS5xD(117)(1);
  CNStageIntLLRInputS6xD(111)(1) <= VNStageIntLLROutputS5xD(117)(2);
  CNStageIntLLRInputS6xD(196)(1) <= VNStageIntLLROutputS5xD(117)(3);
  CNStageIntLLRInputS6xD(2)(1) <= VNStageIntLLROutputS5xD(118)(0);
  CNStageIntLLRInputS6xD(89)(1) <= VNStageIntLLROutputS5xD(118)(1);
  CNStageIntLLRInputS6xD(152)(1) <= VNStageIntLLROutputS5xD(118)(2);
  CNStageIntLLRInputS6xD(249)(1) <= VNStageIntLLROutputS5xD(118)(3);
  CNStageIntLLRInputS6xD(282)(1) <= VNStageIntLLROutputS5xD(118)(4);
  CNStageIntLLRInputS6xD(359)(1) <= VNStageIntLLROutputS5xD(118)(5);
  CNStageIntLLRInputS6xD(1)(1) <= VNStageIntLLROutputS5xD(119)(0);
  CNStageIntLLRInputS6xD(107)(1) <= VNStageIntLLROutputS5xD(119)(1);
  CNStageIntLLRInputS6xD(154)(1) <= VNStageIntLLROutputS5xD(119)(2);
  CNStageIntLLRInputS6xD(227)(1) <= VNStageIntLLROutputS5xD(119)(3);
  CNStageIntLLRInputS6xD(319)(1) <= VNStageIntLLROutputS5xD(119)(4);
  CNStageIntLLRInputS6xD(0)(1) <= VNStageIntLLROutputS5xD(120)(0);
  CNStageIntLLRInputS6xD(80)(1) <= VNStageIntLLROutputS5xD(120)(1);
  CNStageIntLLRInputS6xD(321)(1) <= VNStageIntLLROutputS5xD(120)(2);
  CNStageIntLLRInputS6xD(360)(1) <= VNStageIntLLROutputS5xD(120)(3);
  CNStageIntLLRInputS6xD(64)(1) <= VNStageIntLLROutputS5xD(121)(0);
  CNStageIntLLRInputS6xD(161)(1) <= VNStageIntLLROutputS5xD(121)(1);
  CNStageIntLLRInputS6xD(217)(1) <= VNStageIntLLROutputS5xD(121)(2);
  CNStageIntLLRInputS6xD(236)(1) <= VNStageIntLLROutputS5xD(121)(3);
  CNStageIntLLRInputS6xD(291)(1) <= VNStageIntLLROutputS5xD(121)(4);
  CNStageIntLLRInputS6xD(350)(1) <= VNStageIntLLROutputS5xD(121)(5);
  CNStageIntLLRInputS6xD(91)(1) <= VNStageIntLLROutputS5xD(122)(0);
  CNStageIntLLRInputS6xD(114)(1) <= VNStageIntLLROutputS5xD(122)(1);
  CNStageIntLLRInputS6xD(201)(1) <= VNStageIntLLROutputS5xD(122)(2);
  CNStageIntLLRInputS6xD(241)(1) <= VNStageIntLLROutputS5xD(122)(3);
  CNStageIntLLRInputS6xD(327)(1) <= VNStageIntLLROutputS5xD(122)(4);
  CNStageIntLLRInputS6xD(375)(1) <= VNStageIntLLROutputS5xD(122)(5);
  CNStageIntLLRInputS6xD(82)(1) <= VNStageIntLLROutputS5xD(123)(0);
  CNStageIntLLRInputS6xD(122)(1) <= VNStageIntLLROutputS5xD(123)(1);
  CNStageIntLLRInputS6xD(213)(1) <= VNStageIntLLROutputS5xD(123)(2);
  CNStageIntLLRInputS6xD(279)(1) <= VNStageIntLLROutputS5xD(123)(3);
  CNStageIntLLRInputS6xD(382)(1) <= VNStageIntLLROutputS5xD(123)(4);
  CNStageIntLLRInputS6xD(69)(1) <= VNStageIntLLROutputS5xD(124)(0);
  CNStageIntLLRInputS6xD(153)(1) <= VNStageIntLLROutputS5xD(124)(1);
  CNStageIntLLRInputS6xD(240)(1) <= VNStageIntLLROutputS5xD(124)(2);
  CNStageIntLLRInputS6xD(292)(1) <= VNStageIntLLROutputS5xD(124)(3);
  CNStageIntLLRInputS6xD(364)(1) <= VNStageIntLLROutputS5xD(124)(4);
  CNStageIntLLRInputS6xD(87)(1) <= VNStageIntLLROutputS5xD(125)(0);
  CNStageIntLLRInputS6xD(169)(1) <= VNStageIntLLROutputS5xD(125)(1);
  CNStageIntLLRInputS6xD(320)(1) <= VNStageIntLLROutputS5xD(125)(2);
  CNStageIntLLRInputS6xD(366)(1) <= VNStageIntLLROutputS5xD(125)(3);
  CNStageIntLLRInputS6xD(60)(1) <= VNStageIntLLROutputS5xD(126)(0);
  CNStageIntLLRInputS6xD(139)(1) <= VNStageIntLLROutputS5xD(126)(1);
  CNStageIntLLRInputS6xD(186)(1) <= VNStageIntLLROutputS5xD(126)(2);
  CNStageIntLLRInputS6xD(271)(1) <= VNStageIntLLROutputS5xD(126)(3);
  CNStageIntLLRInputS6xD(281)(1) <= VNStageIntLLROutputS5xD(126)(4);
  CNStageIntLLRInputS6xD(334)(1) <= VNStageIntLLROutputS5xD(126)(5);
  CNStageIntLLRInputS6xD(52)(1) <= VNStageIntLLROutputS5xD(127)(0);
  CNStageIntLLRInputS6xD(57)(1) <= VNStageIntLLROutputS5xD(127)(1);
  CNStageIntLLRInputS6xD(117)(1) <= VNStageIntLLROutputS5xD(127)(2);
  CNStageIntLLRInputS6xD(173)(1) <= VNStageIntLLROutputS5xD(127)(3);
  CNStageIntLLRInputS6xD(277)(1) <= VNStageIntLLROutputS5xD(127)(4);
  CNStageIntLLRInputS6xD(306)(1) <= VNStageIntLLROutputS5xD(127)(5);
  CNStageIntLLRInputS6xD(373)(1) <= VNStageIntLLROutputS5xD(127)(6);
  CNStageIntLLRInputS6xD(53)(2) <= VNStageIntLLROutputS5xD(128)(0);
  CNStageIntLLRInputS6xD(108)(2) <= VNStageIntLLROutputS5xD(128)(1);
  CNStageIntLLRInputS6xD(129)(2) <= VNStageIntLLROutputS5xD(128)(2);
  CNStageIntLLRInputS6xD(198)(2) <= VNStageIntLLROutputS5xD(128)(3);
  CNStageIntLLRInputS6xD(244)(2) <= VNStageIntLLROutputS5xD(128)(4);
  CNStageIntLLRInputS6xD(298)(2) <= VNStageIntLLROutputS5xD(128)(5);
  CNStageIntLLRInputS6xD(341)(2) <= VNStageIntLLROutputS5xD(128)(6);
  CNStageIntLLRInputS6xD(51)(2) <= VNStageIntLLROutputS5xD(129)(0);
  CNStageIntLLRInputS6xD(56)(2) <= VNStageIntLLROutputS5xD(129)(1);
  CNStageIntLLRInputS6xD(116)(2) <= VNStageIntLLROutputS5xD(129)(2);
  CNStageIntLLRInputS6xD(172)(2) <= VNStageIntLLROutputS5xD(129)(3);
  CNStageIntLLRInputS6xD(276)(2) <= VNStageIntLLROutputS5xD(129)(4);
  CNStageIntLLRInputS6xD(305)(2) <= VNStageIntLLROutputS5xD(129)(5);
  CNStageIntLLRInputS6xD(372)(2) <= VNStageIntLLROutputS5xD(129)(6);
  CNStageIntLLRInputS6xD(50)(2) <= VNStageIntLLROutputS5xD(130)(0);
  CNStageIntLLRInputS6xD(73)(2) <= VNStageIntLLROutputS5xD(130)(1);
  CNStageIntLLRInputS6xD(140)(2) <= VNStageIntLLROutputS5xD(130)(2);
  CNStageIntLLRInputS6xD(188)(2) <= VNStageIntLLROutputS5xD(130)(3);
  CNStageIntLLRInputS6xD(245)(2) <= VNStageIntLLROutputS5xD(130)(4);
  CNStageIntLLRInputS6xD(285)(2) <= VNStageIntLLROutputS5xD(130)(5);
  CNStageIntLLRInputS6xD(65)(2) <= VNStageIntLLROutputS5xD(131)(0);
  CNStageIntLLRInputS6xD(154)(2) <= VNStageIntLLROutputS5xD(131)(1);
  CNStageIntLLRInputS6xD(206)(2) <= VNStageIntLLROutputS5xD(131)(2);
  CNStageIntLLRInputS6xD(243)(2) <= VNStageIntLLROutputS5xD(131)(3);
  CNStageIntLLRInputS6xD(307)(2) <= VNStageIntLLROutputS5xD(131)(4);
  CNStageIntLLRInputS6xD(334)(2) <= VNStageIntLLROutputS5xD(131)(5);
  CNStageIntLLRInputS6xD(49)(2) <= VNStageIntLLROutputS5xD(132)(0);
  CNStageIntLLRInputS6xD(151)(2) <= VNStageIntLLROutputS5xD(132)(1);
  CNStageIntLLRInputS6xD(214)(2) <= VNStageIntLLROutputS5xD(132)(2);
  CNStageIntLLRInputS6xD(274)(2) <= VNStageIntLLROutputS5xD(132)(3);
  CNStageIntLLRInputS6xD(321)(2) <= VNStageIntLLROutputS5xD(132)(4);
  CNStageIntLLRInputS6xD(364)(2) <= VNStageIntLLROutputS5xD(132)(5);
  CNStageIntLLRInputS6xD(48)(2) <= VNStageIntLLROutputS5xD(133)(0);
  CNStageIntLLRInputS6xD(209)(2) <= VNStageIntLLROutputS5xD(133)(1);
  CNStageIntLLRInputS6xD(255)(2) <= VNStageIntLLROutputS5xD(133)(2);
  CNStageIntLLRInputS6xD(317)(2) <= VNStageIntLLROutputS5xD(133)(3);
  CNStageIntLLRInputS6xD(380)(2) <= VNStageIntLLROutputS5xD(133)(4);
  CNStageIntLLRInputS6xD(47)(2) <= VNStageIntLLROutputS5xD(134)(0);
  CNStageIntLLRInputS6xD(100)(2) <= VNStageIntLLROutputS5xD(134)(1);
  CNStageIntLLRInputS6xD(134)(2) <= VNStageIntLLROutputS5xD(134)(2);
  CNStageIntLLRInputS6xD(258)(2) <= VNStageIntLLROutputS5xD(134)(3);
  CNStageIntLLRInputS6xD(46)(2) <= VNStageIntLLROutputS5xD(135)(0);
  CNStageIntLLRInputS6xD(103)(2) <= VNStageIntLLROutputS5xD(135)(1);
  CNStageIntLLRInputS6xD(135)(2) <= VNStageIntLLROutputS5xD(135)(2);
  CNStageIntLLRInputS6xD(205)(2) <= VNStageIntLLROutputS5xD(135)(3);
  CNStageIntLLRInputS6xD(45)(2) <= VNStageIntLLROutputS5xD(136)(0);
  CNStageIntLLRInputS6xD(94)(2) <= VNStageIntLLROutputS5xD(136)(1);
  CNStageIntLLRInputS6xD(111)(2) <= VNStageIntLLROutputS5xD(136)(2);
  CNStageIntLLRInputS6xD(175)(2) <= VNStageIntLLROutputS5xD(136)(3);
  CNStageIntLLRInputS6xD(275)(2) <= VNStageIntLLROutputS5xD(136)(4);
  CNStageIntLLRInputS6xD(301)(2) <= VNStageIntLLROutputS5xD(136)(5);
  CNStageIntLLRInputS6xD(352)(2) <= VNStageIntLLROutputS5xD(136)(6);
  CNStageIntLLRInputS6xD(44)(2) <= VNStageIntLLROutputS5xD(137)(0);
  CNStageIntLLRInputS6xD(74)(2) <= VNStageIntLLROutputS5xD(137)(1);
  CNStageIntLLRInputS6xD(161)(2) <= VNStageIntLLROutputS5xD(137)(2);
  CNStageIntLLRInputS6xD(182)(2) <= VNStageIntLLROutputS5xD(137)(3);
  CNStageIntLLRInputS6xD(242)(2) <= VNStageIntLLROutputS5xD(137)(4);
  CNStageIntLLRInputS6xD(282)(2) <= VNStageIntLLROutputS5xD(137)(5);
  CNStageIntLLRInputS6xD(366)(2) <= VNStageIntLLROutputS5xD(137)(6);
  CNStageIntLLRInputS6xD(43)(2) <= VNStageIntLLROutputS5xD(138)(0);
  CNStageIntLLRInputS6xD(55)(2) <= VNStageIntLLROutputS5xD(138)(1);
  CNStageIntLLRInputS6xD(120)(2) <= VNStageIntLLROutputS5xD(138)(2);
  CNStageIntLLRInputS6xD(218)(2) <= VNStageIntLLROutputS5xD(138)(3);
  CNStageIntLLRInputS6xD(268)(2) <= VNStageIntLLROutputS5xD(138)(4);
  CNStageIntLLRInputS6xD(327)(2) <= VNStageIntLLROutputS5xD(138)(5);
  CNStageIntLLRInputS6xD(362)(2) <= VNStageIntLLROutputS5xD(138)(6);
  CNStageIntLLRInputS6xD(42)(2) <= VNStageIntLLROutputS5xD(139)(0);
  CNStageIntLLRInputS6xD(69)(2) <= VNStageIntLLROutputS5xD(139)(1);
  CNStageIntLLRInputS6xD(124)(2) <= VNStageIntLLROutputS5xD(139)(2);
  CNStageIntLLRInputS6xD(220)(2) <= VNStageIntLLROutputS5xD(139)(3);
  CNStageIntLLRInputS6xD(252)(2) <= VNStageIntLLROutputS5xD(139)(4);
  CNStageIntLLRInputS6xD(289)(2) <= VNStageIntLLROutputS5xD(139)(5);
  CNStageIntLLRInputS6xD(383)(2) <= VNStageIntLLROutputS5xD(139)(6);
  CNStageIntLLRInputS6xD(41)(2) <= VNStageIntLLROutputS5xD(140)(0);
  CNStageIntLLRInputS6xD(80)(2) <= VNStageIntLLROutputS5xD(140)(1);
  CNStageIntLLRInputS6xD(170)(2) <= VNStageIntLLROutputS5xD(140)(2);
  CNStageIntLLRInputS6xD(191)(2) <= VNStageIntLLROutputS5xD(140)(3);
  CNStageIntLLRInputS6xD(277)(2) <= VNStageIntLLROutputS5xD(140)(4);
  CNStageIntLLRInputS6xD(293)(2) <= VNStageIntLLROutputS5xD(140)(5);
  CNStageIntLLRInputS6xD(346)(2) <= VNStageIntLLROutputS5xD(140)(6);
  CNStageIntLLRInputS6xD(123)(2) <= VNStageIntLLROutputS5xD(141)(0);
  CNStageIntLLRInputS6xD(173)(2) <= VNStageIntLLROutputS5xD(141)(1);
  CNStageIntLLRInputS6xD(269)(2) <= VNStageIntLLROutputS5xD(141)(2);
  CNStageIntLLRInputS6xD(332)(2) <= VNStageIntLLROutputS5xD(141)(3);
  CNStageIntLLRInputS6xD(347)(2) <= VNStageIntLLROutputS5xD(141)(4);
  CNStageIntLLRInputS6xD(40)(2) <= VNStageIntLLROutputS5xD(142)(0);
  CNStageIntLLRInputS6xD(96)(2) <= VNStageIntLLROutputS5xD(142)(1);
  CNStageIntLLRInputS6xD(118)(2) <= VNStageIntLLROutputS5xD(142)(2);
  CNStageIntLLRInputS6xD(256)(2) <= VNStageIntLLROutputS5xD(142)(3);
  CNStageIntLLRInputS6xD(382)(2) <= VNStageIntLLROutputS5xD(142)(4);
  CNStageIntLLRInputS6xD(39)(2) <= VNStageIntLLROutputS5xD(143)(0);
  CNStageIntLLRInputS6xD(83)(2) <= VNStageIntLLROutputS5xD(143)(1);
  CNStageIntLLRInputS6xD(158)(2) <= VNStageIntLLROutputS5xD(143)(2);
  CNStageIntLLRInputS6xD(192)(2) <= VNStageIntLLROutputS5xD(143)(3);
  CNStageIntLLRInputS6xD(273)(2) <= VNStageIntLLROutputS5xD(143)(4);
  CNStageIntLLRInputS6xD(287)(2) <= VNStageIntLLROutputS5xD(143)(5);
  CNStageIntLLRInputS6xD(373)(2) <= VNStageIntLLROutputS5xD(143)(6);
  CNStageIntLLRInputS6xD(38)(2) <= VNStageIntLLROutputS5xD(144)(0);
  CNStageIntLLRInputS6xD(98)(2) <= VNStageIntLLROutputS5xD(144)(1);
  CNStageIntLLRInputS6xD(166)(2) <= VNStageIntLLROutputS5xD(144)(2);
  CNStageIntLLRInputS6xD(219)(2) <= VNStageIntLLROutputS5xD(144)(3);
  CNStageIntLLRInputS6xD(249)(2) <= VNStageIntLLROutputS5xD(144)(4);
  CNStageIntLLRInputS6xD(324)(2) <= VNStageIntLLROutputS5xD(144)(5);
  CNStageIntLLRInputS6xD(333)(2) <= VNStageIntLLROutputS5xD(144)(6);
  CNStageIntLLRInputS6xD(37)(2) <= VNStageIntLLROutputS5xD(145)(0);
  CNStageIntLLRInputS6xD(61)(2) <= VNStageIntLLROutputS5xD(145)(1);
  CNStageIntLLRInputS6xD(130)(2) <= VNStageIntLLROutputS5xD(145)(2);
  CNStageIntLLRInputS6xD(181)(2) <= VNStageIntLLROutputS5xD(145)(3);
  CNStageIntLLRInputS6xD(247)(2) <= VNStageIntLLROutputS5xD(145)(4);
  CNStageIntLLRInputS6xD(331)(2) <= VNStageIntLLROutputS5xD(145)(5);
  CNStageIntLLRInputS6xD(336)(2) <= VNStageIntLLROutputS5xD(145)(6);
  CNStageIntLLRInputS6xD(36)(2) <= VNStageIntLLROutputS5xD(146)(0);
  CNStageIntLLRInputS6xD(71)(2) <= VNStageIntLLROutputS5xD(146)(1);
  CNStageIntLLRInputS6xD(128)(2) <= VNStageIntLLROutputS5xD(146)(2);
  CNStageIntLLRInputS6xD(261)(2) <= VNStageIntLLROutputS5xD(146)(3);
  CNStageIntLLRInputS6xD(299)(2) <= VNStageIntLLROutputS5xD(146)(4);
  CNStageIntLLRInputS6xD(35)(2) <= VNStageIntLLROutputS5xD(147)(0);
  CNStageIntLLRInputS6xD(66)(2) <= VNStageIntLLROutputS5xD(147)(1);
  CNStageIntLLRInputS6xD(164)(2) <= VNStageIntLLROutputS5xD(147)(2);
  CNStageIntLLRInputS6xD(187)(2) <= VNStageIntLLROutputS5xD(147)(3);
  CNStageIntLLRInputS6xD(253)(2) <= VNStageIntLLROutputS5xD(147)(4);
  CNStageIntLLRInputS6xD(297)(2) <= VNStageIntLLROutputS5xD(147)(5);
  CNStageIntLLRInputS6xD(335)(2) <= VNStageIntLLROutputS5xD(147)(6);
  CNStageIntLLRInputS6xD(34)(2) <= VNStageIntLLROutputS5xD(148)(0);
  CNStageIntLLRInputS6xD(72)(2) <= VNStageIntLLROutputS5xD(148)(1);
  CNStageIntLLRInputS6xD(143)(2) <= VNStageIntLLROutputS5xD(148)(2);
  CNStageIntLLRInputS6xD(207)(2) <= VNStageIntLLROutputS5xD(148)(3);
  CNStageIntLLRInputS6xD(231)(2) <= VNStageIntLLROutputS5xD(148)(4);
  CNStageIntLLRInputS6xD(329)(2) <= VNStageIntLLROutputS5xD(148)(5);
  CNStageIntLLRInputS6xD(33)(2) <= VNStageIntLLROutputS5xD(149)(0);
  CNStageIntLLRInputS6xD(60)(2) <= VNStageIntLLROutputS5xD(149)(1);
  CNStageIntLLRInputS6xD(146)(2) <= VNStageIntLLROutputS5xD(149)(2);
  CNStageIntLLRInputS6xD(221)(2) <= VNStageIntLLROutputS5xD(149)(3);
  CNStageIntLLRInputS6xD(241)(2) <= VNStageIntLLROutputS5xD(149)(4);
  CNStageIntLLRInputS6xD(309)(2) <= VNStageIntLLROutputS5xD(149)(5);
  CNStageIntLLRInputS6xD(370)(2) <= VNStageIntLLROutputS5xD(149)(6);
  CNStageIntLLRInputS6xD(32)(2) <= VNStageIntLLROutputS5xD(150)(0);
  CNStageIntLLRInputS6xD(86)(2) <= VNStageIntLLROutputS5xD(150)(1);
  CNStageIntLLRInputS6xD(131)(2) <= VNStageIntLLROutputS5xD(150)(2);
  CNStageIntLLRInputS6xD(217)(2) <= VNStageIntLLROutputS5xD(150)(3);
  CNStageIntLLRInputS6xD(312)(2) <= VNStageIntLLROutputS5xD(150)(4);
  CNStageIntLLRInputS6xD(378)(2) <= VNStageIntLLROutputS5xD(150)(5);
  CNStageIntLLRInputS6xD(31)(2) <= VNStageIntLLROutputS5xD(151)(0);
  CNStageIntLLRInputS6xD(92)(2) <= VNStageIntLLROutputS5xD(151)(1);
  CNStageIntLLRInputS6xD(165)(2) <= VNStageIntLLROutputS5xD(151)(2);
  CNStageIntLLRInputS6xD(184)(2) <= VNStageIntLLROutputS5xD(151)(3);
  CNStageIntLLRInputS6xD(238)(2) <= VNStageIntLLROutputS5xD(151)(4);
  CNStageIntLLRInputS6xD(342)(2) <= VNStageIntLLROutputS5xD(151)(5);
  CNStageIntLLRInputS6xD(30)(2) <= VNStageIntLLROutputS5xD(152)(0);
  CNStageIntLLRInputS6xD(76)(2) <= VNStageIntLLROutputS5xD(152)(1);
  CNStageIntLLRInputS6xD(127)(2) <= VNStageIntLLROutputS5xD(152)(2);
  CNStageIntLLRInputS6xD(202)(2) <= VNStageIntLLROutputS5xD(152)(3);
  CNStageIntLLRInputS6xD(228)(2) <= VNStageIntLLROutputS5xD(152)(4);
  CNStageIntLLRInputS6xD(330)(2) <= VNStageIntLLROutputS5xD(152)(5);
  CNStageIntLLRInputS6xD(340)(2) <= VNStageIntLLROutputS5xD(152)(6);
  CNStageIntLLRInputS6xD(29)(2) <= VNStageIntLLROutputS5xD(153)(0);
  CNStageIntLLRInputS6xD(78)(2) <= VNStageIntLLROutputS5xD(153)(1);
  CNStageIntLLRInputS6xD(155)(2) <= VNStageIntLLROutputS5xD(153)(2);
  CNStageIntLLRInputS6xD(203)(2) <= VNStageIntLLROutputS5xD(153)(3);
  CNStageIntLLRInputS6xD(262)(2) <= VNStageIntLLROutputS5xD(153)(4);
  CNStageIntLLRInputS6xD(296)(2) <= VNStageIntLLROutputS5xD(153)(5);
  CNStageIntLLRInputS6xD(376)(2) <= VNStageIntLLROutputS5xD(153)(6);
  CNStageIntLLRInputS6xD(28)(2) <= VNStageIntLLROutputS5xD(154)(0);
  CNStageIntLLRInputS6xD(139)(2) <= VNStageIntLLROutputS5xD(154)(1);
  CNStageIntLLRInputS6xD(183)(2) <= VNStageIntLLROutputS5xD(154)(2);
  CNStageIntLLRInputS6xD(246)(2) <= VNStageIntLLROutputS5xD(154)(3);
  CNStageIntLLRInputS6xD(322)(2) <= VNStageIntLLROutputS5xD(154)(4);
  CNStageIntLLRInputS6xD(27)(2) <= VNStageIntLLROutputS5xD(155)(0);
  CNStageIntLLRInputS6xD(84)(2) <= VNStageIntLLROutputS5xD(155)(1);
  CNStageIntLLRInputS6xD(167)(2) <= VNStageIntLLROutputS5xD(155)(2);
  CNStageIntLLRInputS6xD(174)(2) <= VNStageIntLLROutputS5xD(155)(3);
  CNStageIntLLRInputS6xD(257)(2) <= VNStageIntLLROutputS5xD(155)(4);
  CNStageIntLLRInputS6xD(306)(2) <= VNStageIntLLROutputS5xD(155)(5);
  CNStageIntLLRInputS6xD(357)(2) <= VNStageIntLLROutputS5xD(155)(6);
  CNStageIntLLRInputS6xD(26)(2) <= VNStageIntLLROutputS5xD(156)(0);
  CNStageIntLLRInputS6xD(95)(2) <= VNStageIntLLROutputS5xD(156)(1);
  CNStageIntLLRInputS6xD(157)(2) <= VNStageIntLLROutputS5xD(156)(2);
  CNStageIntLLRInputS6xD(343)(2) <= VNStageIntLLROutputS5xD(156)(3);
  CNStageIntLLRInputS6xD(25)(2) <= VNStageIntLLROutputS5xD(157)(0);
  CNStageIntLLRInputS6xD(102)(2) <= VNStageIntLLROutputS5xD(157)(1);
  CNStageIntLLRInputS6xD(144)(2) <= VNStageIntLLROutputS5xD(157)(2);
  CNStageIntLLRInputS6xD(194)(2) <= VNStageIntLLROutputS5xD(157)(3);
  CNStageIntLLRInputS6xD(323)(2) <= VNStageIntLLROutputS5xD(157)(4);
  CNStageIntLLRInputS6xD(377)(2) <= VNStageIntLLROutputS5xD(157)(5);
  CNStageIntLLRInputS6xD(24)(2) <= VNStageIntLLROutputS5xD(158)(0);
  CNStageIntLLRInputS6xD(77)(2) <= VNStageIntLLROutputS5xD(158)(1);
  CNStageIntLLRInputS6xD(163)(2) <= VNStageIntLLROutputS5xD(158)(2);
  CNStageIntLLRInputS6xD(224)(2) <= VNStageIntLLROutputS5xD(158)(3);
  CNStageIntLLRInputS6xD(230)(2) <= VNStageIntLLROutputS5xD(158)(4);
  CNStageIntLLRInputS6xD(310)(2) <= VNStageIntLLROutputS5xD(158)(5);
  CNStageIntLLRInputS6xD(339)(2) <= VNStageIntLLROutputS5xD(158)(6);
  CNStageIntLLRInputS6xD(23)(2) <= VNStageIntLLROutputS5xD(159)(0);
  CNStageIntLLRInputS6xD(91)(2) <= VNStageIntLLROutputS5xD(159)(1);
  CNStageIntLLRInputS6xD(136)(2) <= VNStageIntLLROutputS5xD(159)(2);
  CNStageIntLLRInputS6xD(271)(2) <= VNStageIntLLROutputS5xD(159)(3);
  CNStageIntLLRInputS6xD(367)(2) <= VNStageIntLLROutputS5xD(159)(4);
  CNStageIntLLRInputS6xD(22)(2) <= VNStageIntLLROutputS5xD(160)(0);
  CNStageIntLLRInputS6xD(62)(2) <= VNStageIntLLROutputS5xD(160)(1);
  CNStageIntLLRInputS6xD(133)(2) <= VNStageIntLLROutputS5xD(160)(2);
  CNStageIntLLRInputS6xD(189)(2) <= VNStageIntLLROutputS5xD(160)(3);
  CNStageIntLLRInputS6xD(233)(2) <= VNStageIntLLROutputS5xD(160)(4);
  CNStageIntLLRInputS6xD(302)(2) <= VNStageIntLLROutputS5xD(160)(5);
  CNStageIntLLRInputS6xD(351)(2) <= VNStageIntLLROutputS5xD(160)(6);
  CNStageIntLLRInputS6xD(21)(2) <= VNStageIntLLROutputS5xD(161)(0);
  CNStageIntLLRInputS6xD(97)(2) <= VNStageIntLLROutputS5xD(161)(1);
  CNStageIntLLRInputS6xD(149)(2) <= VNStageIntLLROutputS5xD(161)(2);
  CNStageIntLLRInputS6xD(171)(2) <= VNStageIntLLROutputS5xD(161)(3);
  CNStageIntLLRInputS6xD(250)(2) <= VNStageIntLLROutputS5xD(161)(4);
  CNStageIntLLRInputS6xD(300)(2) <= VNStageIntLLROutputS5xD(161)(5);
  CNStageIntLLRInputS6xD(379)(2) <= VNStageIntLLROutputS5xD(161)(6);
  CNStageIntLLRInputS6xD(20)(2) <= VNStageIntLLROutputS5xD(162)(0);
  CNStageIntLLRInputS6xD(64)(2) <= VNStageIntLLROutputS5xD(162)(1);
  CNStageIntLLRInputS6xD(141)(2) <= VNStageIntLLROutputS5xD(162)(2);
  CNStageIntLLRInputS6xD(179)(2) <= VNStageIntLLROutputS5xD(162)(3);
  CNStageIntLLRInputS6xD(259)(2) <= VNStageIntLLROutputS5xD(162)(4);
  CNStageIntLLRInputS6xD(315)(2) <= VNStageIntLLROutputS5xD(162)(5);
  CNStageIntLLRInputS6xD(369)(2) <= VNStageIntLLROutputS5xD(162)(6);
  CNStageIntLLRInputS6xD(19)(2) <= VNStageIntLLROutputS5xD(163)(0);
  CNStageIntLLRInputS6xD(79)(2) <= VNStageIntLLROutputS5xD(163)(1);
  CNStageIntLLRInputS6xD(115)(2) <= VNStageIntLLROutputS5xD(163)(2);
  CNStageIntLLRInputS6xD(254)(2) <= VNStageIntLLROutputS5xD(163)(3);
  CNStageIntLLRInputS6xD(355)(2) <= VNStageIntLLROutputS5xD(163)(4);
  CNStageIntLLRInputS6xD(18)(2) <= VNStageIntLLROutputS5xD(164)(0);
  CNStageIntLLRInputS6xD(75)(2) <= VNStageIntLLROutputS5xD(164)(1);
  CNStageIntLLRInputS6xD(125)(2) <= VNStageIntLLROutputS5xD(164)(2);
  CNStageIntLLRInputS6xD(197)(2) <= VNStageIntLLROutputS5xD(164)(3);
  CNStageIntLLRInputS6xD(260)(2) <= VNStageIntLLROutputS5xD(164)(4);
  CNStageIntLLRInputS6xD(375)(2) <= VNStageIntLLROutputS5xD(164)(5);
  CNStageIntLLRInputS6xD(17)(2) <= VNStageIntLLROutputS5xD(165)(0);
  CNStageIntLLRInputS6xD(93)(2) <= VNStageIntLLROutputS5xD(165)(1);
  CNStageIntLLRInputS6xD(119)(2) <= VNStageIntLLROutputS5xD(165)(2);
  CNStageIntLLRInputS6xD(177)(2) <= VNStageIntLLROutputS5xD(165)(3);
  CNStageIntLLRInputS6xD(294)(2) <= VNStageIntLLROutputS5xD(165)(4);
  CNStageIntLLRInputS6xD(348)(2) <= VNStageIntLLROutputS5xD(165)(5);
  CNStageIntLLRInputS6xD(16)(2) <= VNStageIntLLROutputS5xD(166)(0);
  CNStageIntLLRInputS6xD(57)(2) <= VNStageIntLLROutputS5xD(166)(1);
  CNStageIntLLRInputS6xD(122)(2) <= VNStageIntLLROutputS5xD(166)(2);
  CNStageIntLLRInputS6xD(210)(2) <= VNStageIntLLROutputS5xD(166)(3);
  CNStageIntLLRInputS6xD(288)(2) <= VNStageIntLLROutputS5xD(166)(4);
  CNStageIntLLRInputS6xD(345)(2) <= VNStageIntLLROutputS5xD(166)(5);
  CNStageIntLLRInputS6xD(15)(2) <= VNStageIntLLROutputS5xD(167)(0);
  CNStageIntLLRInputS6xD(58)(2) <= VNStageIntLLROutputS5xD(167)(1);
  CNStageIntLLRInputS6xD(112)(2) <= VNStageIntLLROutputS5xD(167)(2);
  CNStageIntLLRInputS6xD(213)(2) <= VNStageIntLLROutputS5xD(167)(3);
  CNStageIntLLRInputS6xD(225)(2) <= VNStageIntLLROutputS5xD(167)(4);
  CNStageIntLLRInputS6xD(292)(2) <= VNStageIntLLROutputS5xD(167)(5);
  CNStageIntLLRInputS6xD(360)(2) <= VNStageIntLLROutputS5xD(167)(6);
  CNStageIntLLRInputS6xD(14)(2) <= VNStageIntLLROutputS5xD(168)(0);
  CNStageIntLLRInputS6xD(150)(2) <= VNStageIntLLROutputS5xD(168)(1);
  CNStageIntLLRInputS6xD(199)(2) <= VNStageIntLLROutputS5xD(168)(2);
  CNStageIntLLRInputS6xD(264)(2) <= VNStageIntLLROutputS5xD(168)(3);
  CNStageIntLLRInputS6xD(283)(2) <= VNStageIntLLROutputS5xD(168)(4);
  CNStageIntLLRInputS6xD(353)(2) <= VNStageIntLLROutputS5xD(168)(5);
  CNStageIntLLRInputS6xD(13)(2) <= VNStageIntLLROutputS5xD(169)(0);
  CNStageIntLLRInputS6xD(85)(2) <= VNStageIntLLROutputS5xD(169)(1);
  CNStageIntLLRInputS6xD(132)(2) <= VNStageIntLLROutputS5xD(169)(2);
  CNStageIntLLRInputS6xD(178)(2) <= VNStageIntLLROutputS5xD(169)(3);
  CNStageIntLLRInputS6xD(266)(2) <= VNStageIntLLROutputS5xD(169)(4);
  CNStageIntLLRInputS6xD(316)(2) <= VNStageIntLLROutputS5xD(169)(5);
  CNStageIntLLRInputS6xD(12)(2) <= VNStageIntLLROutputS5xD(170)(0);
  CNStageIntLLRInputS6xD(101)(2) <= VNStageIntLLROutputS5xD(170)(1);
  CNStageIntLLRInputS6xD(145)(2) <= VNStageIntLLROutputS5xD(170)(2);
  CNStageIntLLRInputS6xD(236)(2) <= VNStageIntLLROutputS5xD(170)(3);
  CNStageIntLLRInputS6xD(337)(2) <= VNStageIntLLROutputS5xD(170)(4);
  CNStageIntLLRInputS6xD(105)(2) <= VNStageIntLLROutputS5xD(171)(0);
  CNStageIntLLRInputS6xD(156)(2) <= VNStageIntLLROutputS5xD(171)(1);
  CNStageIntLLRInputS6xD(222)(2) <= VNStageIntLLROutputS5xD(171)(2);
  CNStageIntLLRInputS6xD(311)(2) <= VNStageIntLLROutputS5xD(171)(3);
  CNStageIntLLRInputS6xD(11)(2) <= VNStageIntLLROutputS5xD(172)(0);
  CNStageIntLLRInputS6xD(110)(2) <= VNStageIntLLROutputS5xD(172)(1);
  CNStageIntLLRInputS6xD(126)(2) <= VNStageIntLLROutputS5xD(172)(2);
  CNStageIntLLRInputS6xD(229)(2) <= VNStageIntLLROutputS5xD(172)(3);
  CNStageIntLLRInputS6xD(10)(2) <= VNStageIntLLROutputS5xD(173)(0);
  CNStageIntLLRInputS6xD(104)(2) <= VNStageIntLLROutputS5xD(173)(1);
  CNStageIntLLRInputS6xD(114)(2) <= VNStageIntLLROutputS5xD(173)(2);
  CNStageIntLLRInputS6xD(180)(2) <= VNStageIntLLROutputS5xD(173)(3);
  CNStageIntLLRInputS6xD(237)(2) <= VNStageIntLLROutputS5xD(173)(4);
  CNStageIntLLRInputS6xD(295)(2) <= VNStageIntLLROutputS5xD(173)(5);
  CNStageIntLLRInputS6xD(9)(2) <= VNStageIntLLROutputS5xD(174)(0);
  CNStageIntLLRInputS6xD(99)(2) <= VNStageIntLLROutputS5xD(174)(1);
  CNStageIntLLRInputS6xD(159)(2) <= VNStageIntLLROutputS5xD(174)(2);
  CNStageIntLLRInputS6xD(265)(2) <= VNStageIntLLROutputS5xD(174)(3);
  CNStageIntLLRInputS6xD(361)(2) <= VNStageIntLLROutputS5xD(174)(4);
  CNStageIntLLRInputS6xD(8)(2) <= VNStageIntLLROutputS5xD(175)(0);
  CNStageIntLLRInputS6xD(82)(2) <= VNStageIntLLROutputS5xD(175)(1);
  CNStageIntLLRInputS6xD(117)(2) <= VNStageIntLLROutputS5xD(175)(2);
  CNStageIntLLRInputS6xD(211)(2) <= VNStageIntLLROutputS5xD(175)(3);
  CNStageIntLLRInputS6xD(278)(2) <= VNStageIntLLROutputS5xD(175)(4);
  CNStageIntLLRInputS6xD(325)(2) <= VNStageIntLLROutputS5xD(175)(5);
  CNStageIntLLRInputS6xD(344)(2) <= VNStageIntLLROutputS5xD(175)(6);
  CNStageIntLLRInputS6xD(7)(2) <= VNStageIntLLROutputS5xD(176)(0);
  CNStageIntLLRInputS6xD(89)(2) <= VNStageIntLLROutputS5xD(176)(1);
  CNStageIntLLRInputS6xD(137)(2) <= VNStageIntLLROutputS5xD(176)(2);
  CNStageIntLLRInputS6xD(176)(2) <= VNStageIntLLROutputS5xD(176)(3);
  CNStageIntLLRInputS6xD(251)(2) <= VNStageIntLLROutputS5xD(176)(4);
  CNStageIntLLRInputS6xD(286)(2) <= VNStageIntLLROutputS5xD(176)(5);
  CNStageIntLLRInputS6xD(356)(2) <= VNStageIntLLROutputS5xD(176)(6);
  CNStageIntLLRInputS6xD(6)(2) <= VNStageIntLLROutputS5xD(177)(0);
  CNStageIntLLRInputS6xD(109)(2) <= VNStageIntLLROutputS5xD(177)(1);
  CNStageIntLLRInputS6xD(147)(2) <= VNStageIntLLROutputS5xD(177)(2);
  CNStageIntLLRInputS6xD(204)(2) <= VNStageIntLLROutputS5xD(177)(3);
  CNStageIntLLRInputS6xD(232)(2) <= VNStageIntLLROutputS5xD(177)(4);
  CNStageIntLLRInputS6xD(304)(2) <= VNStageIntLLROutputS5xD(177)(5);
  CNStageIntLLRInputS6xD(368)(2) <= VNStageIntLLROutputS5xD(177)(6);
  CNStageIntLLRInputS6xD(5)(2) <= VNStageIntLLROutputS5xD(178)(0);
  CNStageIntLLRInputS6xD(107)(2) <= VNStageIntLLROutputS5xD(178)(1);
  CNStageIntLLRInputS6xD(142)(2) <= VNStageIntLLROutputS5xD(178)(2);
  CNStageIntLLRInputS6xD(201)(2) <= VNStageIntLLROutputS5xD(178)(3);
  CNStageIntLLRInputS6xD(313)(2) <= VNStageIntLLROutputS5xD(178)(4);
  CNStageIntLLRInputS6xD(338)(2) <= VNStageIntLLROutputS5xD(178)(5);
  CNStageIntLLRInputS6xD(4)(2) <= VNStageIntLLROutputS5xD(179)(0);
  CNStageIntLLRInputS6xD(87)(2) <= VNStageIntLLROutputS5xD(179)(1);
  CNStageIntLLRInputS6xD(148)(2) <= VNStageIntLLROutputS5xD(179)(2);
  CNStageIntLLRInputS6xD(215)(2) <= VNStageIntLLROutputS5xD(179)(3);
  CNStageIntLLRInputS6xD(267)(2) <= VNStageIntLLROutputS5xD(179)(4);
  CNStageIntLLRInputS6xD(308)(2) <= VNStageIntLLROutputS5xD(179)(5);
  CNStageIntLLRInputS6xD(67)(2) <= VNStageIntLLROutputS5xD(180)(0);
  CNStageIntLLRInputS6xD(208)(2) <= VNStageIntLLROutputS5xD(180)(1);
  CNStageIntLLRInputS6xD(263)(2) <= VNStageIntLLROutputS5xD(180)(2);
  CNStageIntLLRInputS6xD(314)(2) <= VNStageIntLLROutputS5xD(180)(3);
  CNStageIntLLRInputS6xD(371)(2) <= VNStageIntLLROutputS5xD(180)(4);
  CNStageIntLLRInputS6xD(3)(2) <= VNStageIntLLROutputS5xD(181)(0);
  CNStageIntLLRInputS6xD(70)(2) <= VNStageIntLLROutputS5xD(181)(1);
  CNStageIntLLRInputS6xD(162)(2) <= VNStageIntLLROutputS5xD(181)(2);
  CNStageIntLLRInputS6xD(186)(2) <= VNStageIntLLROutputS5xD(181)(3);
  CNStageIntLLRInputS6xD(227)(2) <= VNStageIntLLROutputS5xD(181)(4);
  CNStageIntLLRInputS6xD(303)(2) <= VNStageIntLLROutputS5xD(181)(5);
  CNStageIntLLRInputS6xD(2)(2) <= VNStageIntLLROutputS5xD(182)(0);
  CNStageIntLLRInputS6xD(54)(2) <= VNStageIntLLROutputS5xD(182)(1);
  CNStageIntLLRInputS6xD(169)(2) <= VNStageIntLLROutputS5xD(182)(2);
  CNStageIntLLRInputS6xD(195)(2) <= VNStageIntLLROutputS5xD(182)(3);
  CNStageIntLLRInputS6xD(248)(2) <= VNStageIntLLROutputS5xD(182)(4);
  CNStageIntLLRInputS6xD(328)(2) <= VNStageIntLLROutputS5xD(182)(5);
  CNStageIntLLRInputS6xD(350)(2) <= VNStageIntLLROutputS5xD(182)(6);
  CNStageIntLLRInputS6xD(1)(2) <= VNStageIntLLROutputS5xD(183)(0);
  CNStageIntLLRInputS6xD(88)(2) <= VNStageIntLLROutputS5xD(183)(1);
  CNStageIntLLRInputS6xD(190)(2) <= VNStageIntLLROutputS5xD(183)(2);
  CNStageIntLLRInputS6xD(281)(2) <= VNStageIntLLROutputS5xD(183)(3);
  CNStageIntLLRInputS6xD(358)(2) <= VNStageIntLLROutputS5xD(183)(4);
  CNStageIntLLRInputS6xD(0)(2) <= VNStageIntLLROutputS5xD(184)(0);
  CNStageIntLLRInputS6xD(106)(2) <= VNStageIntLLROutputS5xD(184)(1);
  CNStageIntLLRInputS6xD(153)(2) <= VNStageIntLLROutputS5xD(184)(2);
  CNStageIntLLRInputS6xD(193)(2) <= VNStageIntLLROutputS5xD(184)(3);
  CNStageIntLLRInputS6xD(226)(2) <= VNStageIntLLROutputS5xD(184)(4);
  CNStageIntLLRInputS6xD(318)(2) <= VNStageIntLLROutputS5xD(184)(5);
  CNStageIntLLRInputS6xD(354)(2) <= VNStageIntLLROutputS5xD(184)(6);
  CNStageIntLLRInputS6xD(121)(2) <= VNStageIntLLROutputS5xD(185)(0);
  CNStageIntLLRInputS6xD(272)(2) <= VNStageIntLLROutputS5xD(185)(1);
  CNStageIntLLRInputS6xD(320)(2) <= VNStageIntLLROutputS5xD(185)(2);
  CNStageIntLLRInputS6xD(359)(2) <= VNStageIntLLROutputS5xD(185)(3);
  CNStageIntLLRInputS6xD(63)(2) <= VNStageIntLLROutputS5xD(186)(0);
  CNStageIntLLRInputS6xD(160)(2) <= VNStageIntLLROutputS5xD(186)(1);
  CNStageIntLLRInputS6xD(216)(2) <= VNStageIntLLROutputS5xD(186)(2);
  CNStageIntLLRInputS6xD(235)(2) <= VNStageIntLLROutputS5xD(186)(3);
  CNStageIntLLRInputS6xD(290)(2) <= VNStageIntLLROutputS5xD(186)(4);
  CNStageIntLLRInputS6xD(349)(2) <= VNStageIntLLROutputS5xD(186)(5);
  CNStageIntLLRInputS6xD(90)(2) <= VNStageIntLLROutputS5xD(187)(0);
  CNStageIntLLRInputS6xD(113)(2) <= VNStageIntLLROutputS5xD(187)(1);
  CNStageIntLLRInputS6xD(200)(2) <= VNStageIntLLROutputS5xD(187)(2);
  CNStageIntLLRInputS6xD(240)(2) <= VNStageIntLLROutputS5xD(187)(3);
  CNStageIntLLRInputS6xD(326)(2) <= VNStageIntLLROutputS5xD(187)(4);
  CNStageIntLLRInputS6xD(374)(2) <= VNStageIntLLROutputS5xD(187)(5);
  CNStageIntLLRInputS6xD(81)(2) <= VNStageIntLLROutputS5xD(188)(0);
  CNStageIntLLRInputS6xD(212)(2) <= VNStageIntLLROutputS5xD(188)(1);
  CNStageIntLLRInputS6xD(279)(2) <= VNStageIntLLROutputS5xD(188)(2);
  CNStageIntLLRInputS6xD(284)(2) <= VNStageIntLLROutputS5xD(188)(3);
  CNStageIntLLRInputS6xD(381)(2) <= VNStageIntLLROutputS5xD(188)(4);
  CNStageIntLLRInputS6xD(68)(2) <= VNStageIntLLROutputS5xD(189)(0);
  CNStageIntLLRInputS6xD(152)(2) <= VNStageIntLLROutputS5xD(189)(1);
  CNStageIntLLRInputS6xD(223)(2) <= VNStageIntLLROutputS5xD(189)(2);
  CNStageIntLLRInputS6xD(239)(2) <= VNStageIntLLROutputS5xD(189)(3);
  CNStageIntLLRInputS6xD(291)(2) <= VNStageIntLLROutputS5xD(189)(4);
  CNStageIntLLRInputS6xD(363)(2) <= VNStageIntLLROutputS5xD(189)(5);
  CNStageIntLLRInputS6xD(168)(2) <= VNStageIntLLROutputS5xD(190)(0);
  CNStageIntLLRInputS6xD(196)(2) <= VNStageIntLLROutputS5xD(190)(1);
  CNStageIntLLRInputS6xD(234)(2) <= VNStageIntLLROutputS5xD(190)(2);
  CNStageIntLLRInputS6xD(319)(2) <= VNStageIntLLROutputS5xD(190)(3);
  CNStageIntLLRInputS6xD(365)(2) <= VNStageIntLLROutputS5xD(190)(4);
  CNStageIntLLRInputS6xD(52)(2) <= VNStageIntLLROutputS5xD(191)(0);
  CNStageIntLLRInputS6xD(59)(2) <= VNStageIntLLROutputS5xD(191)(1);
  CNStageIntLLRInputS6xD(138)(2) <= VNStageIntLLROutputS5xD(191)(2);
  CNStageIntLLRInputS6xD(185)(2) <= VNStageIntLLROutputS5xD(191)(3);
  CNStageIntLLRInputS6xD(270)(2) <= VNStageIntLLROutputS5xD(191)(4);
  CNStageIntLLRInputS6xD(280)(2) <= VNStageIntLLROutputS5xD(191)(5);
  CNStageIntLLRInputS6xD(53)(3) <= VNStageIntLLROutputS5xD(192)(0);
  CNStageIntLLRInputS6xD(107)(3) <= VNStageIntLLROutputS5xD(192)(1);
  CNStageIntLLRInputS6xD(128)(3) <= VNStageIntLLROutputS5xD(192)(2);
  CNStageIntLLRInputS6xD(197)(3) <= VNStageIntLLROutputS5xD(192)(3);
  CNStageIntLLRInputS6xD(243)(3) <= VNStageIntLLROutputS5xD(192)(4);
  CNStageIntLLRInputS6xD(297)(3) <= VNStageIntLLROutputS5xD(192)(5);
  CNStageIntLLRInputS6xD(340)(3) <= VNStageIntLLROutputS5xD(192)(6);
  CNStageIntLLRInputS6xD(51)(3) <= VNStageIntLLROutputS5xD(193)(0);
  CNStageIntLLRInputS6xD(58)(3) <= VNStageIntLLROutputS5xD(193)(1);
  CNStageIntLLRInputS6xD(137)(3) <= VNStageIntLLROutputS5xD(193)(2);
  CNStageIntLLRInputS6xD(269)(3) <= VNStageIntLLROutputS5xD(193)(3);
  CNStageIntLLRInputS6xD(333)(3) <= VNStageIntLLROutputS5xD(193)(4);
  CNStageIntLLRInputS6xD(50)(3) <= VNStageIntLLROutputS5xD(194)(0);
  CNStageIntLLRInputS6xD(55)(3) <= VNStageIntLLROutputS5xD(194)(1);
  CNStageIntLLRInputS6xD(115)(3) <= VNStageIntLLROutputS5xD(194)(2);
  CNStageIntLLRInputS6xD(171)(3) <= VNStageIntLLROutputS5xD(194)(3);
  CNStageIntLLRInputS6xD(275)(3) <= VNStageIntLLROutputS5xD(194)(4);
  CNStageIntLLRInputS6xD(304)(3) <= VNStageIntLLROutputS5xD(194)(5);
  CNStageIntLLRInputS6xD(371)(3) <= VNStageIntLLROutputS5xD(194)(6);
  CNStageIntLLRInputS6xD(72)(3) <= VNStageIntLLROutputS5xD(195)(0);
  CNStageIntLLRInputS6xD(139)(3) <= VNStageIntLLROutputS5xD(195)(1);
  CNStageIntLLRInputS6xD(187)(3) <= VNStageIntLLROutputS5xD(195)(2);
  CNStageIntLLRInputS6xD(244)(3) <= VNStageIntLLROutputS5xD(195)(3);
  CNStageIntLLRInputS6xD(49)(3) <= VNStageIntLLROutputS5xD(196)(0);
  CNStageIntLLRInputS6xD(64)(3) <= VNStageIntLLROutputS5xD(196)(1);
  CNStageIntLLRInputS6xD(153)(3) <= VNStageIntLLROutputS5xD(196)(2);
  CNStageIntLLRInputS6xD(205)(3) <= VNStageIntLLROutputS5xD(196)(3);
  CNStageIntLLRInputS6xD(242)(3) <= VNStageIntLLROutputS5xD(196)(4);
  CNStageIntLLRInputS6xD(306)(3) <= VNStageIntLLROutputS5xD(196)(5);
  CNStageIntLLRInputS6xD(48)(3) <= VNStageIntLLROutputS5xD(197)(0);
  CNStageIntLLRInputS6xD(96)(3) <= VNStageIntLLROutputS5xD(197)(1);
  CNStageIntLLRInputS6xD(150)(3) <= VNStageIntLLROutputS5xD(197)(2);
  CNStageIntLLRInputS6xD(213)(3) <= VNStageIntLLROutputS5xD(197)(3);
  CNStageIntLLRInputS6xD(273)(3) <= VNStageIntLLROutputS5xD(197)(4);
  CNStageIntLLRInputS6xD(320)(3) <= VNStageIntLLROutputS5xD(197)(5);
  CNStageIntLLRInputS6xD(363)(3) <= VNStageIntLLROutputS5xD(197)(6);
  CNStageIntLLRInputS6xD(47)(3) <= VNStageIntLLROutputS5xD(198)(0);
  CNStageIntLLRInputS6xD(105)(3) <= VNStageIntLLROutputS5xD(198)(1);
  CNStageIntLLRInputS6xD(111)(3) <= VNStageIntLLROutputS5xD(198)(2);
  CNStageIntLLRInputS6xD(208)(3) <= VNStageIntLLROutputS5xD(198)(3);
  CNStageIntLLRInputS6xD(254)(3) <= VNStageIntLLROutputS5xD(198)(4);
  CNStageIntLLRInputS6xD(316)(3) <= VNStageIntLLROutputS5xD(198)(5);
  CNStageIntLLRInputS6xD(379)(3) <= VNStageIntLLROutputS5xD(198)(6);
  CNStageIntLLRInputS6xD(46)(3) <= VNStageIntLLROutputS5xD(199)(0);
  CNStageIntLLRInputS6xD(99)(3) <= VNStageIntLLROutputS5xD(199)(1);
  CNStageIntLLRInputS6xD(133)(3) <= VNStageIntLLROutputS5xD(199)(2);
  CNStageIntLLRInputS6xD(214)(3) <= VNStageIntLLROutputS5xD(199)(3);
  CNStageIntLLRInputS6xD(257)(3) <= VNStageIntLLROutputS5xD(199)(4);
  CNStageIntLLRInputS6xD(282)(3) <= VNStageIntLLROutputS5xD(199)(5);
  CNStageIntLLRInputS6xD(350)(3) <= VNStageIntLLROutputS5xD(199)(6);
  CNStageIntLLRInputS6xD(45)(3) <= VNStageIntLLROutputS5xD(200)(0);
  CNStageIntLLRInputS6xD(102)(3) <= VNStageIntLLROutputS5xD(200)(1);
  CNStageIntLLRInputS6xD(134)(3) <= VNStageIntLLROutputS5xD(200)(2);
  CNStageIntLLRInputS6xD(204)(3) <= VNStageIntLLROutputS5xD(200)(3);
  CNStageIntLLRInputS6xD(245)(3) <= VNStageIntLLROutputS5xD(200)(4);
  CNStageIntLLRInputS6xD(300)(3) <= VNStageIntLLROutputS5xD(200)(5);
  CNStageIntLLRInputS6xD(44)(3) <= VNStageIntLLROutputS5xD(201)(0);
  CNStageIntLLRInputS6xD(93)(3) <= VNStageIntLLROutputS5xD(201)(1);
  CNStageIntLLRInputS6xD(169)(3) <= VNStageIntLLROutputS5xD(201)(2);
  CNStageIntLLRInputS6xD(174)(3) <= VNStageIntLLROutputS5xD(201)(3);
  CNStageIntLLRInputS6xD(274)(3) <= VNStageIntLLROutputS5xD(201)(4);
  CNStageIntLLRInputS6xD(351)(3) <= VNStageIntLLROutputS5xD(201)(5);
  CNStageIntLLRInputS6xD(43)(3) <= VNStageIntLLROutputS5xD(202)(0);
  CNStageIntLLRInputS6xD(73)(3) <= VNStageIntLLROutputS5xD(202)(1);
  CNStageIntLLRInputS6xD(160)(3) <= VNStageIntLLROutputS5xD(202)(2);
  CNStageIntLLRInputS6xD(181)(3) <= VNStageIntLLROutputS5xD(202)(3);
  CNStageIntLLRInputS6xD(281)(3) <= VNStageIntLLROutputS5xD(202)(4);
  CNStageIntLLRInputS6xD(365)(3) <= VNStageIntLLROutputS5xD(202)(5);
  CNStageIntLLRInputS6xD(42)(3) <= VNStageIntLLROutputS5xD(203)(0);
  CNStageIntLLRInputS6xD(54)(3) <= VNStageIntLLROutputS5xD(203)(1);
  CNStageIntLLRInputS6xD(119)(3) <= VNStageIntLLROutputS5xD(203)(2);
  CNStageIntLLRInputS6xD(217)(3) <= VNStageIntLLROutputS5xD(203)(3);
  CNStageIntLLRInputS6xD(267)(3) <= VNStageIntLLROutputS5xD(203)(4);
  CNStageIntLLRInputS6xD(326)(3) <= VNStageIntLLROutputS5xD(203)(5);
  CNStageIntLLRInputS6xD(361)(3) <= VNStageIntLLROutputS5xD(203)(6);
  CNStageIntLLRInputS6xD(41)(3) <= VNStageIntLLROutputS5xD(204)(0);
  CNStageIntLLRInputS6xD(68)(3) <= VNStageIntLLROutputS5xD(204)(1);
  CNStageIntLLRInputS6xD(123)(3) <= VNStageIntLLROutputS5xD(204)(2);
  CNStageIntLLRInputS6xD(219)(3) <= VNStageIntLLROutputS5xD(204)(3);
  CNStageIntLLRInputS6xD(251)(3) <= VNStageIntLLROutputS5xD(204)(4);
  CNStageIntLLRInputS6xD(288)(3) <= VNStageIntLLROutputS5xD(204)(5);
  CNStageIntLLRInputS6xD(382)(3) <= VNStageIntLLROutputS5xD(204)(6);
  CNStageIntLLRInputS6xD(170)(3) <= VNStageIntLLROutputS5xD(205)(0);
  CNStageIntLLRInputS6xD(276)(3) <= VNStageIntLLROutputS5xD(205)(1);
  CNStageIntLLRInputS6xD(345)(3) <= VNStageIntLLROutputS5xD(205)(2);
  CNStageIntLLRInputS6xD(40)(3) <= VNStageIntLLROutputS5xD(206)(0);
  CNStageIntLLRInputS6xD(122)(3) <= VNStageIntLLROutputS5xD(206)(1);
  CNStageIntLLRInputS6xD(172)(3) <= VNStageIntLLROutputS5xD(206)(2);
  CNStageIntLLRInputS6xD(332)(3) <= VNStageIntLLROutputS5xD(206)(3);
  CNStageIntLLRInputS6xD(346)(3) <= VNStageIntLLROutputS5xD(206)(4);
  CNStageIntLLRInputS6xD(39)(3) <= VNStageIntLLROutputS5xD(207)(0);
  CNStageIntLLRInputS6xD(95)(3) <= VNStageIntLLROutputS5xD(207)(1);
  CNStageIntLLRInputS6xD(117)(3) <= VNStageIntLLROutputS5xD(207)(2);
  CNStageIntLLRInputS6xD(255)(3) <= VNStageIntLLROutputS5xD(207)(3);
  CNStageIntLLRInputS6xD(292)(3) <= VNStageIntLLROutputS5xD(207)(4);
  CNStageIntLLRInputS6xD(381)(3) <= VNStageIntLLROutputS5xD(207)(5);
  CNStageIntLLRInputS6xD(38)(3) <= VNStageIntLLROutputS5xD(208)(0);
  CNStageIntLLRInputS6xD(82)(3) <= VNStageIntLLROutputS5xD(208)(1);
  CNStageIntLLRInputS6xD(157)(3) <= VNStageIntLLROutputS5xD(208)(2);
  CNStageIntLLRInputS6xD(191)(3) <= VNStageIntLLROutputS5xD(208)(3);
  CNStageIntLLRInputS6xD(286)(3) <= VNStageIntLLROutputS5xD(208)(4);
  CNStageIntLLRInputS6xD(372)(3) <= VNStageIntLLROutputS5xD(208)(5);
  CNStageIntLLRInputS6xD(37)(3) <= VNStageIntLLROutputS5xD(209)(0);
  CNStageIntLLRInputS6xD(97)(3) <= VNStageIntLLROutputS5xD(209)(1);
  CNStageIntLLRInputS6xD(165)(3) <= VNStageIntLLROutputS5xD(209)(2);
  CNStageIntLLRInputS6xD(218)(3) <= VNStageIntLLROutputS5xD(209)(3);
  CNStageIntLLRInputS6xD(323)(3) <= VNStageIntLLROutputS5xD(209)(4);
  CNStageIntLLRInputS6xD(36)(3) <= VNStageIntLLROutputS5xD(210)(0);
  CNStageIntLLRInputS6xD(60)(3) <= VNStageIntLLROutputS5xD(210)(1);
  CNStageIntLLRInputS6xD(129)(3) <= VNStageIntLLROutputS5xD(210)(2);
  CNStageIntLLRInputS6xD(180)(3) <= VNStageIntLLROutputS5xD(210)(3);
  CNStageIntLLRInputS6xD(246)(3) <= VNStageIntLLROutputS5xD(210)(4);
  CNStageIntLLRInputS6xD(330)(3) <= VNStageIntLLROutputS5xD(210)(5);
  CNStageIntLLRInputS6xD(335)(3) <= VNStageIntLLROutputS5xD(210)(6);
  CNStageIntLLRInputS6xD(35)(3) <= VNStageIntLLROutputS5xD(211)(0);
  CNStageIntLLRInputS6xD(70)(3) <= VNStageIntLLROutputS5xD(211)(1);
  CNStageIntLLRInputS6xD(127)(3) <= VNStageIntLLROutputS5xD(211)(2);
  CNStageIntLLRInputS6xD(206)(3) <= VNStageIntLLROutputS5xD(211)(3);
  CNStageIntLLRInputS6xD(260)(3) <= VNStageIntLLROutputS5xD(211)(4);
  CNStageIntLLRInputS6xD(298)(3) <= VNStageIntLLROutputS5xD(211)(5);
  CNStageIntLLRInputS6xD(34)(3) <= VNStageIntLLROutputS5xD(212)(0);
  CNStageIntLLRInputS6xD(65)(3) <= VNStageIntLLROutputS5xD(212)(1);
  CNStageIntLLRInputS6xD(163)(3) <= VNStageIntLLROutputS5xD(212)(2);
  CNStageIntLLRInputS6xD(186)(3) <= VNStageIntLLROutputS5xD(212)(3);
  CNStageIntLLRInputS6xD(296)(3) <= VNStageIntLLROutputS5xD(212)(4);
  CNStageIntLLRInputS6xD(33)(3) <= VNStageIntLLROutputS5xD(213)(0);
  CNStageIntLLRInputS6xD(71)(3) <= VNStageIntLLROutputS5xD(213)(1);
  CNStageIntLLRInputS6xD(142)(3) <= VNStageIntLLROutputS5xD(213)(2);
  CNStageIntLLRInputS6xD(230)(3) <= VNStageIntLLROutputS5xD(213)(3);
  CNStageIntLLRInputS6xD(32)(3) <= VNStageIntLLROutputS5xD(214)(0);
  CNStageIntLLRInputS6xD(59)(3) <= VNStageIntLLROutputS5xD(214)(1);
  CNStageIntLLRInputS6xD(145)(3) <= VNStageIntLLROutputS5xD(214)(2);
  CNStageIntLLRInputS6xD(220)(3) <= VNStageIntLLROutputS5xD(214)(3);
  CNStageIntLLRInputS6xD(240)(3) <= VNStageIntLLROutputS5xD(214)(4);
  CNStageIntLLRInputS6xD(308)(3) <= VNStageIntLLROutputS5xD(214)(5);
  CNStageIntLLRInputS6xD(369)(3) <= VNStageIntLLROutputS5xD(214)(6);
  CNStageIntLLRInputS6xD(31)(3) <= VNStageIntLLROutputS5xD(215)(0);
  CNStageIntLLRInputS6xD(85)(3) <= VNStageIntLLROutputS5xD(215)(1);
  CNStageIntLLRInputS6xD(130)(3) <= VNStageIntLLROutputS5xD(215)(2);
  CNStageIntLLRInputS6xD(216)(3) <= VNStageIntLLROutputS5xD(215)(3);
  CNStageIntLLRInputS6xD(234)(3) <= VNStageIntLLROutputS5xD(215)(4);
  CNStageIntLLRInputS6xD(311)(3) <= VNStageIntLLROutputS5xD(215)(5);
  CNStageIntLLRInputS6xD(377)(3) <= VNStageIntLLROutputS5xD(215)(6);
  CNStageIntLLRInputS6xD(30)(3) <= VNStageIntLLROutputS5xD(216)(0);
  CNStageIntLLRInputS6xD(91)(3) <= VNStageIntLLROutputS5xD(216)(1);
  CNStageIntLLRInputS6xD(164)(3) <= VNStageIntLLROutputS5xD(216)(2);
  CNStageIntLLRInputS6xD(183)(3) <= VNStageIntLLROutputS5xD(216)(3);
  CNStageIntLLRInputS6xD(237)(3) <= VNStageIntLLROutputS5xD(216)(4);
  CNStageIntLLRInputS6xD(299)(3) <= VNStageIntLLROutputS5xD(216)(5);
  CNStageIntLLRInputS6xD(341)(3) <= VNStageIntLLROutputS5xD(216)(6);
  CNStageIntLLRInputS6xD(29)(3) <= VNStageIntLLROutputS5xD(217)(0);
  CNStageIntLLRInputS6xD(75)(3) <= VNStageIntLLROutputS5xD(217)(1);
  CNStageIntLLRInputS6xD(126)(3) <= VNStageIntLLROutputS5xD(217)(2);
  CNStageIntLLRInputS6xD(201)(3) <= VNStageIntLLROutputS5xD(217)(3);
  CNStageIntLLRInputS6xD(227)(3) <= VNStageIntLLROutputS5xD(217)(4);
  CNStageIntLLRInputS6xD(329)(3) <= VNStageIntLLROutputS5xD(217)(5);
  CNStageIntLLRInputS6xD(339)(3) <= VNStageIntLLROutputS5xD(217)(6);
  CNStageIntLLRInputS6xD(28)(3) <= VNStageIntLLROutputS5xD(218)(0);
  CNStageIntLLRInputS6xD(77)(3) <= VNStageIntLLROutputS5xD(218)(1);
  CNStageIntLLRInputS6xD(154)(3) <= VNStageIntLLROutputS5xD(218)(2);
  CNStageIntLLRInputS6xD(202)(3) <= VNStageIntLLROutputS5xD(218)(3);
  CNStageIntLLRInputS6xD(261)(3) <= VNStageIntLLROutputS5xD(218)(4);
  CNStageIntLLRInputS6xD(295)(3) <= VNStageIntLLROutputS5xD(218)(5);
  CNStageIntLLRInputS6xD(375)(3) <= VNStageIntLLROutputS5xD(218)(6);
  CNStageIntLLRInputS6xD(27)(3) <= VNStageIntLLROutputS5xD(219)(0);
  CNStageIntLLRInputS6xD(101)(3) <= VNStageIntLLROutputS5xD(219)(1);
  CNStageIntLLRInputS6xD(138)(3) <= VNStageIntLLROutputS5xD(219)(2);
  CNStageIntLLRInputS6xD(182)(3) <= VNStageIntLLROutputS5xD(219)(3);
  CNStageIntLLRInputS6xD(321)(3) <= VNStageIntLLROutputS5xD(219)(4);
  CNStageIntLLRInputS6xD(354)(3) <= VNStageIntLLROutputS5xD(219)(5);
  CNStageIntLLRInputS6xD(26)(3) <= VNStageIntLLROutputS5xD(220)(0);
  CNStageIntLLRInputS6xD(83)(3) <= VNStageIntLLROutputS5xD(220)(1);
  CNStageIntLLRInputS6xD(166)(3) <= VNStageIntLLROutputS5xD(220)(2);
  CNStageIntLLRInputS6xD(173)(3) <= VNStageIntLLROutputS5xD(220)(3);
  CNStageIntLLRInputS6xD(256)(3) <= VNStageIntLLROutputS5xD(220)(4);
  CNStageIntLLRInputS6xD(305)(3) <= VNStageIntLLROutputS5xD(220)(5);
  CNStageIntLLRInputS6xD(356)(3) <= VNStageIntLLROutputS5xD(220)(6);
  CNStageIntLLRInputS6xD(25)(3) <= VNStageIntLLROutputS5xD(221)(0);
  CNStageIntLLRInputS6xD(94)(3) <= VNStageIntLLROutputS5xD(221)(1);
  CNStageIntLLRInputS6xD(156)(3) <= VNStageIntLLROutputS5xD(221)(2);
  CNStageIntLLRInputS6xD(190)(3) <= VNStageIntLLROutputS5xD(221)(3);
  CNStageIntLLRInputS6xD(268)(3) <= VNStageIntLLROutputS5xD(221)(4);
  CNStageIntLLRInputS6xD(331)(3) <= VNStageIntLLROutputS5xD(221)(5);
  CNStageIntLLRInputS6xD(342)(3) <= VNStageIntLLROutputS5xD(221)(6);
  CNStageIntLLRInputS6xD(24)(3) <= VNStageIntLLROutputS5xD(222)(0);
  CNStageIntLLRInputS6xD(143)(3) <= VNStageIntLLROutputS5xD(222)(1);
  CNStageIntLLRInputS6xD(241)(3) <= VNStageIntLLROutputS5xD(222)(2);
  CNStageIntLLRInputS6xD(376)(3) <= VNStageIntLLROutputS5xD(222)(3);
  CNStageIntLLRInputS6xD(23)(3) <= VNStageIntLLROutputS5xD(223)(0);
  CNStageIntLLRInputS6xD(76)(3) <= VNStageIntLLROutputS5xD(223)(1);
  CNStageIntLLRInputS6xD(162)(3) <= VNStageIntLLROutputS5xD(223)(2);
  CNStageIntLLRInputS6xD(224)(3) <= VNStageIntLLROutputS5xD(223)(3);
  CNStageIntLLRInputS6xD(229)(3) <= VNStageIntLLROutputS5xD(223)(4);
  CNStageIntLLRInputS6xD(309)(3) <= VNStageIntLLROutputS5xD(223)(5);
  CNStageIntLLRInputS6xD(338)(3) <= VNStageIntLLROutputS5xD(223)(6);
  CNStageIntLLRInputS6xD(22)(3) <= VNStageIntLLROutputS5xD(224)(0);
  CNStageIntLLRInputS6xD(90)(3) <= VNStageIntLLROutputS5xD(224)(1);
  CNStageIntLLRInputS6xD(135)(3) <= VNStageIntLLROutputS5xD(224)(2);
  CNStageIntLLRInputS6xD(193)(3) <= VNStageIntLLROutputS5xD(224)(3);
  CNStageIntLLRInputS6xD(270)(3) <= VNStageIntLLROutputS5xD(224)(4);
  CNStageIntLLRInputS6xD(328)(3) <= VNStageIntLLROutputS5xD(224)(5);
  CNStageIntLLRInputS6xD(366)(3) <= VNStageIntLLROutputS5xD(224)(6);
  CNStageIntLLRInputS6xD(21)(3) <= VNStageIntLLROutputS5xD(225)(0);
  CNStageIntLLRInputS6xD(61)(3) <= VNStageIntLLROutputS5xD(225)(1);
  CNStageIntLLRInputS6xD(132)(3) <= VNStageIntLLROutputS5xD(225)(2);
  CNStageIntLLRInputS6xD(188)(3) <= VNStageIntLLROutputS5xD(225)(3);
  CNStageIntLLRInputS6xD(232)(3) <= VNStageIntLLROutputS5xD(225)(4);
  CNStageIntLLRInputS6xD(301)(3) <= VNStageIntLLROutputS5xD(225)(5);
  CNStageIntLLRInputS6xD(20)(3) <= VNStageIntLLROutputS5xD(226)(0);
  CNStageIntLLRInputS6xD(148)(3) <= VNStageIntLLROutputS5xD(226)(1);
  CNStageIntLLRInputS6xD(378)(3) <= VNStageIntLLROutputS5xD(226)(2);
  CNStageIntLLRInputS6xD(19)(3) <= VNStageIntLLROutputS5xD(227)(0);
  CNStageIntLLRInputS6xD(63)(3) <= VNStageIntLLROutputS5xD(227)(1);
  CNStageIntLLRInputS6xD(140)(3) <= VNStageIntLLROutputS5xD(227)(2);
  CNStageIntLLRInputS6xD(178)(3) <= VNStageIntLLROutputS5xD(227)(3);
  CNStageIntLLRInputS6xD(258)(3) <= VNStageIntLLROutputS5xD(227)(4);
  CNStageIntLLRInputS6xD(314)(3) <= VNStageIntLLROutputS5xD(227)(5);
  CNStageIntLLRInputS6xD(368)(3) <= VNStageIntLLROutputS5xD(227)(6);
  CNStageIntLLRInputS6xD(18)(3) <= VNStageIntLLROutputS5xD(228)(0);
  CNStageIntLLRInputS6xD(78)(3) <= VNStageIntLLROutputS5xD(228)(1);
  CNStageIntLLRInputS6xD(114)(3) <= VNStageIntLLROutputS5xD(228)(2);
  CNStageIntLLRInputS6xD(198)(3) <= VNStageIntLLROutputS5xD(228)(3);
  CNStageIntLLRInputS6xD(253)(3) <= VNStageIntLLROutputS5xD(228)(4);
  CNStageIntLLRInputS6xD(307)(3) <= VNStageIntLLROutputS5xD(228)(5);
  CNStageIntLLRInputS6xD(17)(3) <= VNStageIntLLROutputS5xD(229)(0);
  CNStageIntLLRInputS6xD(74)(3) <= VNStageIntLLROutputS5xD(229)(1);
  CNStageIntLLRInputS6xD(124)(3) <= VNStageIntLLROutputS5xD(229)(2);
  CNStageIntLLRInputS6xD(259)(3) <= VNStageIntLLROutputS5xD(229)(3);
  CNStageIntLLRInputS6xD(374)(3) <= VNStageIntLLROutputS5xD(229)(4);
  CNStageIntLLRInputS6xD(16)(3) <= VNStageIntLLROutputS5xD(230)(0);
  CNStageIntLLRInputS6xD(118)(3) <= VNStageIntLLROutputS5xD(230)(1);
  CNStageIntLLRInputS6xD(176)(3) <= VNStageIntLLROutputS5xD(230)(2);
  CNStageIntLLRInputS6xD(249)(3) <= VNStageIntLLROutputS5xD(230)(3);
  CNStageIntLLRInputS6xD(293)(3) <= VNStageIntLLROutputS5xD(230)(4);
  CNStageIntLLRInputS6xD(347)(3) <= VNStageIntLLROutputS5xD(230)(5);
  CNStageIntLLRInputS6xD(15)(3) <= VNStageIntLLROutputS5xD(231)(0);
  CNStageIntLLRInputS6xD(56)(3) <= VNStageIntLLROutputS5xD(231)(1);
  CNStageIntLLRInputS6xD(209)(3) <= VNStageIntLLROutputS5xD(231)(2);
  CNStageIntLLRInputS6xD(272)(3) <= VNStageIntLLROutputS5xD(231)(3);
  CNStageIntLLRInputS6xD(287)(3) <= VNStageIntLLROutputS5xD(231)(4);
  CNStageIntLLRInputS6xD(344)(3) <= VNStageIntLLROutputS5xD(231)(5);
  CNStageIntLLRInputS6xD(14)(3) <= VNStageIntLLROutputS5xD(232)(0);
  CNStageIntLLRInputS6xD(57)(3) <= VNStageIntLLROutputS5xD(232)(1);
  CNStageIntLLRInputS6xD(212)(3) <= VNStageIntLLROutputS5xD(232)(2);
  CNStageIntLLRInputS6xD(278)(3) <= VNStageIntLLROutputS5xD(232)(3);
  CNStageIntLLRInputS6xD(291)(3) <= VNStageIntLLROutputS5xD(232)(4);
  CNStageIntLLRInputS6xD(359)(3) <= VNStageIntLLROutputS5xD(232)(5);
  CNStageIntLLRInputS6xD(13)(3) <= VNStageIntLLROutputS5xD(233)(0);
  CNStageIntLLRInputS6xD(92)(3) <= VNStageIntLLROutputS5xD(233)(1);
  CNStageIntLLRInputS6xD(149)(3) <= VNStageIntLLROutputS5xD(233)(2);
  CNStageIntLLRInputS6xD(263)(3) <= VNStageIntLLROutputS5xD(233)(3);
  CNStageIntLLRInputS6xD(352)(3) <= VNStageIntLLROutputS5xD(233)(4);
  CNStageIntLLRInputS6xD(12)(3) <= VNStageIntLLROutputS5xD(234)(0);
  CNStageIntLLRInputS6xD(84)(3) <= VNStageIntLLROutputS5xD(234)(1);
  CNStageIntLLRInputS6xD(131)(3) <= VNStageIntLLROutputS5xD(234)(2);
  CNStageIntLLRInputS6xD(177)(3) <= VNStageIntLLROutputS5xD(234)(3);
  CNStageIntLLRInputS6xD(265)(3) <= VNStageIntLLROutputS5xD(234)(4);
  CNStageIntLLRInputS6xD(315)(3) <= VNStageIntLLROutputS5xD(234)(5);
  CNStageIntLLRInputS6xD(100)(3) <= VNStageIntLLROutputS5xD(235)(0);
  CNStageIntLLRInputS6xD(144)(3) <= VNStageIntLLROutputS5xD(235)(1);
  CNStageIntLLRInputS6xD(196)(3) <= VNStageIntLLROutputS5xD(235)(2);
  CNStageIntLLRInputS6xD(235)(3) <= VNStageIntLLROutputS5xD(235)(3);
  CNStageIntLLRInputS6xD(336)(3) <= VNStageIntLLROutputS5xD(235)(4);
  CNStageIntLLRInputS6xD(11)(3) <= VNStageIntLLROutputS5xD(236)(0);
  CNStageIntLLRInputS6xD(104)(3) <= VNStageIntLLROutputS5xD(236)(1);
  CNStageIntLLRInputS6xD(155)(3) <= VNStageIntLLROutputS5xD(236)(2);
  CNStageIntLLRInputS6xD(221)(3) <= VNStageIntLLROutputS5xD(236)(3);
  CNStageIntLLRInputS6xD(271)(3) <= VNStageIntLLROutputS5xD(236)(4);
  CNStageIntLLRInputS6xD(310)(3) <= VNStageIntLLROutputS5xD(236)(5);
  CNStageIntLLRInputS6xD(10)(3) <= VNStageIntLLROutputS5xD(237)(0);
  CNStageIntLLRInputS6xD(110)(3) <= VNStageIntLLROutputS5xD(237)(1);
  CNStageIntLLRInputS6xD(125)(3) <= VNStageIntLLROutputS5xD(237)(2);
  CNStageIntLLRInputS6xD(228)(3) <= VNStageIntLLROutputS5xD(237)(3);
  CNStageIntLLRInputS6xD(322)(3) <= VNStageIntLLROutputS5xD(237)(4);
  CNStageIntLLRInputS6xD(334)(3) <= VNStageIntLLROutputS5xD(237)(5);
  CNStageIntLLRInputS6xD(9)(3) <= VNStageIntLLROutputS5xD(238)(0);
  CNStageIntLLRInputS6xD(103)(3) <= VNStageIntLLROutputS5xD(238)(1);
  CNStageIntLLRInputS6xD(113)(3) <= VNStageIntLLROutputS5xD(238)(2);
  CNStageIntLLRInputS6xD(179)(3) <= VNStageIntLLROutputS5xD(238)(3);
  CNStageIntLLRInputS6xD(236)(3) <= VNStageIntLLROutputS5xD(238)(4);
  CNStageIntLLRInputS6xD(294)(3) <= VNStageIntLLROutputS5xD(238)(5);
  CNStageIntLLRInputS6xD(383)(3) <= VNStageIntLLROutputS5xD(238)(6);
  CNStageIntLLRInputS6xD(8)(3) <= VNStageIntLLROutputS5xD(239)(0);
  CNStageIntLLRInputS6xD(98)(3) <= VNStageIntLLROutputS5xD(239)(1);
  CNStageIntLLRInputS6xD(158)(3) <= VNStageIntLLROutputS5xD(239)(2);
  CNStageIntLLRInputS6xD(223)(3) <= VNStageIntLLROutputS5xD(239)(3);
  CNStageIntLLRInputS6xD(264)(3) <= VNStageIntLLROutputS5xD(239)(4);
  CNStageIntLLRInputS6xD(284)(3) <= VNStageIntLLROutputS5xD(239)(5);
  CNStageIntLLRInputS6xD(360)(3) <= VNStageIntLLROutputS5xD(239)(6);
  CNStageIntLLRInputS6xD(7)(3) <= VNStageIntLLROutputS5xD(240)(0);
  CNStageIntLLRInputS6xD(81)(3) <= VNStageIntLLROutputS5xD(240)(1);
  CNStageIntLLRInputS6xD(116)(3) <= VNStageIntLLROutputS5xD(240)(2);
  CNStageIntLLRInputS6xD(210)(3) <= VNStageIntLLROutputS5xD(240)(3);
  CNStageIntLLRInputS6xD(277)(3) <= VNStageIntLLROutputS5xD(240)(4);
  CNStageIntLLRInputS6xD(324)(3) <= VNStageIntLLROutputS5xD(240)(5);
  CNStageIntLLRInputS6xD(343)(3) <= VNStageIntLLROutputS5xD(240)(6);
  CNStageIntLLRInputS6xD(6)(3) <= VNStageIntLLROutputS5xD(241)(0);
  CNStageIntLLRInputS6xD(88)(3) <= VNStageIntLLROutputS5xD(241)(1);
  CNStageIntLLRInputS6xD(175)(3) <= VNStageIntLLROutputS5xD(241)(2);
  CNStageIntLLRInputS6xD(250)(3) <= VNStageIntLLROutputS5xD(241)(3);
  CNStageIntLLRInputS6xD(285)(3) <= VNStageIntLLROutputS5xD(241)(4);
  CNStageIntLLRInputS6xD(355)(3) <= VNStageIntLLROutputS5xD(241)(5);
  CNStageIntLLRInputS6xD(5)(3) <= VNStageIntLLROutputS5xD(242)(0);
  CNStageIntLLRInputS6xD(108)(3) <= VNStageIntLLROutputS5xD(242)(1);
  CNStageIntLLRInputS6xD(146)(3) <= VNStageIntLLROutputS5xD(242)(2);
  CNStageIntLLRInputS6xD(203)(3) <= VNStageIntLLROutputS5xD(242)(3);
  CNStageIntLLRInputS6xD(231)(3) <= VNStageIntLLROutputS5xD(242)(4);
  CNStageIntLLRInputS6xD(303)(3) <= VNStageIntLLROutputS5xD(242)(5);
  CNStageIntLLRInputS6xD(367)(3) <= VNStageIntLLROutputS5xD(242)(6);
  CNStageIntLLRInputS6xD(4)(3) <= VNStageIntLLROutputS5xD(243)(0);
  CNStageIntLLRInputS6xD(106)(3) <= VNStageIntLLROutputS5xD(243)(1);
  CNStageIntLLRInputS6xD(141)(3) <= VNStageIntLLROutputS5xD(243)(2);
  CNStageIntLLRInputS6xD(200)(3) <= VNStageIntLLROutputS5xD(243)(3);
  CNStageIntLLRInputS6xD(252)(3) <= VNStageIntLLROutputS5xD(243)(4);
  CNStageIntLLRInputS6xD(312)(3) <= VNStageIntLLROutputS5xD(243)(5);
  CNStageIntLLRInputS6xD(337)(3) <= VNStageIntLLROutputS5xD(243)(6);
  CNStageIntLLRInputS6xD(147)(3) <= VNStageIntLLROutputS5xD(244)(0);
  CNStageIntLLRInputS6xD(266)(3) <= VNStageIntLLROutputS5xD(244)(1);
  CNStageIntLLRInputS6xD(3)(3) <= VNStageIntLLROutputS5xD(245)(0);
  CNStageIntLLRInputS6xD(66)(3) <= VNStageIntLLROutputS5xD(245)(1);
  CNStageIntLLRInputS6xD(136)(3) <= VNStageIntLLROutputS5xD(245)(2);
  CNStageIntLLRInputS6xD(207)(3) <= VNStageIntLLROutputS5xD(245)(3);
  CNStageIntLLRInputS6xD(262)(3) <= VNStageIntLLROutputS5xD(245)(4);
  CNStageIntLLRInputS6xD(313)(3) <= VNStageIntLLROutputS5xD(245)(5);
  CNStageIntLLRInputS6xD(370)(3) <= VNStageIntLLROutputS5xD(245)(6);
  CNStageIntLLRInputS6xD(2)(3) <= VNStageIntLLROutputS5xD(246)(0);
  CNStageIntLLRInputS6xD(69)(3) <= VNStageIntLLROutputS5xD(246)(1);
  CNStageIntLLRInputS6xD(161)(3) <= VNStageIntLLROutputS5xD(246)(2);
  CNStageIntLLRInputS6xD(185)(3) <= VNStageIntLLROutputS5xD(246)(3);
  CNStageIntLLRInputS6xD(226)(3) <= VNStageIntLLROutputS5xD(246)(4);
  CNStageIntLLRInputS6xD(302)(3) <= VNStageIntLLROutputS5xD(246)(5);
  CNStageIntLLRInputS6xD(1)(3) <= VNStageIntLLROutputS5xD(247)(0);
  CNStageIntLLRInputS6xD(109)(3) <= VNStageIntLLROutputS5xD(247)(1);
  CNStageIntLLRInputS6xD(168)(3) <= VNStageIntLLROutputS5xD(247)(2);
  CNStageIntLLRInputS6xD(194)(3) <= VNStageIntLLROutputS5xD(247)(3);
  CNStageIntLLRInputS6xD(247)(3) <= VNStageIntLLROutputS5xD(247)(4);
  CNStageIntLLRInputS6xD(327)(3) <= VNStageIntLLROutputS5xD(247)(5);
  CNStageIntLLRInputS6xD(349)(3) <= VNStageIntLLROutputS5xD(247)(6);
  CNStageIntLLRInputS6xD(0)(3) <= VNStageIntLLROutputS5xD(248)(0);
  CNStageIntLLRInputS6xD(87)(3) <= VNStageIntLLROutputS5xD(248)(1);
  CNStageIntLLRInputS6xD(151)(3) <= VNStageIntLLROutputS5xD(248)(2);
  CNStageIntLLRInputS6xD(189)(3) <= VNStageIntLLROutputS5xD(248)(3);
  CNStageIntLLRInputS6xD(248)(3) <= VNStageIntLLROutputS5xD(248)(4);
  CNStageIntLLRInputS6xD(280)(3) <= VNStageIntLLROutputS5xD(248)(5);
  CNStageIntLLRInputS6xD(357)(3) <= VNStageIntLLROutputS5xD(248)(6);
  CNStageIntLLRInputS6xD(152)(3) <= VNStageIntLLROutputS5xD(249)(0);
  CNStageIntLLRInputS6xD(192)(3) <= VNStageIntLLROutputS5xD(249)(1);
  CNStageIntLLRInputS6xD(225)(3) <= VNStageIntLLROutputS5xD(249)(2);
  CNStageIntLLRInputS6xD(317)(3) <= VNStageIntLLROutputS5xD(249)(3);
  CNStageIntLLRInputS6xD(353)(3) <= VNStageIntLLROutputS5xD(249)(4);
  CNStageIntLLRInputS6xD(79)(3) <= VNStageIntLLROutputS5xD(250)(0);
  CNStageIntLLRInputS6xD(120)(3) <= VNStageIntLLROutputS5xD(250)(1);
  CNStageIntLLRInputS6xD(184)(3) <= VNStageIntLLROutputS5xD(250)(2);
  CNStageIntLLRInputS6xD(319)(3) <= VNStageIntLLROutputS5xD(250)(3);
  CNStageIntLLRInputS6xD(358)(3) <= VNStageIntLLROutputS5xD(250)(4);
  CNStageIntLLRInputS6xD(62)(3) <= VNStageIntLLROutputS5xD(251)(0);
  CNStageIntLLRInputS6xD(159)(3) <= VNStageIntLLROutputS5xD(251)(1);
  CNStageIntLLRInputS6xD(215)(3) <= VNStageIntLLROutputS5xD(251)(2);
  CNStageIntLLRInputS6xD(289)(3) <= VNStageIntLLROutputS5xD(251)(3);
  CNStageIntLLRInputS6xD(348)(3) <= VNStageIntLLROutputS5xD(251)(4);
  CNStageIntLLRInputS6xD(89)(3) <= VNStageIntLLROutputS5xD(252)(0);
  CNStageIntLLRInputS6xD(112)(3) <= VNStageIntLLROutputS5xD(252)(1);
  CNStageIntLLRInputS6xD(199)(3) <= VNStageIntLLROutputS5xD(252)(2);
  CNStageIntLLRInputS6xD(239)(3) <= VNStageIntLLROutputS5xD(252)(3);
  CNStageIntLLRInputS6xD(325)(3) <= VNStageIntLLROutputS5xD(252)(4);
  CNStageIntLLRInputS6xD(373)(3) <= VNStageIntLLROutputS5xD(252)(5);
  CNStageIntLLRInputS6xD(80)(3) <= VNStageIntLLROutputS5xD(253)(0);
  CNStageIntLLRInputS6xD(121)(3) <= VNStageIntLLROutputS5xD(253)(1);
  CNStageIntLLRInputS6xD(211)(3) <= VNStageIntLLROutputS5xD(253)(2);
  CNStageIntLLRInputS6xD(279)(3) <= VNStageIntLLROutputS5xD(253)(3);
  CNStageIntLLRInputS6xD(283)(3) <= VNStageIntLLROutputS5xD(253)(4);
  CNStageIntLLRInputS6xD(380)(3) <= VNStageIntLLROutputS5xD(253)(5);
  CNStageIntLLRInputS6xD(67)(3) <= VNStageIntLLROutputS5xD(254)(0);
  CNStageIntLLRInputS6xD(222)(3) <= VNStageIntLLROutputS5xD(254)(1);
  CNStageIntLLRInputS6xD(238)(3) <= VNStageIntLLROutputS5xD(254)(2);
  CNStageIntLLRInputS6xD(290)(3) <= VNStageIntLLROutputS5xD(254)(3);
  CNStageIntLLRInputS6xD(362)(3) <= VNStageIntLLROutputS5xD(254)(4);
  CNStageIntLLRInputS6xD(52)(3) <= VNStageIntLLROutputS5xD(255)(0);
  CNStageIntLLRInputS6xD(86)(3) <= VNStageIntLLROutputS5xD(255)(1);
  CNStageIntLLRInputS6xD(167)(3) <= VNStageIntLLROutputS5xD(255)(2);
  CNStageIntLLRInputS6xD(195)(3) <= VNStageIntLLROutputS5xD(255)(3);
  CNStageIntLLRInputS6xD(233)(3) <= VNStageIntLLROutputS5xD(255)(4);
  CNStageIntLLRInputS6xD(318)(3) <= VNStageIntLLROutputS5xD(255)(5);
  CNStageIntLLRInputS6xD(364)(3) <= VNStageIntLLROutputS5xD(255)(6);
  CNStageIntLLRInputS6xD(53)(4) <= VNStageIntLLROutputS5xD(256)(0);
  CNStageIntLLRInputS6xD(106)(4) <= VNStageIntLLROutputS5xD(256)(1);
  CNStageIntLLRInputS6xD(127)(4) <= VNStageIntLLROutputS5xD(256)(2);
  CNStageIntLLRInputS6xD(242)(4) <= VNStageIntLLROutputS5xD(256)(3);
  CNStageIntLLRInputS6xD(296)(4) <= VNStageIntLLROutputS5xD(256)(4);
  CNStageIntLLRInputS6xD(339)(4) <= VNStageIntLLROutputS5xD(256)(5);
  CNStageIntLLRInputS6xD(51)(4) <= VNStageIntLLROutputS5xD(257)(0);
  CNStageIntLLRInputS6xD(85)(4) <= VNStageIntLLROutputS5xD(257)(1);
  CNStageIntLLRInputS6xD(166)(4) <= VNStageIntLLROutputS5xD(257)(2);
  CNStageIntLLRInputS6xD(194)(4) <= VNStageIntLLROutputS5xD(257)(3);
  CNStageIntLLRInputS6xD(232)(4) <= VNStageIntLLROutputS5xD(257)(4);
  CNStageIntLLRInputS6xD(317)(4) <= VNStageIntLLROutputS5xD(257)(5);
  CNStageIntLLRInputS6xD(363)(4) <= VNStageIntLLROutputS5xD(257)(6);
  CNStageIntLLRInputS6xD(50)(4) <= VNStageIntLLROutputS5xD(258)(0);
  CNStageIntLLRInputS6xD(57)(4) <= VNStageIntLLROutputS5xD(258)(1);
  CNStageIntLLRInputS6xD(331)(4) <= VNStageIntLLROutputS5xD(258)(2);
  CNStageIntLLRInputS6xD(54)(4) <= VNStageIntLLROutputS5xD(259)(0);
  CNStageIntLLRInputS6xD(114)(4) <= VNStageIntLLROutputS5xD(259)(1);
  CNStageIntLLRInputS6xD(274)(4) <= VNStageIntLLROutputS5xD(259)(2);
  CNStageIntLLRInputS6xD(303)(4) <= VNStageIntLLROutputS5xD(259)(3);
  CNStageIntLLRInputS6xD(370)(4) <= VNStageIntLLROutputS5xD(259)(4);
  CNStageIntLLRInputS6xD(49)(4) <= VNStageIntLLROutputS5xD(260)(0);
  CNStageIntLLRInputS6xD(71)(4) <= VNStageIntLLROutputS5xD(260)(1);
  CNStageIntLLRInputS6xD(138)(4) <= VNStageIntLLROutputS5xD(260)(2);
  CNStageIntLLRInputS6xD(186)(4) <= VNStageIntLLROutputS5xD(260)(3);
  CNStageIntLLRInputS6xD(243)(4) <= VNStageIntLLROutputS5xD(260)(4);
  CNStageIntLLRInputS6xD(383)(4) <= VNStageIntLLROutputS5xD(260)(5);
  CNStageIntLLRInputS6xD(48)(4) <= VNStageIntLLROutputS5xD(261)(0);
  CNStageIntLLRInputS6xD(63)(4) <= VNStageIntLLROutputS5xD(261)(1);
  CNStageIntLLRInputS6xD(152)(4) <= VNStageIntLLROutputS5xD(261)(2);
  CNStageIntLLRInputS6xD(204)(4) <= VNStageIntLLROutputS5xD(261)(3);
  CNStageIntLLRInputS6xD(305)(4) <= VNStageIntLLROutputS5xD(261)(4);
  CNStageIntLLRInputS6xD(333)(4) <= VNStageIntLLROutputS5xD(261)(5);
  CNStageIntLLRInputS6xD(47)(4) <= VNStageIntLLROutputS5xD(262)(0);
  CNStageIntLLRInputS6xD(95)(4) <= VNStageIntLLROutputS5xD(262)(1);
  CNStageIntLLRInputS6xD(149)(4) <= VNStageIntLLROutputS5xD(262)(2);
  CNStageIntLLRInputS6xD(212)(4) <= VNStageIntLLROutputS5xD(262)(3);
  CNStageIntLLRInputS6xD(319)(4) <= VNStageIntLLROutputS5xD(262)(4);
  CNStageIntLLRInputS6xD(362)(4) <= VNStageIntLLROutputS5xD(262)(5);
  CNStageIntLLRInputS6xD(46)(4) <= VNStageIntLLROutputS5xD(263)(0);
  CNStageIntLLRInputS6xD(104)(4) <= VNStageIntLLROutputS5xD(263)(1);
  CNStageIntLLRInputS6xD(169)(4) <= VNStageIntLLROutputS5xD(263)(2);
  CNStageIntLLRInputS6xD(207)(4) <= VNStageIntLLROutputS5xD(263)(3);
  CNStageIntLLRInputS6xD(253)(4) <= VNStageIntLLROutputS5xD(263)(4);
  CNStageIntLLRInputS6xD(315)(4) <= VNStageIntLLROutputS5xD(263)(5);
  CNStageIntLLRInputS6xD(378)(4) <= VNStageIntLLROutputS5xD(263)(6);
  CNStageIntLLRInputS6xD(45)(4) <= VNStageIntLLROutputS5xD(264)(0);
  CNStageIntLLRInputS6xD(98)(4) <= VNStageIntLLROutputS5xD(264)(1);
  CNStageIntLLRInputS6xD(132)(4) <= VNStageIntLLROutputS5xD(264)(2);
  CNStageIntLLRInputS6xD(213)(4) <= VNStageIntLLROutputS5xD(264)(3);
  CNStageIntLLRInputS6xD(256)(4) <= VNStageIntLLROutputS5xD(264)(4);
  CNStageIntLLRInputS6xD(281)(4) <= VNStageIntLLROutputS5xD(264)(5);
  CNStageIntLLRInputS6xD(349)(4) <= VNStageIntLLROutputS5xD(264)(6);
  CNStageIntLLRInputS6xD(44)(4) <= VNStageIntLLROutputS5xD(265)(0);
  CNStageIntLLRInputS6xD(133)(4) <= VNStageIntLLROutputS5xD(265)(1);
  CNStageIntLLRInputS6xD(203)(4) <= VNStageIntLLROutputS5xD(265)(2);
  CNStageIntLLRInputS6xD(244)(4) <= VNStageIntLLROutputS5xD(265)(3);
  CNStageIntLLRInputS6xD(43)(4) <= VNStageIntLLROutputS5xD(266)(0);
  CNStageIntLLRInputS6xD(168)(4) <= VNStageIntLLROutputS5xD(266)(1);
  CNStageIntLLRInputS6xD(173)(4) <= VNStageIntLLROutputS5xD(266)(2);
  CNStageIntLLRInputS6xD(273)(4) <= VNStageIntLLROutputS5xD(266)(3);
  CNStageIntLLRInputS6xD(300)(4) <= VNStageIntLLROutputS5xD(266)(4);
  CNStageIntLLRInputS6xD(42)(4) <= VNStageIntLLROutputS5xD(267)(0);
  CNStageIntLLRInputS6xD(72)(4) <= VNStageIntLLROutputS5xD(267)(1);
  CNStageIntLLRInputS6xD(159)(4) <= VNStageIntLLROutputS5xD(267)(2);
  CNStageIntLLRInputS6xD(180)(4) <= VNStageIntLLROutputS5xD(267)(3);
  CNStageIntLLRInputS6xD(241)(4) <= VNStageIntLLROutputS5xD(267)(4);
  CNStageIntLLRInputS6xD(280)(4) <= VNStageIntLLROutputS5xD(267)(5);
  CNStageIntLLRInputS6xD(364)(4) <= VNStageIntLLROutputS5xD(267)(6);
  CNStageIntLLRInputS6xD(41)(4) <= VNStageIntLLROutputS5xD(268)(0);
  CNStageIntLLRInputS6xD(109)(4) <= VNStageIntLLROutputS5xD(268)(1);
  CNStageIntLLRInputS6xD(118)(4) <= VNStageIntLLROutputS5xD(268)(2);
  CNStageIntLLRInputS6xD(216)(4) <= VNStageIntLLROutputS5xD(268)(3);
  CNStageIntLLRInputS6xD(266)(4) <= VNStageIntLLROutputS5xD(268)(4);
  CNStageIntLLRInputS6xD(325)(4) <= VNStageIntLLROutputS5xD(268)(5);
  CNStageIntLLRInputS6xD(360)(4) <= VNStageIntLLROutputS5xD(268)(6);
  CNStageIntLLRInputS6xD(67)(4) <= VNStageIntLLROutputS5xD(269)(0);
  CNStageIntLLRInputS6xD(122)(4) <= VNStageIntLLROutputS5xD(269)(1);
  CNStageIntLLRInputS6xD(218)(4) <= VNStageIntLLROutputS5xD(269)(2);
  CNStageIntLLRInputS6xD(250)(4) <= VNStageIntLLROutputS5xD(269)(3);
  CNStageIntLLRInputS6xD(287)(4) <= VNStageIntLLROutputS5xD(269)(4);
  CNStageIntLLRInputS6xD(381)(4) <= VNStageIntLLROutputS5xD(269)(5);
  CNStageIntLLRInputS6xD(40)(4) <= VNStageIntLLROutputS5xD(270)(0);
  CNStageIntLLRInputS6xD(79)(4) <= VNStageIntLLROutputS5xD(270)(1);
  CNStageIntLLRInputS6xD(170)(4) <= VNStageIntLLROutputS5xD(270)(2);
  CNStageIntLLRInputS6xD(190)(4) <= VNStageIntLLROutputS5xD(270)(3);
  CNStageIntLLRInputS6xD(275)(4) <= VNStageIntLLROutputS5xD(270)(4);
  CNStageIntLLRInputS6xD(292)(4) <= VNStageIntLLROutputS5xD(270)(5);
  CNStageIntLLRInputS6xD(344)(4) <= VNStageIntLLROutputS5xD(270)(6);
  CNStageIntLLRInputS6xD(39)(4) <= VNStageIntLLROutputS5xD(271)(0);
  CNStageIntLLRInputS6xD(105)(4) <= VNStageIntLLROutputS5xD(271)(1);
  CNStageIntLLRInputS6xD(171)(4) <= VNStageIntLLROutputS5xD(271)(2);
  CNStageIntLLRInputS6xD(268)(4) <= VNStageIntLLROutputS5xD(271)(3);
  CNStageIntLLRInputS6xD(332)(4) <= VNStageIntLLROutputS5xD(271)(4);
  CNStageIntLLRInputS6xD(345)(4) <= VNStageIntLLROutputS5xD(271)(5);
  CNStageIntLLRInputS6xD(38)(4) <= VNStageIntLLROutputS5xD(272)(0);
  CNStageIntLLRInputS6xD(94)(4) <= VNStageIntLLROutputS5xD(272)(1);
  CNStageIntLLRInputS6xD(116)(4) <= VNStageIntLLROutputS5xD(272)(2);
  CNStageIntLLRInputS6xD(184)(4) <= VNStageIntLLROutputS5xD(272)(3);
  CNStageIntLLRInputS6xD(254)(4) <= VNStageIntLLROutputS5xD(272)(4);
  CNStageIntLLRInputS6xD(291)(4) <= VNStageIntLLROutputS5xD(272)(5);
  CNStageIntLLRInputS6xD(380)(4) <= VNStageIntLLROutputS5xD(272)(6);
  CNStageIntLLRInputS6xD(37)(4) <= VNStageIntLLROutputS5xD(273)(0);
  CNStageIntLLRInputS6xD(81)(4) <= VNStageIntLLROutputS5xD(273)(1);
  CNStageIntLLRInputS6xD(156)(4) <= VNStageIntLLROutputS5xD(273)(2);
  CNStageIntLLRInputS6xD(272)(4) <= VNStageIntLLROutputS5xD(273)(3);
  CNStageIntLLRInputS6xD(285)(4) <= VNStageIntLLROutputS5xD(273)(4);
  CNStageIntLLRInputS6xD(371)(4) <= VNStageIntLLROutputS5xD(273)(5);
  CNStageIntLLRInputS6xD(36)(4) <= VNStageIntLLROutputS5xD(274)(0);
  CNStageIntLLRInputS6xD(164)(4) <= VNStageIntLLROutputS5xD(274)(1);
  CNStageIntLLRInputS6xD(217)(4) <= VNStageIntLLROutputS5xD(274)(2);
  CNStageIntLLRInputS6xD(248)(4) <= VNStageIntLLROutputS5xD(274)(3);
  CNStageIntLLRInputS6xD(35)(4) <= VNStageIntLLROutputS5xD(275)(0);
  CNStageIntLLRInputS6xD(59)(4) <= VNStageIntLLROutputS5xD(275)(1);
  CNStageIntLLRInputS6xD(128)(4) <= VNStageIntLLROutputS5xD(275)(2);
  CNStageIntLLRInputS6xD(179)(4) <= VNStageIntLLROutputS5xD(275)(3);
  CNStageIntLLRInputS6xD(329)(4) <= VNStageIntLLROutputS5xD(275)(4);
  CNStageIntLLRInputS6xD(34)(4) <= VNStageIntLLROutputS5xD(276)(0);
  CNStageIntLLRInputS6xD(69)(4) <= VNStageIntLLROutputS5xD(276)(1);
  CNStageIntLLRInputS6xD(126)(4) <= VNStageIntLLROutputS5xD(276)(2);
  CNStageIntLLRInputS6xD(205)(4) <= VNStageIntLLROutputS5xD(276)(3);
  CNStageIntLLRInputS6xD(259)(4) <= VNStageIntLLROutputS5xD(276)(4);
  CNStageIntLLRInputS6xD(297)(4) <= VNStageIntLLROutputS5xD(276)(5);
  CNStageIntLLRInputS6xD(33)(4) <= VNStageIntLLROutputS5xD(277)(0);
  CNStageIntLLRInputS6xD(64)(4) <= VNStageIntLLROutputS5xD(277)(1);
  CNStageIntLLRInputS6xD(162)(4) <= VNStageIntLLROutputS5xD(277)(2);
  CNStageIntLLRInputS6xD(185)(4) <= VNStageIntLLROutputS5xD(277)(3);
  CNStageIntLLRInputS6xD(252)(4) <= VNStageIntLLROutputS5xD(277)(4);
  CNStageIntLLRInputS6xD(295)(4) <= VNStageIntLLROutputS5xD(277)(5);
  CNStageIntLLRInputS6xD(334)(4) <= VNStageIntLLROutputS5xD(277)(6);
  CNStageIntLLRInputS6xD(32)(4) <= VNStageIntLLROutputS5xD(278)(0);
  CNStageIntLLRInputS6xD(70)(4) <= VNStageIntLLROutputS5xD(278)(1);
  CNStageIntLLRInputS6xD(141)(4) <= VNStageIntLLROutputS5xD(278)(2);
  CNStageIntLLRInputS6xD(229)(4) <= VNStageIntLLROutputS5xD(278)(3);
  CNStageIntLLRInputS6xD(328)(4) <= VNStageIntLLROutputS5xD(278)(4);
  CNStageIntLLRInputS6xD(31)(4) <= VNStageIntLLROutputS5xD(279)(0);
  CNStageIntLLRInputS6xD(58)(4) <= VNStageIntLLROutputS5xD(279)(1);
  CNStageIntLLRInputS6xD(144)(4) <= VNStageIntLLROutputS5xD(279)(2);
  CNStageIntLLRInputS6xD(219)(4) <= VNStageIntLLROutputS5xD(279)(3);
  CNStageIntLLRInputS6xD(239)(4) <= VNStageIntLLROutputS5xD(279)(4);
  CNStageIntLLRInputS6xD(368)(4) <= VNStageIntLLROutputS5xD(279)(5);
  CNStageIntLLRInputS6xD(30)(4) <= VNStageIntLLROutputS5xD(280)(0);
  CNStageIntLLRInputS6xD(84)(4) <= VNStageIntLLROutputS5xD(280)(1);
  CNStageIntLLRInputS6xD(129)(4) <= VNStageIntLLROutputS5xD(280)(2);
  CNStageIntLLRInputS6xD(215)(4) <= VNStageIntLLROutputS5xD(280)(3);
  CNStageIntLLRInputS6xD(233)(4) <= VNStageIntLLROutputS5xD(280)(4);
  CNStageIntLLRInputS6xD(310)(4) <= VNStageIntLLROutputS5xD(280)(5);
  CNStageIntLLRInputS6xD(376)(4) <= VNStageIntLLROutputS5xD(280)(6);
  CNStageIntLLRInputS6xD(29)(4) <= VNStageIntLLROutputS5xD(281)(0);
  CNStageIntLLRInputS6xD(90)(4) <= VNStageIntLLROutputS5xD(281)(1);
  CNStageIntLLRInputS6xD(163)(4) <= VNStageIntLLROutputS5xD(281)(2);
  CNStageIntLLRInputS6xD(182)(4) <= VNStageIntLLROutputS5xD(281)(3);
  CNStageIntLLRInputS6xD(236)(4) <= VNStageIntLLROutputS5xD(281)(4);
  CNStageIntLLRInputS6xD(298)(4) <= VNStageIntLLROutputS5xD(281)(5);
  CNStageIntLLRInputS6xD(340)(4) <= VNStageIntLLROutputS5xD(281)(6);
  CNStageIntLLRInputS6xD(28)(4) <= VNStageIntLLROutputS5xD(282)(0);
  CNStageIntLLRInputS6xD(74)(4) <= VNStageIntLLROutputS5xD(282)(1);
  CNStageIntLLRInputS6xD(125)(4) <= VNStageIntLLROutputS5xD(282)(2);
  CNStageIntLLRInputS6xD(200)(4) <= VNStageIntLLROutputS5xD(282)(3);
  CNStageIntLLRInputS6xD(226)(4) <= VNStageIntLLROutputS5xD(282)(4);
  CNStageIntLLRInputS6xD(338)(4) <= VNStageIntLLROutputS5xD(282)(5);
  CNStageIntLLRInputS6xD(27)(4) <= VNStageIntLLROutputS5xD(283)(0);
  CNStageIntLLRInputS6xD(76)(4) <= VNStageIntLLROutputS5xD(283)(1);
  CNStageIntLLRInputS6xD(153)(4) <= VNStageIntLLROutputS5xD(283)(2);
  CNStageIntLLRInputS6xD(201)(4) <= VNStageIntLLROutputS5xD(283)(3);
  CNStageIntLLRInputS6xD(260)(4) <= VNStageIntLLROutputS5xD(283)(4);
  CNStageIntLLRInputS6xD(294)(4) <= VNStageIntLLROutputS5xD(283)(5);
  CNStageIntLLRInputS6xD(374)(4) <= VNStageIntLLROutputS5xD(283)(6);
  CNStageIntLLRInputS6xD(26)(4) <= VNStageIntLLROutputS5xD(284)(0);
  CNStageIntLLRInputS6xD(100)(4) <= VNStageIntLLROutputS5xD(284)(1);
  CNStageIntLLRInputS6xD(137)(4) <= VNStageIntLLROutputS5xD(284)(2);
  CNStageIntLLRInputS6xD(181)(4) <= VNStageIntLLROutputS5xD(284)(3);
  CNStageIntLLRInputS6xD(245)(4) <= VNStageIntLLROutputS5xD(284)(4);
  CNStageIntLLRInputS6xD(320)(4) <= VNStageIntLLROutputS5xD(284)(5);
  CNStageIntLLRInputS6xD(353)(4) <= VNStageIntLLROutputS5xD(284)(6);
  CNStageIntLLRInputS6xD(25)(4) <= VNStageIntLLROutputS5xD(285)(0);
  CNStageIntLLRInputS6xD(82)(4) <= VNStageIntLLROutputS5xD(285)(1);
  CNStageIntLLRInputS6xD(165)(4) <= VNStageIntLLROutputS5xD(285)(2);
  CNStageIntLLRInputS6xD(172)(4) <= VNStageIntLLROutputS5xD(285)(3);
  CNStageIntLLRInputS6xD(255)(4) <= VNStageIntLLROutputS5xD(285)(4);
  CNStageIntLLRInputS6xD(304)(4) <= VNStageIntLLROutputS5xD(285)(5);
  CNStageIntLLRInputS6xD(355)(4) <= VNStageIntLLROutputS5xD(285)(6);
  CNStageIntLLRInputS6xD(24)(4) <= VNStageIntLLROutputS5xD(286)(0);
  CNStageIntLLRInputS6xD(93)(4) <= VNStageIntLLROutputS5xD(286)(1);
  CNStageIntLLRInputS6xD(155)(4) <= VNStageIntLLROutputS5xD(286)(2);
  CNStageIntLLRInputS6xD(189)(4) <= VNStageIntLLROutputS5xD(286)(3);
  CNStageIntLLRInputS6xD(267)(4) <= VNStageIntLLROutputS5xD(286)(4);
  CNStageIntLLRInputS6xD(330)(4) <= VNStageIntLLROutputS5xD(286)(5);
  CNStageIntLLRInputS6xD(341)(4) <= VNStageIntLLROutputS5xD(286)(6);
  CNStageIntLLRInputS6xD(23)(4) <= VNStageIntLLROutputS5xD(287)(0);
  CNStageIntLLRInputS6xD(101)(4) <= VNStageIntLLROutputS5xD(287)(1);
  CNStageIntLLRInputS6xD(142)(4) <= VNStageIntLLROutputS5xD(287)(2);
  CNStageIntLLRInputS6xD(193)(4) <= VNStageIntLLROutputS5xD(287)(3);
  CNStageIntLLRInputS6xD(240)(4) <= VNStageIntLLROutputS5xD(287)(4);
  CNStageIntLLRInputS6xD(322)(4) <= VNStageIntLLROutputS5xD(287)(5);
  CNStageIntLLRInputS6xD(375)(4) <= VNStageIntLLROutputS5xD(287)(6);
  CNStageIntLLRInputS6xD(22)(4) <= VNStageIntLLROutputS5xD(288)(0);
  CNStageIntLLRInputS6xD(75)(4) <= VNStageIntLLROutputS5xD(288)(1);
  CNStageIntLLRInputS6xD(161)(4) <= VNStageIntLLROutputS5xD(288)(2);
  CNStageIntLLRInputS6xD(224)(4) <= VNStageIntLLROutputS5xD(288)(3);
  CNStageIntLLRInputS6xD(228)(4) <= VNStageIntLLROutputS5xD(288)(4);
  CNStageIntLLRInputS6xD(308)(4) <= VNStageIntLLROutputS5xD(288)(5);
  CNStageIntLLRInputS6xD(337)(4) <= VNStageIntLLROutputS5xD(288)(6);
  CNStageIntLLRInputS6xD(21)(4) <= VNStageIntLLROutputS5xD(289)(0);
  CNStageIntLLRInputS6xD(89)(4) <= VNStageIntLLROutputS5xD(289)(1);
  CNStageIntLLRInputS6xD(134)(4) <= VNStageIntLLROutputS5xD(289)(2);
  CNStageIntLLRInputS6xD(192)(4) <= VNStageIntLLROutputS5xD(289)(3);
  CNStageIntLLRInputS6xD(269)(4) <= VNStageIntLLROutputS5xD(289)(4);
  CNStageIntLLRInputS6xD(327)(4) <= VNStageIntLLROutputS5xD(289)(5);
  CNStageIntLLRInputS6xD(365)(4) <= VNStageIntLLROutputS5xD(289)(6);
  CNStageIntLLRInputS6xD(20)(4) <= VNStageIntLLROutputS5xD(290)(0);
  CNStageIntLLRInputS6xD(60)(4) <= VNStageIntLLROutputS5xD(290)(1);
  CNStageIntLLRInputS6xD(131)(4) <= VNStageIntLLROutputS5xD(290)(2);
  CNStageIntLLRInputS6xD(187)(4) <= VNStageIntLLROutputS5xD(290)(3);
  CNStageIntLLRInputS6xD(231)(4) <= VNStageIntLLROutputS5xD(290)(4);
  CNStageIntLLRInputS6xD(350)(4) <= VNStageIntLLROutputS5xD(290)(5);
  CNStageIntLLRInputS6xD(19)(4) <= VNStageIntLLROutputS5xD(291)(0);
  CNStageIntLLRInputS6xD(96)(4) <= VNStageIntLLROutputS5xD(291)(1);
  CNStageIntLLRInputS6xD(147)(4) <= VNStageIntLLROutputS5xD(291)(2);
  CNStageIntLLRInputS6xD(223)(4) <= VNStageIntLLROutputS5xD(291)(3);
  CNStageIntLLRInputS6xD(249)(4) <= VNStageIntLLROutputS5xD(291)(4);
  CNStageIntLLRInputS6xD(377)(4) <= VNStageIntLLROutputS5xD(291)(5);
  CNStageIntLLRInputS6xD(18)(4) <= VNStageIntLLROutputS5xD(292)(0);
  CNStageIntLLRInputS6xD(62)(4) <= VNStageIntLLROutputS5xD(292)(1);
  CNStageIntLLRInputS6xD(139)(4) <= VNStageIntLLROutputS5xD(292)(2);
  CNStageIntLLRInputS6xD(177)(4) <= VNStageIntLLROutputS5xD(292)(3);
  CNStageIntLLRInputS6xD(257)(4) <= VNStageIntLLROutputS5xD(292)(4);
  CNStageIntLLRInputS6xD(313)(4) <= VNStageIntLLROutputS5xD(292)(5);
  CNStageIntLLRInputS6xD(367)(4) <= VNStageIntLLROutputS5xD(292)(6);
  CNStageIntLLRInputS6xD(17)(4) <= VNStageIntLLROutputS5xD(293)(0);
  CNStageIntLLRInputS6xD(77)(4) <= VNStageIntLLROutputS5xD(293)(1);
  CNStageIntLLRInputS6xD(113)(4) <= VNStageIntLLROutputS5xD(293)(2);
  CNStageIntLLRInputS6xD(197)(4) <= VNStageIntLLROutputS5xD(293)(3);
  CNStageIntLLRInputS6xD(306)(4) <= VNStageIntLLROutputS5xD(293)(4);
  CNStageIntLLRInputS6xD(354)(4) <= VNStageIntLLROutputS5xD(293)(5);
  CNStageIntLLRInputS6xD(16)(4) <= VNStageIntLLROutputS5xD(294)(0);
  CNStageIntLLRInputS6xD(73)(4) <= VNStageIntLLROutputS5xD(294)(1);
  CNStageIntLLRInputS6xD(123)(4) <= VNStageIntLLROutputS5xD(294)(2);
  CNStageIntLLRInputS6xD(196)(4) <= VNStageIntLLROutputS5xD(294)(3);
  CNStageIntLLRInputS6xD(258)(4) <= VNStageIntLLROutputS5xD(294)(4);
  CNStageIntLLRInputS6xD(284)(4) <= VNStageIntLLROutputS5xD(294)(5);
  CNStageIntLLRInputS6xD(373)(4) <= VNStageIntLLROutputS5xD(294)(6);
  CNStageIntLLRInputS6xD(15)(4) <= VNStageIntLLROutputS5xD(295)(0);
  CNStageIntLLRInputS6xD(92)(4) <= VNStageIntLLROutputS5xD(295)(1);
  CNStageIntLLRInputS6xD(117)(4) <= VNStageIntLLROutputS5xD(295)(2);
  CNStageIntLLRInputS6xD(175)(4) <= VNStageIntLLROutputS5xD(295)(3);
  CNStageIntLLRInputS6xD(346)(4) <= VNStageIntLLROutputS5xD(295)(4);
  CNStageIntLLRInputS6xD(14)(4) <= VNStageIntLLROutputS5xD(296)(0);
  CNStageIntLLRInputS6xD(55)(4) <= VNStageIntLLROutputS5xD(296)(1);
  CNStageIntLLRInputS6xD(121)(4) <= VNStageIntLLROutputS5xD(296)(2);
  CNStageIntLLRInputS6xD(208)(4) <= VNStageIntLLROutputS5xD(296)(3);
  CNStageIntLLRInputS6xD(286)(4) <= VNStageIntLLROutputS5xD(296)(4);
  CNStageIntLLRInputS6xD(343)(4) <= VNStageIntLLROutputS5xD(296)(5);
  CNStageIntLLRInputS6xD(13)(4) <= VNStageIntLLROutputS5xD(297)(0);
  CNStageIntLLRInputS6xD(56)(4) <= VNStageIntLLROutputS5xD(297)(1);
  CNStageIntLLRInputS6xD(111)(4) <= VNStageIntLLROutputS5xD(297)(2);
  CNStageIntLLRInputS6xD(211)(4) <= VNStageIntLLROutputS5xD(297)(3);
  CNStageIntLLRInputS6xD(277)(4) <= VNStageIntLLROutputS5xD(297)(4);
  CNStageIntLLRInputS6xD(290)(4) <= VNStageIntLLROutputS5xD(297)(5);
  CNStageIntLLRInputS6xD(358)(4) <= VNStageIntLLROutputS5xD(297)(6);
  CNStageIntLLRInputS6xD(12)(4) <= VNStageIntLLROutputS5xD(298)(0);
  CNStageIntLLRInputS6xD(91)(4) <= VNStageIntLLROutputS5xD(298)(1);
  CNStageIntLLRInputS6xD(148)(4) <= VNStageIntLLROutputS5xD(298)(2);
  CNStageIntLLRInputS6xD(198)(4) <= VNStageIntLLROutputS5xD(298)(3);
  CNStageIntLLRInputS6xD(262)(4) <= VNStageIntLLROutputS5xD(298)(4);
  CNStageIntLLRInputS6xD(282)(4) <= VNStageIntLLROutputS5xD(298)(5);
  CNStageIntLLRInputS6xD(351)(4) <= VNStageIntLLROutputS5xD(298)(6);
  CNStageIntLLRInputS6xD(83)(4) <= VNStageIntLLROutputS5xD(299)(0);
  CNStageIntLLRInputS6xD(130)(4) <= VNStageIntLLROutputS5xD(299)(1);
  CNStageIntLLRInputS6xD(176)(4) <= VNStageIntLLROutputS5xD(299)(2);
  CNStageIntLLRInputS6xD(264)(4) <= VNStageIntLLROutputS5xD(299)(3);
  CNStageIntLLRInputS6xD(314)(4) <= VNStageIntLLROutputS5xD(299)(4);
  CNStageIntLLRInputS6xD(11)(4) <= VNStageIntLLROutputS5xD(300)(0);
  CNStageIntLLRInputS6xD(99)(4) <= VNStageIntLLROutputS5xD(300)(1);
  CNStageIntLLRInputS6xD(143)(4) <= VNStageIntLLROutputS5xD(300)(2);
  CNStageIntLLRInputS6xD(195)(4) <= VNStageIntLLROutputS5xD(300)(3);
  CNStageIntLLRInputS6xD(299)(4) <= VNStageIntLLROutputS5xD(300)(4);
  CNStageIntLLRInputS6xD(335)(4) <= VNStageIntLLROutputS5xD(300)(5);
  CNStageIntLLRInputS6xD(10)(4) <= VNStageIntLLROutputS5xD(301)(0);
  CNStageIntLLRInputS6xD(103)(4) <= VNStageIntLLROutputS5xD(301)(1);
  CNStageIntLLRInputS6xD(154)(4) <= VNStageIntLLROutputS5xD(301)(2);
  CNStageIntLLRInputS6xD(220)(4) <= VNStageIntLLROutputS5xD(301)(3);
  CNStageIntLLRInputS6xD(270)(4) <= VNStageIntLLROutputS5xD(301)(4);
  CNStageIntLLRInputS6xD(309)(4) <= VNStageIntLLROutputS5xD(301)(5);
  CNStageIntLLRInputS6xD(9)(4) <= VNStageIntLLROutputS5xD(302)(0);
  CNStageIntLLRInputS6xD(110)(4) <= VNStageIntLLROutputS5xD(302)(1);
  CNStageIntLLRInputS6xD(124)(4) <= VNStageIntLLROutputS5xD(302)(2);
  CNStageIntLLRInputS6xD(206)(4) <= VNStageIntLLROutputS5xD(302)(3);
  CNStageIntLLRInputS6xD(227)(4) <= VNStageIntLLROutputS5xD(302)(4);
  CNStageIntLLRInputS6xD(321)(4) <= VNStageIntLLROutputS5xD(302)(5);
  CNStageIntLLRInputS6xD(8)(4) <= VNStageIntLLROutputS5xD(303)(0);
  CNStageIntLLRInputS6xD(102)(4) <= VNStageIntLLROutputS5xD(303)(1);
  CNStageIntLLRInputS6xD(112)(4) <= VNStageIntLLROutputS5xD(303)(2);
  CNStageIntLLRInputS6xD(178)(4) <= VNStageIntLLROutputS5xD(303)(3);
  CNStageIntLLRInputS6xD(235)(4) <= VNStageIntLLROutputS5xD(303)(4);
  CNStageIntLLRInputS6xD(293)(4) <= VNStageIntLLROutputS5xD(303)(5);
  CNStageIntLLRInputS6xD(382)(4) <= VNStageIntLLROutputS5xD(303)(6);
  CNStageIntLLRInputS6xD(7)(4) <= VNStageIntLLROutputS5xD(304)(0);
  CNStageIntLLRInputS6xD(97)(4) <= VNStageIntLLROutputS5xD(304)(1);
  CNStageIntLLRInputS6xD(157)(4) <= VNStageIntLLROutputS5xD(304)(2);
  CNStageIntLLRInputS6xD(222)(4) <= VNStageIntLLROutputS5xD(304)(3);
  CNStageIntLLRInputS6xD(263)(4) <= VNStageIntLLROutputS5xD(304)(4);
  CNStageIntLLRInputS6xD(283)(4) <= VNStageIntLLROutputS5xD(304)(5);
  CNStageIntLLRInputS6xD(359)(4) <= VNStageIntLLROutputS5xD(304)(6);
  CNStageIntLLRInputS6xD(6)(4) <= VNStageIntLLROutputS5xD(305)(0);
  CNStageIntLLRInputS6xD(80)(4) <= VNStageIntLLROutputS5xD(305)(1);
  CNStageIntLLRInputS6xD(115)(4) <= VNStageIntLLROutputS5xD(305)(2);
  CNStageIntLLRInputS6xD(209)(4) <= VNStageIntLLROutputS5xD(305)(3);
  CNStageIntLLRInputS6xD(276)(4) <= VNStageIntLLROutputS5xD(305)(4);
  CNStageIntLLRInputS6xD(323)(4) <= VNStageIntLLROutputS5xD(305)(5);
  CNStageIntLLRInputS6xD(342)(4) <= VNStageIntLLROutputS5xD(305)(6);
  CNStageIntLLRInputS6xD(5)(4) <= VNStageIntLLROutputS5xD(306)(0);
  CNStageIntLLRInputS6xD(87)(4) <= VNStageIntLLROutputS5xD(306)(1);
  CNStageIntLLRInputS6xD(136)(4) <= VNStageIntLLROutputS5xD(306)(2);
  CNStageIntLLRInputS6xD(174)(4) <= VNStageIntLLROutputS5xD(306)(3);
  CNStageIntLLRInputS6xD(4)(4) <= VNStageIntLLROutputS5xD(307)(0);
  CNStageIntLLRInputS6xD(107)(4) <= VNStageIntLLROutputS5xD(307)(1);
  CNStageIntLLRInputS6xD(145)(4) <= VNStageIntLLROutputS5xD(307)(2);
  CNStageIntLLRInputS6xD(202)(4) <= VNStageIntLLROutputS5xD(307)(3);
  CNStageIntLLRInputS6xD(230)(4) <= VNStageIntLLROutputS5xD(307)(4);
  CNStageIntLLRInputS6xD(302)(4) <= VNStageIntLLROutputS5xD(307)(5);
  CNStageIntLLRInputS6xD(366)(4) <= VNStageIntLLROutputS5xD(307)(6);
  CNStageIntLLRInputS6xD(140)(4) <= VNStageIntLLROutputS5xD(308)(0);
  CNStageIntLLRInputS6xD(199)(4) <= VNStageIntLLROutputS5xD(308)(1);
  CNStageIntLLRInputS6xD(251)(4) <= VNStageIntLLROutputS5xD(308)(2);
  CNStageIntLLRInputS6xD(311)(4) <= VNStageIntLLROutputS5xD(308)(3);
  CNStageIntLLRInputS6xD(336)(4) <= VNStageIntLLROutputS5xD(308)(4);
  CNStageIntLLRInputS6xD(3)(4) <= VNStageIntLLROutputS5xD(309)(0);
  CNStageIntLLRInputS6xD(86)(4) <= VNStageIntLLROutputS5xD(309)(1);
  CNStageIntLLRInputS6xD(146)(4) <= VNStageIntLLROutputS5xD(309)(2);
  CNStageIntLLRInputS6xD(214)(4) <= VNStageIntLLROutputS5xD(309)(3);
  CNStageIntLLRInputS6xD(265)(4) <= VNStageIntLLROutputS5xD(309)(4);
  CNStageIntLLRInputS6xD(307)(4) <= VNStageIntLLROutputS5xD(309)(5);
  CNStageIntLLRInputS6xD(2)(4) <= VNStageIntLLROutputS5xD(310)(0);
  CNStageIntLLRInputS6xD(65)(4) <= VNStageIntLLROutputS5xD(310)(1);
  CNStageIntLLRInputS6xD(135)(4) <= VNStageIntLLROutputS5xD(310)(2);
  CNStageIntLLRInputS6xD(261)(4) <= VNStageIntLLROutputS5xD(310)(3);
  CNStageIntLLRInputS6xD(312)(4) <= VNStageIntLLROutputS5xD(310)(4);
  CNStageIntLLRInputS6xD(369)(4) <= VNStageIntLLROutputS5xD(310)(5);
  CNStageIntLLRInputS6xD(1)(4) <= VNStageIntLLROutputS5xD(311)(0);
  CNStageIntLLRInputS6xD(68)(4) <= VNStageIntLLROutputS5xD(311)(1);
  CNStageIntLLRInputS6xD(160)(4) <= VNStageIntLLROutputS5xD(311)(2);
  CNStageIntLLRInputS6xD(225)(4) <= VNStageIntLLROutputS5xD(311)(3);
  CNStageIntLLRInputS6xD(301)(4) <= VNStageIntLLROutputS5xD(311)(4);
  CNStageIntLLRInputS6xD(0)(4) <= VNStageIntLLROutputS5xD(312)(0);
  CNStageIntLLRInputS6xD(108)(4) <= VNStageIntLLROutputS5xD(312)(1);
  CNStageIntLLRInputS6xD(167)(4) <= VNStageIntLLROutputS5xD(312)(2);
  CNStageIntLLRInputS6xD(246)(4) <= VNStageIntLLROutputS5xD(312)(3);
  CNStageIntLLRInputS6xD(326)(4) <= VNStageIntLLROutputS5xD(312)(4);
  CNStageIntLLRInputS6xD(348)(4) <= VNStageIntLLROutputS5xD(312)(5);
  CNStageIntLLRInputS6xD(150)(4) <= VNStageIntLLROutputS5xD(313)(0);
  CNStageIntLLRInputS6xD(188)(4) <= VNStageIntLLROutputS5xD(313)(1);
  CNStageIntLLRInputS6xD(247)(4) <= VNStageIntLLROutputS5xD(313)(2);
  CNStageIntLLRInputS6xD(356)(4) <= VNStageIntLLROutputS5xD(313)(3);
  CNStageIntLLRInputS6xD(191)(4) <= VNStageIntLLROutputS5xD(314)(0);
  CNStageIntLLRInputS6xD(278)(4) <= VNStageIntLLROutputS5xD(314)(1);
  CNStageIntLLRInputS6xD(316)(4) <= VNStageIntLLROutputS5xD(314)(2);
  CNStageIntLLRInputS6xD(352)(4) <= VNStageIntLLROutputS5xD(314)(3);
  CNStageIntLLRInputS6xD(78)(4) <= VNStageIntLLROutputS5xD(315)(0);
  CNStageIntLLRInputS6xD(119)(4) <= VNStageIntLLROutputS5xD(315)(1);
  CNStageIntLLRInputS6xD(183)(4) <= VNStageIntLLROutputS5xD(315)(2);
  CNStageIntLLRInputS6xD(271)(4) <= VNStageIntLLROutputS5xD(315)(3);
  CNStageIntLLRInputS6xD(318)(4) <= VNStageIntLLROutputS5xD(315)(4);
  CNStageIntLLRInputS6xD(357)(4) <= VNStageIntLLROutputS5xD(315)(5);
  CNStageIntLLRInputS6xD(61)(4) <= VNStageIntLLROutputS5xD(316)(0);
  CNStageIntLLRInputS6xD(158)(4) <= VNStageIntLLROutputS5xD(316)(1);
  CNStageIntLLRInputS6xD(234)(4) <= VNStageIntLLROutputS5xD(316)(2);
  CNStageIntLLRInputS6xD(288)(4) <= VNStageIntLLROutputS5xD(316)(3);
  CNStageIntLLRInputS6xD(347)(4) <= VNStageIntLLROutputS5xD(316)(4);
  CNStageIntLLRInputS6xD(88)(4) <= VNStageIntLLROutputS5xD(317)(0);
  CNStageIntLLRInputS6xD(238)(4) <= VNStageIntLLROutputS5xD(317)(1);
  CNStageIntLLRInputS6xD(324)(4) <= VNStageIntLLROutputS5xD(317)(2);
  CNStageIntLLRInputS6xD(372)(4) <= VNStageIntLLROutputS5xD(317)(3);
  CNStageIntLLRInputS6xD(120)(4) <= VNStageIntLLROutputS5xD(318)(0);
  CNStageIntLLRInputS6xD(210)(4) <= VNStageIntLLROutputS5xD(318)(1);
  CNStageIntLLRInputS6xD(279)(4) <= VNStageIntLLROutputS5xD(318)(2);
  CNStageIntLLRInputS6xD(379)(4) <= VNStageIntLLROutputS5xD(318)(3);
  CNStageIntLLRInputS6xD(52)(4) <= VNStageIntLLROutputS5xD(319)(0);
  CNStageIntLLRInputS6xD(66)(4) <= VNStageIntLLROutputS5xD(319)(1);
  CNStageIntLLRInputS6xD(151)(4) <= VNStageIntLLROutputS5xD(319)(2);
  CNStageIntLLRInputS6xD(221)(4) <= VNStageIntLLROutputS5xD(319)(3);
  CNStageIntLLRInputS6xD(237)(4) <= VNStageIntLLROutputS5xD(319)(4);
  CNStageIntLLRInputS6xD(289)(4) <= VNStageIntLLROutputS5xD(319)(5);
  CNStageIntLLRInputS6xD(361)(4) <= VNStageIntLLROutputS5xD(319)(6);
  CNStageIntLLRInputS6xD(53)(5) <= VNStageIntLLROutputS5xD(320)(0);
  CNStageIntLLRInputS6xD(126)(5) <= VNStageIntLLROutputS5xD(320)(1);
  CNStageIntLLRInputS6xD(196)(5) <= VNStageIntLLROutputS5xD(320)(2);
  CNStageIntLLRInputS6xD(295)(5) <= VNStageIntLLROutputS5xD(320)(3);
  CNStageIntLLRInputS6xD(338)(5) <= VNStageIntLLROutputS5xD(320)(4);
  CNStageIntLLRInputS6xD(51)(5) <= VNStageIntLLROutputS5xD(321)(0);
  CNStageIntLLRInputS6xD(65)(5) <= VNStageIntLLROutputS5xD(321)(1);
  CNStageIntLLRInputS6xD(150)(5) <= VNStageIntLLROutputS5xD(321)(2);
  CNStageIntLLRInputS6xD(220)(5) <= VNStageIntLLROutputS5xD(321)(3);
  CNStageIntLLRInputS6xD(236)(5) <= VNStageIntLLROutputS5xD(321)(4);
  CNStageIntLLRInputS6xD(288)(5) <= VNStageIntLLROutputS5xD(321)(5);
  CNStageIntLLRInputS6xD(360)(5) <= VNStageIntLLROutputS5xD(321)(6);
  CNStageIntLLRInputS6xD(50)(5) <= VNStageIntLLROutputS5xD(322)(0);
  CNStageIntLLRInputS6xD(84)(5) <= VNStageIntLLROutputS5xD(322)(1);
  CNStageIntLLRInputS6xD(165)(5) <= VNStageIntLLROutputS5xD(322)(2);
  CNStageIntLLRInputS6xD(231)(5) <= VNStageIntLLROutputS5xD(322)(3);
  CNStageIntLLRInputS6xD(316)(5) <= VNStageIntLLROutputS5xD(322)(4);
  CNStageIntLLRInputS6xD(362)(5) <= VNStageIntLLROutputS5xD(322)(5);
  CNStageIntLLRInputS6xD(56)(5) <= VNStageIntLLROutputS5xD(323)(0);
  CNStageIntLLRInputS6xD(136)(5) <= VNStageIntLLROutputS5xD(323)(1);
  CNStageIntLLRInputS6xD(184)(5) <= VNStageIntLLROutputS5xD(323)(2);
  CNStageIntLLRInputS6xD(268)(5) <= VNStageIntLLROutputS5xD(323)(3);
  CNStageIntLLRInputS6xD(330)(5) <= VNStageIntLLROutputS5xD(323)(4);
  CNStageIntLLRInputS6xD(49)(5) <= VNStageIntLLROutputS5xD(324)(0);
  CNStageIntLLRInputS6xD(109)(5) <= VNStageIntLLROutputS5xD(324)(1);
  CNStageIntLLRInputS6xD(113)(5) <= VNStageIntLLROutputS5xD(324)(2);
  CNStageIntLLRInputS6xD(223)(5) <= VNStageIntLLROutputS5xD(324)(3);
  CNStageIntLLRInputS6xD(273)(5) <= VNStageIntLLROutputS5xD(324)(4);
  CNStageIntLLRInputS6xD(302)(5) <= VNStageIntLLROutputS5xD(324)(5);
  CNStageIntLLRInputS6xD(369)(5) <= VNStageIntLLROutputS5xD(324)(6);
  CNStageIntLLRInputS6xD(48)(5) <= VNStageIntLLROutputS5xD(325)(0);
  CNStageIntLLRInputS6xD(70)(5) <= VNStageIntLLROutputS5xD(325)(1);
  CNStageIntLLRInputS6xD(137)(5) <= VNStageIntLLROutputS5xD(325)(2);
  CNStageIntLLRInputS6xD(185)(5) <= VNStageIntLLROutputS5xD(325)(3);
  CNStageIntLLRInputS6xD(242)(5) <= VNStageIntLLROutputS5xD(325)(4);
  CNStageIntLLRInputS6xD(284)(5) <= VNStageIntLLROutputS5xD(325)(5);
  CNStageIntLLRInputS6xD(382)(5) <= VNStageIntLLROutputS5xD(325)(6);
  CNStageIntLLRInputS6xD(47)(5) <= VNStageIntLLROutputS5xD(326)(0);
  CNStageIntLLRInputS6xD(62)(5) <= VNStageIntLLROutputS5xD(326)(1);
  CNStageIntLLRInputS6xD(203)(5) <= VNStageIntLLROutputS5xD(326)(2);
  CNStageIntLLRInputS6xD(241)(5) <= VNStageIntLLROutputS5xD(326)(3);
  CNStageIntLLRInputS6xD(304)(5) <= VNStageIntLLROutputS5xD(326)(4);
  CNStageIntLLRInputS6xD(46)(5) <= VNStageIntLLROutputS5xD(327)(0);
  CNStageIntLLRInputS6xD(94)(5) <= VNStageIntLLROutputS5xD(327)(1);
  CNStageIntLLRInputS6xD(148)(5) <= VNStageIntLLROutputS5xD(327)(2);
  CNStageIntLLRInputS6xD(211)(5) <= VNStageIntLLROutputS5xD(327)(3);
  CNStageIntLLRInputS6xD(272)(5) <= VNStageIntLLROutputS5xD(327)(4);
  CNStageIntLLRInputS6xD(318)(5) <= VNStageIntLLROutputS5xD(327)(5);
  CNStageIntLLRInputS6xD(361)(5) <= VNStageIntLLROutputS5xD(327)(6);
  CNStageIntLLRInputS6xD(45)(5) <= VNStageIntLLROutputS5xD(328)(0);
  CNStageIntLLRInputS6xD(103)(5) <= VNStageIntLLROutputS5xD(328)(1);
  CNStageIntLLRInputS6xD(168)(5) <= VNStageIntLLROutputS5xD(328)(2);
  CNStageIntLLRInputS6xD(314)(5) <= VNStageIntLLROutputS5xD(328)(3);
  CNStageIntLLRInputS6xD(377)(5) <= VNStageIntLLROutputS5xD(328)(4);
  CNStageIntLLRInputS6xD(44)(5) <= VNStageIntLLROutputS5xD(329)(0);
  CNStageIntLLRInputS6xD(97)(5) <= VNStageIntLLROutputS5xD(329)(1);
  CNStageIntLLRInputS6xD(131)(5) <= VNStageIntLLROutputS5xD(329)(2);
  CNStageIntLLRInputS6xD(212)(5) <= VNStageIntLLROutputS5xD(329)(3);
  CNStageIntLLRInputS6xD(255)(5) <= VNStageIntLLROutputS5xD(329)(4);
  CNStageIntLLRInputS6xD(280)(5) <= VNStageIntLLROutputS5xD(329)(5);
  CNStageIntLLRInputS6xD(348)(5) <= VNStageIntLLROutputS5xD(329)(6);
  CNStageIntLLRInputS6xD(43)(5) <= VNStageIntLLROutputS5xD(330)(0);
  CNStageIntLLRInputS6xD(101)(5) <= VNStageIntLLROutputS5xD(330)(1);
  CNStageIntLLRInputS6xD(132)(5) <= VNStageIntLLROutputS5xD(330)(2);
  CNStageIntLLRInputS6xD(202)(5) <= VNStageIntLLROutputS5xD(330)(3);
  CNStageIntLLRInputS6xD(243)(5) <= VNStageIntLLROutputS5xD(330)(4);
  CNStageIntLLRInputS6xD(42)(5) <= VNStageIntLLROutputS5xD(331)(0);
  CNStageIntLLRInputS6xD(92)(5) <= VNStageIntLLROutputS5xD(331)(1);
  CNStageIntLLRInputS6xD(167)(5) <= VNStageIntLLROutputS5xD(331)(2);
  CNStageIntLLRInputS6xD(172)(5) <= VNStageIntLLROutputS5xD(331)(3);
  CNStageIntLLRInputS6xD(350)(5) <= VNStageIntLLROutputS5xD(331)(4);
  CNStageIntLLRInputS6xD(41)(5) <= VNStageIntLLROutputS5xD(332)(0);
  CNStageIntLLRInputS6xD(71)(5) <= VNStageIntLLROutputS5xD(332)(1);
  CNStageIntLLRInputS6xD(158)(5) <= VNStageIntLLROutputS5xD(332)(2);
  CNStageIntLLRInputS6xD(179)(5) <= VNStageIntLLROutputS5xD(332)(3);
  CNStageIntLLRInputS6xD(240)(5) <= VNStageIntLLROutputS5xD(332)(4);
  CNStageIntLLRInputS6xD(363)(5) <= VNStageIntLLROutputS5xD(332)(5);
  CNStageIntLLRInputS6xD(108)(5) <= VNStageIntLLROutputS5xD(333)(0);
  CNStageIntLLRInputS6xD(117)(5) <= VNStageIntLLROutputS5xD(333)(1);
  CNStageIntLLRInputS6xD(215)(5) <= VNStageIntLLROutputS5xD(333)(2);
  CNStageIntLLRInputS6xD(265)(5) <= VNStageIntLLROutputS5xD(333)(3);
  CNStageIntLLRInputS6xD(324)(5) <= VNStageIntLLROutputS5xD(333)(4);
  CNStageIntLLRInputS6xD(359)(5) <= VNStageIntLLROutputS5xD(333)(5);
  CNStageIntLLRInputS6xD(40)(5) <= VNStageIntLLROutputS5xD(334)(0);
  CNStageIntLLRInputS6xD(66)(5) <= VNStageIntLLROutputS5xD(334)(1);
  CNStageIntLLRInputS6xD(217)(5) <= VNStageIntLLROutputS5xD(334)(2);
  CNStageIntLLRInputS6xD(286)(5) <= VNStageIntLLROutputS5xD(334)(3);
  CNStageIntLLRInputS6xD(380)(5) <= VNStageIntLLROutputS5xD(334)(4);
  CNStageIntLLRInputS6xD(39)(5) <= VNStageIntLLROutputS5xD(335)(0);
  CNStageIntLLRInputS6xD(78)(5) <= VNStageIntLLROutputS5xD(335)(1);
  CNStageIntLLRInputS6xD(170)(5) <= VNStageIntLLROutputS5xD(335)(2);
  CNStageIntLLRInputS6xD(189)(5) <= VNStageIntLLROutputS5xD(335)(3);
  CNStageIntLLRInputS6xD(274)(5) <= VNStageIntLLROutputS5xD(335)(4);
  CNStageIntLLRInputS6xD(291)(5) <= VNStageIntLLROutputS5xD(335)(5);
  CNStageIntLLRInputS6xD(343)(5) <= VNStageIntLLROutputS5xD(335)(6);
  CNStageIntLLRInputS6xD(38)(5) <= VNStageIntLLROutputS5xD(336)(0);
  CNStageIntLLRInputS6xD(104)(5) <= VNStageIntLLROutputS5xD(336)(1);
  CNStageIntLLRInputS6xD(121)(5) <= VNStageIntLLROutputS5xD(336)(2);
  CNStageIntLLRInputS6xD(267)(5) <= VNStageIntLLROutputS5xD(336)(3);
  CNStageIntLLRInputS6xD(332)(5) <= VNStageIntLLROutputS5xD(336)(4);
  CNStageIntLLRInputS6xD(344)(5) <= VNStageIntLLROutputS5xD(336)(5);
  CNStageIntLLRInputS6xD(37)(5) <= VNStageIntLLROutputS5xD(337)(0);
  CNStageIntLLRInputS6xD(93)(5) <= VNStageIntLLROutputS5xD(337)(1);
  CNStageIntLLRInputS6xD(115)(5) <= VNStageIntLLROutputS5xD(337)(2);
  CNStageIntLLRInputS6xD(183)(5) <= VNStageIntLLROutputS5xD(337)(3);
  CNStageIntLLRInputS6xD(253)(5) <= VNStageIntLLROutputS5xD(337)(4);
  CNStageIntLLRInputS6xD(290)(5) <= VNStageIntLLROutputS5xD(337)(5);
  CNStageIntLLRInputS6xD(379)(5) <= VNStageIntLLROutputS5xD(337)(6);
  CNStageIntLLRInputS6xD(36)(5) <= VNStageIntLLROutputS5xD(338)(0);
  CNStageIntLLRInputS6xD(80)(5) <= VNStageIntLLROutputS5xD(338)(1);
  CNStageIntLLRInputS6xD(155)(5) <= VNStageIntLLROutputS5xD(338)(2);
  CNStageIntLLRInputS6xD(190)(5) <= VNStageIntLLROutputS5xD(338)(3);
  CNStageIntLLRInputS6xD(370)(5) <= VNStageIntLLROutputS5xD(338)(4);
  CNStageIntLLRInputS6xD(35)(5) <= VNStageIntLLROutputS5xD(339)(0);
  CNStageIntLLRInputS6xD(96)(5) <= VNStageIntLLROutputS5xD(339)(1);
  CNStageIntLLRInputS6xD(163)(5) <= VNStageIntLLROutputS5xD(339)(2);
  CNStageIntLLRInputS6xD(216)(5) <= VNStageIntLLROutputS5xD(339)(3);
  CNStageIntLLRInputS6xD(247)(5) <= VNStageIntLLROutputS5xD(339)(4);
  CNStageIntLLRInputS6xD(322)(5) <= VNStageIntLLROutputS5xD(339)(5);
  CNStageIntLLRInputS6xD(34)(5) <= VNStageIntLLROutputS5xD(340)(0);
  CNStageIntLLRInputS6xD(58)(5) <= VNStageIntLLROutputS5xD(340)(1);
  CNStageIntLLRInputS6xD(127)(5) <= VNStageIntLLROutputS5xD(340)(2);
  CNStageIntLLRInputS6xD(178)(5) <= VNStageIntLLROutputS5xD(340)(3);
  CNStageIntLLRInputS6xD(245)(5) <= VNStageIntLLROutputS5xD(340)(4);
  CNStageIntLLRInputS6xD(334)(5) <= VNStageIntLLROutputS5xD(340)(5);
  CNStageIntLLRInputS6xD(33)(5) <= VNStageIntLLROutputS5xD(341)(0);
  CNStageIntLLRInputS6xD(68)(5) <= VNStageIntLLROutputS5xD(341)(1);
  CNStageIntLLRInputS6xD(125)(5) <= VNStageIntLLROutputS5xD(341)(2);
  CNStageIntLLRInputS6xD(204)(5) <= VNStageIntLLROutputS5xD(341)(3);
  CNStageIntLLRInputS6xD(258)(5) <= VNStageIntLLROutputS5xD(341)(4);
  CNStageIntLLRInputS6xD(296)(5) <= VNStageIntLLROutputS5xD(341)(5);
  CNStageIntLLRInputS6xD(32)(5) <= VNStageIntLLROutputS5xD(342)(0);
  CNStageIntLLRInputS6xD(63)(5) <= VNStageIntLLROutputS5xD(342)(1);
  CNStageIntLLRInputS6xD(161)(5) <= VNStageIntLLROutputS5xD(342)(2);
  CNStageIntLLRInputS6xD(251)(5) <= VNStageIntLLROutputS5xD(342)(3);
  CNStageIntLLRInputS6xD(294)(5) <= VNStageIntLLROutputS5xD(342)(4);
  CNStageIntLLRInputS6xD(31)(5) <= VNStageIntLLROutputS5xD(343)(0);
  CNStageIntLLRInputS6xD(69)(5) <= VNStageIntLLROutputS5xD(343)(1);
  CNStageIntLLRInputS6xD(140)(5) <= VNStageIntLLROutputS5xD(343)(2);
  CNStageIntLLRInputS6xD(206)(5) <= VNStageIntLLROutputS5xD(343)(3);
  CNStageIntLLRInputS6xD(228)(5) <= VNStageIntLLROutputS5xD(343)(4);
  CNStageIntLLRInputS6xD(327)(5) <= VNStageIntLLROutputS5xD(343)(5);
  CNStageIntLLRInputS6xD(30)(5) <= VNStageIntLLROutputS5xD(344)(0);
  CNStageIntLLRInputS6xD(57)(5) <= VNStageIntLLROutputS5xD(344)(1);
  CNStageIntLLRInputS6xD(143)(5) <= VNStageIntLLROutputS5xD(344)(2);
  CNStageIntLLRInputS6xD(218)(5) <= VNStageIntLLROutputS5xD(344)(3);
  CNStageIntLLRInputS6xD(238)(5) <= VNStageIntLLROutputS5xD(344)(4);
  CNStageIntLLRInputS6xD(307)(5) <= VNStageIntLLROutputS5xD(344)(5);
  CNStageIntLLRInputS6xD(367)(5) <= VNStageIntLLROutputS5xD(344)(6);
  CNStageIntLLRInputS6xD(29)(5) <= VNStageIntLLROutputS5xD(345)(0);
  CNStageIntLLRInputS6xD(83)(5) <= VNStageIntLLROutputS5xD(345)(1);
  CNStageIntLLRInputS6xD(128)(5) <= VNStageIntLLROutputS5xD(345)(2);
  CNStageIntLLRInputS6xD(232)(5) <= VNStageIntLLROutputS5xD(345)(3);
  CNStageIntLLRInputS6xD(309)(5) <= VNStageIntLLROutputS5xD(345)(4);
  CNStageIntLLRInputS6xD(375)(5) <= VNStageIntLLROutputS5xD(345)(5);
  CNStageIntLLRInputS6xD(28)(5) <= VNStageIntLLROutputS5xD(346)(0);
  CNStageIntLLRInputS6xD(89)(5) <= VNStageIntLLROutputS5xD(346)(1);
  CNStageIntLLRInputS6xD(162)(5) <= VNStageIntLLROutputS5xD(346)(2);
  CNStageIntLLRInputS6xD(181)(5) <= VNStageIntLLROutputS5xD(346)(3);
  CNStageIntLLRInputS6xD(235)(5) <= VNStageIntLLROutputS5xD(346)(4);
  CNStageIntLLRInputS6xD(297)(5) <= VNStageIntLLROutputS5xD(346)(5);
  CNStageIntLLRInputS6xD(339)(5) <= VNStageIntLLROutputS5xD(346)(6);
  CNStageIntLLRInputS6xD(27)(5) <= VNStageIntLLROutputS5xD(347)(0);
  CNStageIntLLRInputS6xD(73)(5) <= VNStageIntLLROutputS5xD(347)(1);
  CNStageIntLLRInputS6xD(124)(5) <= VNStageIntLLROutputS5xD(347)(2);
  CNStageIntLLRInputS6xD(199)(5) <= VNStageIntLLROutputS5xD(347)(3);
  CNStageIntLLRInputS6xD(225)(5) <= VNStageIntLLROutputS5xD(347)(4);
  CNStageIntLLRInputS6xD(328)(5) <= VNStageIntLLROutputS5xD(347)(5);
  CNStageIntLLRInputS6xD(337)(5) <= VNStageIntLLROutputS5xD(347)(6);
  CNStageIntLLRInputS6xD(26)(5) <= VNStageIntLLROutputS5xD(348)(0);
  CNStageIntLLRInputS6xD(75)(5) <= VNStageIntLLROutputS5xD(348)(1);
  CNStageIntLLRInputS6xD(152)(5) <= VNStageIntLLROutputS5xD(348)(2);
  CNStageIntLLRInputS6xD(200)(5) <= VNStageIntLLROutputS5xD(348)(3);
  CNStageIntLLRInputS6xD(259)(5) <= VNStageIntLLROutputS5xD(348)(4);
  CNStageIntLLRInputS6xD(293)(5) <= VNStageIntLLROutputS5xD(348)(5);
  CNStageIntLLRInputS6xD(373)(5) <= VNStageIntLLROutputS5xD(348)(6);
  CNStageIntLLRInputS6xD(25)(5) <= VNStageIntLLROutputS5xD(349)(0);
  CNStageIntLLRInputS6xD(99)(5) <= VNStageIntLLROutputS5xD(349)(1);
  CNStageIntLLRInputS6xD(180)(5) <= VNStageIntLLROutputS5xD(349)(2);
  CNStageIntLLRInputS6xD(244)(5) <= VNStageIntLLROutputS5xD(349)(3);
  CNStageIntLLRInputS6xD(319)(5) <= VNStageIntLLROutputS5xD(349)(4);
  CNStageIntLLRInputS6xD(352)(5) <= VNStageIntLLROutputS5xD(349)(5);
  CNStageIntLLRInputS6xD(24)(5) <= VNStageIntLLROutputS5xD(350)(0);
  CNStageIntLLRInputS6xD(81)(5) <= VNStageIntLLROutputS5xD(350)(1);
  CNStageIntLLRInputS6xD(164)(5) <= VNStageIntLLROutputS5xD(350)(2);
  CNStageIntLLRInputS6xD(171)(5) <= VNStageIntLLROutputS5xD(350)(3);
  CNStageIntLLRInputS6xD(254)(5) <= VNStageIntLLROutputS5xD(350)(4);
  CNStageIntLLRInputS6xD(303)(5) <= VNStageIntLLROutputS5xD(350)(5);
  CNStageIntLLRInputS6xD(23)(5) <= VNStageIntLLROutputS5xD(351)(0);
  CNStageIntLLRInputS6xD(154)(5) <= VNStageIntLLROutputS5xD(351)(1);
  CNStageIntLLRInputS6xD(188)(5) <= VNStageIntLLROutputS5xD(351)(2);
  CNStageIntLLRInputS6xD(266)(5) <= VNStageIntLLROutputS5xD(351)(3);
  CNStageIntLLRInputS6xD(329)(5) <= VNStageIntLLROutputS5xD(351)(4);
  CNStageIntLLRInputS6xD(340)(5) <= VNStageIntLLROutputS5xD(351)(5);
  CNStageIntLLRInputS6xD(22)(5) <= VNStageIntLLROutputS5xD(352)(0);
  CNStageIntLLRInputS6xD(100)(5) <= VNStageIntLLROutputS5xD(352)(1);
  CNStageIntLLRInputS6xD(141)(5) <= VNStageIntLLROutputS5xD(352)(2);
  CNStageIntLLRInputS6xD(192)(5) <= VNStageIntLLROutputS5xD(352)(3);
  CNStageIntLLRInputS6xD(239)(5) <= VNStageIntLLROutputS5xD(352)(4);
  CNStageIntLLRInputS6xD(321)(5) <= VNStageIntLLROutputS5xD(352)(5);
  CNStageIntLLRInputS6xD(374)(5) <= VNStageIntLLROutputS5xD(352)(6);
  CNStageIntLLRInputS6xD(21)(5) <= VNStageIntLLROutputS5xD(353)(0);
  CNStageIntLLRInputS6xD(74)(5) <= VNStageIntLLROutputS5xD(353)(1);
  CNStageIntLLRInputS6xD(160)(5) <= VNStageIntLLROutputS5xD(353)(2);
  CNStageIntLLRInputS6xD(224)(5) <= VNStageIntLLROutputS5xD(353)(3);
  CNStageIntLLRInputS6xD(227)(5) <= VNStageIntLLROutputS5xD(353)(4);
  CNStageIntLLRInputS6xD(336)(5) <= VNStageIntLLROutputS5xD(353)(5);
  CNStageIntLLRInputS6xD(20)(5) <= VNStageIntLLROutputS5xD(354)(0);
  CNStageIntLLRInputS6xD(88)(5) <= VNStageIntLLROutputS5xD(354)(1);
  CNStageIntLLRInputS6xD(133)(5) <= VNStageIntLLROutputS5xD(354)(2);
  CNStageIntLLRInputS6xD(191)(5) <= VNStageIntLLROutputS5xD(354)(3);
  CNStageIntLLRInputS6xD(326)(5) <= VNStageIntLLROutputS5xD(354)(4);
  CNStageIntLLRInputS6xD(364)(5) <= VNStageIntLLROutputS5xD(354)(5);
  CNStageIntLLRInputS6xD(19)(5) <= VNStageIntLLROutputS5xD(355)(0);
  CNStageIntLLRInputS6xD(59)(5) <= VNStageIntLLROutputS5xD(355)(1);
  CNStageIntLLRInputS6xD(130)(5) <= VNStageIntLLROutputS5xD(355)(2);
  CNStageIntLLRInputS6xD(186)(5) <= VNStageIntLLROutputS5xD(355)(3);
  CNStageIntLLRInputS6xD(230)(5) <= VNStageIntLLROutputS5xD(355)(4);
  CNStageIntLLRInputS6xD(300)(5) <= VNStageIntLLROutputS5xD(355)(5);
  CNStageIntLLRInputS6xD(349)(5) <= VNStageIntLLROutputS5xD(355)(6);
  CNStageIntLLRInputS6xD(18)(5) <= VNStageIntLLROutputS5xD(356)(0);
  CNStageIntLLRInputS6xD(95)(5) <= VNStageIntLLROutputS5xD(356)(1);
  CNStageIntLLRInputS6xD(146)(5) <= VNStageIntLLROutputS5xD(356)(2);
  CNStageIntLLRInputS6xD(222)(5) <= VNStageIntLLROutputS5xD(356)(3);
  CNStageIntLLRInputS6xD(299)(5) <= VNStageIntLLROutputS5xD(356)(4);
  CNStageIntLLRInputS6xD(376)(5) <= VNStageIntLLROutputS5xD(356)(5);
  CNStageIntLLRInputS6xD(17)(5) <= VNStageIntLLROutputS5xD(357)(0);
  CNStageIntLLRInputS6xD(61)(5) <= VNStageIntLLROutputS5xD(357)(1);
  CNStageIntLLRInputS6xD(138)(5) <= VNStageIntLLROutputS5xD(357)(2);
  CNStageIntLLRInputS6xD(176)(5) <= VNStageIntLLROutputS5xD(357)(3);
  CNStageIntLLRInputS6xD(256)(5) <= VNStageIntLLROutputS5xD(357)(4);
  CNStageIntLLRInputS6xD(312)(5) <= VNStageIntLLROutputS5xD(357)(5);
  CNStageIntLLRInputS6xD(366)(5) <= VNStageIntLLROutputS5xD(357)(6);
  CNStageIntLLRInputS6xD(16)(5) <= VNStageIntLLROutputS5xD(358)(0);
  CNStageIntLLRInputS6xD(76)(5) <= VNStageIntLLROutputS5xD(358)(1);
  CNStageIntLLRInputS6xD(112)(5) <= VNStageIntLLROutputS5xD(358)(2);
  CNStageIntLLRInputS6xD(252)(5) <= VNStageIntLLROutputS5xD(358)(3);
  CNStageIntLLRInputS6xD(305)(5) <= VNStageIntLLROutputS5xD(358)(4);
  CNStageIntLLRInputS6xD(353)(5) <= VNStageIntLLROutputS5xD(358)(5);
  CNStageIntLLRInputS6xD(15)(5) <= VNStageIntLLROutputS5xD(359)(0);
  CNStageIntLLRInputS6xD(72)(5) <= VNStageIntLLROutputS5xD(359)(1);
  CNStageIntLLRInputS6xD(122)(5) <= VNStageIntLLROutputS5xD(359)(2);
  CNStageIntLLRInputS6xD(195)(5) <= VNStageIntLLROutputS5xD(359)(3);
  CNStageIntLLRInputS6xD(257)(5) <= VNStageIntLLROutputS5xD(359)(4);
  CNStageIntLLRInputS6xD(283)(5) <= VNStageIntLLROutputS5xD(359)(5);
  CNStageIntLLRInputS6xD(372)(5) <= VNStageIntLLROutputS5xD(359)(6);
  CNStageIntLLRInputS6xD(14)(5) <= VNStageIntLLROutputS5xD(360)(0);
  CNStageIntLLRInputS6xD(91)(5) <= VNStageIntLLROutputS5xD(360)(1);
  CNStageIntLLRInputS6xD(116)(5) <= VNStageIntLLROutputS5xD(360)(2);
  CNStageIntLLRInputS6xD(174)(5) <= VNStageIntLLROutputS5xD(360)(3);
  CNStageIntLLRInputS6xD(248)(5) <= VNStageIntLLROutputS5xD(360)(4);
  CNStageIntLLRInputS6xD(292)(5) <= VNStageIntLLROutputS5xD(360)(5);
  CNStageIntLLRInputS6xD(345)(5) <= VNStageIntLLROutputS5xD(360)(6);
  CNStageIntLLRInputS6xD(13)(5) <= VNStageIntLLROutputS5xD(361)(0);
  CNStageIntLLRInputS6xD(54)(5) <= VNStageIntLLROutputS5xD(361)(1);
  CNStageIntLLRInputS6xD(120)(5) <= VNStageIntLLROutputS5xD(361)(2);
  CNStageIntLLRInputS6xD(207)(5) <= VNStageIntLLROutputS5xD(361)(3);
  CNStageIntLLRInputS6xD(271)(5) <= VNStageIntLLROutputS5xD(361)(4);
  CNStageIntLLRInputS6xD(285)(5) <= VNStageIntLLROutputS5xD(361)(5);
  CNStageIntLLRInputS6xD(342)(5) <= VNStageIntLLROutputS5xD(361)(6);
  CNStageIntLLRInputS6xD(12)(5) <= VNStageIntLLROutputS5xD(362)(0);
  CNStageIntLLRInputS6xD(55)(5) <= VNStageIntLLROutputS5xD(362)(1);
  CNStageIntLLRInputS6xD(169)(5) <= VNStageIntLLROutputS5xD(362)(2);
  CNStageIntLLRInputS6xD(210)(5) <= VNStageIntLLROutputS5xD(362)(3);
  CNStageIntLLRInputS6xD(276)(5) <= VNStageIntLLROutputS5xD(362)(4);
  CNStageIntLLRInputS6xD(289)(5) <= VNStageIntLLROutputS5xD(362)(5);
  CNStageIntLLRInputS6xD(357)(5) <= VNStageIntLLROutputS5xD(362)(6);
  CNStageIntLLRInputS6xD(90)(5) <= VNStageIntLLROutputS5xD(363)(0);
  CNStageIntLLRInputS6xD(147)(5) <= VNStageIntLLROutputS5xD(363)(1);
  CNStageIntLLRInputS6xD(197)(5) <= VNStageIntLLROutputS5xD(363)(2);
  CNStageIntLLRInputS6xD(261)(5) <= VNStageIntLLROutputS5xD(363)(3);
  CNStageIntLLRInputS6xD(281)(5) <= VNStageIntLLROutputS5xD(363)(4);
  CNStageIntLLRInputS6xD(11)(5) <= VNStageIntLLROutputS5xD(364)(0);
  CNStageIntLLRInputS6xD(82)(5) <= VNStageIntLLROutputS5xD(364)(1);
  CNStageIntLLRInputS6xD(129)(5) <= VNStageIntLLROutputS5xD(364)(2);
  CNStageIntLLRInputS6xD(175)(5) <= VNStageIntLLROutputS5xD(364)(3);
  CNStageIntLLRInputS6xD(263)(5) <= VNStageIntLLROutputS5xD(364)(4);
  CNStageIntLLRInputS6xD(313)(5) <= VNStageIntLLROutputS5xD(364)(5);
  CNStageIntLLRInputS6xD(10)(5) <= VNStageIntLLROutputS5xD(365)(0);
  CNStageIntLLRInputS6xD(98)(5) <= VNStageIntLLROutputS5xD(365)(1);
  CNStageIntLLRInputS6xD(142)(5) <= VNStageIntLLROutputS5xD(365)(2);
  CNStageIntLLRInputS6xD(194)(5) <= VNStageIntLLROutputS5xD(365)(3);
  CNStageIntLLRInputS6xD(234)(5) <= VNStageIntLLROutputS5xD(365)(4);
  CNStageIntLLRInputS6xD(298)(5) <= VNStageIntLLROutputS5xD(365)(5);
  CNStageIntLLRInputS6xD(9)(5) <= VNStageIntLLROutputS5xD(366)(0);
  CNStageIntLLRInputS6xD(102)(5) <= VNStageIntLLROutputS5xD(366)(1);
  CNStageIntLLRInputS6xD(153)(5) <= VNStageIntLLROutputS5xD(366)(2);
  CNStageIntLLRInputS6xD(219)(5) <= VNStageIntLLROutputS5xD(366)(3);
  CNStageIntLLRInputS6xD(269)(5) <= VNStageIntLLROutputS5xD(366)(4);
  CNStageIntLLRInputS6xD(308)(5) <= VNStageIntLLROutputS5xD(366)(5);
  CNStageIntLLRInputS6xD(8)(5) <= VNStageIntLLROutputS5xD(367)(0);
  CNStageIntLLRInputS6xD(110)(5) <= VNStageIntLLROutputS5xD(367)(1);
  CNStageIntLLRInputS6xD(123)(5) <= VNStageIntLLROutputS5xD(367)(2);
  CNStageIntLLRInputS6xD(205)(5) <= VNStageIntLLROutputS5xD(367)(3);
  CNStageIntLLRInputS6xD(226)(5) <= VNStageIntLLROutputS5xD(367)(4);
  CNStageIntLLRInputS6xD(320)(5) <= VNStageIntLLROutputS5xD(367)(5);
  CNStageIntLLRInputS6xD(333)(5) <= VNStageIntLLROutputS5xD(367)(6);
  CNStageIntLLRInputS6xD(7)(5) <= VNStageIntLLROutputS5xD(368)(0);
  CNStageIntLLRInputS6xD(177)(5) <= VNStageIntLLROutputS5xD(368)(1);
  CNStageIntLLRInputS6xD(381)(5) <= VNStageIntLLROutputS5xD(368)(2);
  CNStageIntLLRInputS6xD(6)(5) <= VNStageIntLLROutputS5xD(369)(0);
  CNStageIntLLRInputS6xD(156)(5) <= VNStageIntLLROutputS5xD(369)(1);
  CNStageIntLLRInputS6xD(221)(5) <= VNStageIntLLROutputS5xD(369)(2);
  CNStageIntLLRInputS6xD(262)(5) <= VNStageIntLLROutputS5xD(369)(3);
  CNStageIntLLRInputS6xD(358)(5) <= VNStageIntLLROutputS5xD(369)(4);
  CNStageIntLLRInputS6xD(5)(5) <= VNStageIntLLROutputS5xD(370)(0);
  CNStageIntLLRInputS6xD(114)(5) <= VNStageIntLLROutputS5xD(370)(1);
  CNStageIntLLRInputS6xD(208)(5) <= VNStageIntLLROutputS5xD(370)(2);
  CNStageIntLLRInputS6xD(275)(5) <= VNStageIntLLROutputS5xD(370)(3);
  CNStageIntLLRInputS6xD(341)(5) <= VNStageIntLLROutputS5xD(370)(4);
  CNStageIntLLRInputS6xD(4)(5) <= VNStageIntLLROutputS5xD(371)(0);
  CNStageIntLLRInputS6xD(135)(5) <= VNStageIntLLROutputS5xD(371)(1);
  CNStageIntLLRInputS6xD(173)(5) <= VNStageIntLLROutputS5xD(371)(2);
  CNStageIntLLRInputS6xD(249)(5) <= VNStageIntLLROutputS5xD(371)(3);
  CNStageIntLLRInputS6xD(354)(5) <= VNStageIntLLROutputS5xD(371)(4);
  CNStageIntLLRInputS6xD(106)(5) <= VNStageIntLLROutputS5xD(372)(0);
  CNStageIntLLRInputS6xD(144)(5) <= VNStageIntLLROutputS5xD(372)(1);
  CNStageIntLLRInputS6xD(201)(5) <= VNStageIntLLROutputS5xD(372)(2);
  CNStageIntLLRInputS6xD(229)(5) <= VNStageIntLLROutputS5xD(372)(3);
  CNStageIntLLRInputS6xD(301)(5) <= VNStageIntLLROutputS5xD(372)(4);
  CNStageIntLLRInputS6xD(365)(5) <= VNStageIntLLROutputS5xD(372)(5);
  CNStageIntLLRInputS6xD(3)(5) <= VNStageIntLLROutputS5xD(373)(0);
  CNStageIntLLRInputS6xD(139)(5) <= VNStageIntLLROutputS5xD(373)(1);
  CNStageIntLLRInputS6xD(250)(5) <= VNStageIntLLROutputS5xD(373)(2);
  CNStageIntLLRInputS6xD(310)(5) <= VNStageIntLLROutputS5xD(373)(3);
  CNStageIntLLRInputS6xD(335)(5) <= VNStageIntLLROutputS5xD(373)(4);
  CNStageIntLLRInputS6xD(2)(5) <= VNStageIntLLROutputS5xD(374)(0);
  CNStageIntLLRInputS6xD(85)(5) <= VNStageIntLLROutputS5xD(374)(1);
  CNStageIntLLRInputS6xD(145)(5) <= VNStageIntLLROutputS5xD(374)(2);
  CNStageIntLLRInputS6xD(213)(5) <= VNStageIntLLROutputS5xD(374)(3);
  CNStageIntLLRInputS6xD(264)(5) <= VNStageIntLLROutputS5xD(374)(4);
  CNStageIntLLRInputS6xD(306)(5) <= VNStageIntLLROutputS5xD(374)(5);
  CNStageIntLLRInputS6xD(383)(5) <= VNStageIntLLROutputS5xD(374)(6);
  CNStageIntLLRInputS6xD(1)(5) <= VNStageIntLLROutputS5xD(375)(0);
  CNStageIntLLRInputS6xD(64)(5) <= VNStageIntLLROutputS5xD(375)(1);
  CNStageIntLLRInputS6xD(134)(5) <= VNStageIntLLROutputS5xD(375)(2);
  CNStageIntLLRInputS6xD(260)(5) <= VNStageIntLLROutputS5xD(375)(3);
  CNStageIntLLRInputS6xD(311)(5) <= VNStageIntLLROutputS5xD(375)(4);
  CNStageIntLLRInputS6xD(368)(5) <= VNStageIntLLROutputS5xD(375)(5);
  CNStageIntLLRInputS6xD(0)(5) <= VNStageIntLLROutputS5xD(376)(0);
  CNStageIntLLRInputS6xD(67)(5) <= VNStageIntLLROutputS5xD(376)(1);
  CNStageIntLLRInputS6xD(159)(5) <= VNStageIntLLROutputS5xD(376)(2);
  CNStageIntLLRInputS6xD(278)(5) <= VNStageIntLLROutputS5xD(376)(3);
  CNStageIntLLRInputS6xD(107)(5) <= VNStageIntLLROutputS5xD(377)(0);
  CNStageIntLLRInputS6xD(166)(5) <= VNStageIntLLROutputS5xD(377)(1);
  CNStageIntLLRInputS6xD(193)(5) <= VNStageIntLLROutputS5xD(377)(2);
  CNStageIntLLRInputS6xD(325)(5) <= VNStageIntLLROutputS5xD(377)(3);
  CNStageIntLLRInputS6xD(347)(5) <= VNStageIntLLROutputS5xD(377)(4);
  CNStageIntLLRInputS6xD(86)(5) <= VNStageIntLLROutputS5xD(378)(0);
  CNStageIntLLRInputS6xD(149)(5) <= VNStageIntLLROutputS5xD(378)(1);
  CNStageIntLLRInputS6xD(187)(5) <= VNStageIntLLROutputS5xD(378)(2);
  CNStageIntLLRInputS6xD(246)(5) <= VNStageIntLLROutputS5xD(378)(3);
  CNStageIntLLRInputS6xD(331)(5) <= VNStageIntLLROutputS5xD(378)(4);
  CNStageIntLLRInputS6xD(355)(5) <= VNStageIntLLROutputS5xD(378)(5);
  CNStageIntLLRInputS6xD(105)(5) <= VNStageIntLLROutputS5xD(379)(0);
  CNStageIntLLRInputS6xD(151)(5) <= VNStageIntLLROutputS5xD(379)(1);
  CNStageIntLLRInputS6xD(277)(5) <= VNStageIntLLROutputS5xD(379)(2);
  CNStageIntLLRInputS6xD(315)(5) <= VNStageIntLLROutputS5xD(379)(3);
  CNStageIntLLRInputS6xD(351)(5) <= VNStageIntLLROutputS5xD(379)(4);
  CNStageIntLLRInputS6xD(77)(5) <= VNStageIntLLROutputS5xD(380)(0);
  CNStageIntLLRInputS6xD(118)(5) <= VNStageIntLLROutputS5xD(380)(1);
  CNStageIntLLRInputS6xD(182)(5) <= VNStageIntLLROutputS5xD(380)(2);
  CNStageIntLLRInputS6xD(270)(5) <= VNStageIntLLROutputS5xD(380)(3);
  CNStageIntLLRInputS6xD(317)(5) <= VNStageIntLLROutputS5xD(380)(4);
  CNStageIntLLRInputS6xD(356)(5) <= VNStageIntLLROutputS5xD(380)(5);
  CNStageIntLLRInputS6xD(60)(5) <= VNStageIntLLROutputS5xD(381)(0);
  CNStageIntLLRInputS6xD(157)(5) <= VNStageIntLLROutputS5xD(381)(1);
  CNStageIntLLRInputS6xD(214)(5) <= VNStageIntLLROutputS5xD(381)(2);
  CNStageIntLLRInputS6xD(233)(5) <= VNStageIntLLROutputS5xD(381)(3);
  CNStageIntLLRInputS6xD(287)(5) <= VNStageIntLLROutputS5xD(381)(4);
  CNStageIntLLRInputS6xD(346)(5) <= VNStageIntLLROutputS5xD(381)(5);
  CNStageIntLLRInputS6xD(87)(5) <= VNStageIntLLROutputS5xD(382)(0);
  CNStageIntLLRInputS6xD(111)(5) <= VNStageIntLLROutputS5xD(382)(1);
  CNStageIntLLRInputS6xD(198)(5) <= VNStageIntLLROutputS5xD(382)(2);
  CNStageIntLLRInputS6xD(237)(5) <= VNStageIntLLROutputS5xD(382)(3);
  CNStageIntLLRInputS6xD(323)(5) <= VNStageIntLLROutputS5xD(382)(4);
  CNStageIntLLRInputS6xD(371)(5) <= VNStageIntLLROutputS5xD(382)(5);
  CNStageIntLLRInputS6xD(52)(5) <= VNStageIntLLROutputS5xD(383)(0);
  CNStageIntLLRInputS6xD(79)(5) <= VNStageIntLLROutputS5xD(383)(1);
  CNStageIntLLRInputS6xD(119)(5) <= VNStageIntLLROutputS5xD(383)(2);
  CNStageIntLLRInputS6xD(209)(5) <= VNStageIntLLROutputS5xD(383)(3);
  CNStageIntLLRInputS6xD(279)(5) <= VNStageIntLLROutputS5xD(383)(4);
  CNStageIntLLRInputS6xD(282)(5) <= VNStageIntLLROutputS5xD(383)(5);
  CNStageIntLLRInputS6xD(378)(5) <= VNStageIntLLROutputS5xD(383)(6);

  -- Variable Nodes (Iteration 6)
  VNStageIntLLRInputS6xD(56)(0) <= CNStageIntLLROutputS6xD(0)(0);
  VNStageIntLLRInputS6xD(120)(0) <= CNStageIntLLROutputS6xD(0)(1);
  VNStageIntLLRInputS6xD(184)(0) <= CNStageIntLLROutputS6xD(0)(2);
  VNStageIntLLRInputS6xD(248)(0) <= CNStageIntLLROutputS6xD(0)(3);
  VNStageIntLLRInputS6xD(312)(0) <= CNStageIntLLROutputS6xD(0)(4);
  VNStageIntLLRInputS6xD(376)(0) <= CNStageIntLLROutputS6xD(0)(5);
  VNStageIntLLRInputS6xD(55)(0) <= CNStageIntLLROutputS6xD(1)(0);
  VNStageIntLLRInputS6xD(119)(0) <= CNStageIntLLROutputS6xD(1)(1);
  VNStageIntLLRInputS6xD(183)(0) <= CNStageIntLLROutputS6xD(1)(2);
  VNStageIntLLRInputS6xD(247)(0) <= CNStageIntLLROutputS6xD(1)(3);
  VNStageIntLLRInputS6xD(311)(0) <= CNStageIntLLROutputS6xD(1)(4);
  VNStageIntLLRInputS6xD(375)(0) <= CNStageIntLLROutputS6xD(1)(5);
  VNStageIntLLRInputS6xD(54)(0) <= CNStageIntLLROutputS6xD(2)(0);
  VNStageIntLLRInputS6xD(118)(0) <= CNStageIntLLROutputS6xD(2)(1);
  VNStageIntLLRInputS6xD(182)(0) <= CNStageIntLLROutputS6xD(2)(2);
  VNStageIntLLRInputS6xD(246)(0) <= CNStageIntLLROutputS6xD(2)(3);
  VNStageIntLLRInputS6xD(310)(0) <= CNStageIntLLROutputS6xD(2)(4);
  VNStageIntLLRInputS6xD(374)(0) <= CNStageIntLLROutputS6xD(2)(5);
  VNStageIntLLRInputS6xD(53)(0) <= CNStageIntLLROutputS6xD(3)(0);
  VNStageIntLLRInputS6xD(117)(0) <= CNStageIntLLROutputS6xD(3)(1);
  VNStageIntLLRInputS6xD(181)(0) <= CNStageIntLLROutputS6xD(3)(2);
  VNStageIntLLRInputS6xD(245)(0) <= CNStageIntLLROutputS6xD(3)(3);
  VNStageIntLLRInputS6xD(309)(0) <= CNStageIntLLROutputS6xD(3)(4);
  VNStageIntLLRInputS6xD(373)(0) <= CNStageIntLLROutputS6xD(3)(5);
  VNStageIntLLRInputS6xD(51)(0) <= CNStageIntLLROutputS6xD(4)(0);
  VNStageIntLLRInputS6xD(115)(0) <= CNStageIntLLROutputS6xD(4)(1);
  VNStageIntLLRInputS6xD(179)(0) <= CNStageIntLLROutputS6xD(4)(2);
  VNStageIntLLRInputS6xD(243)(0) <= CNStageIntLLROutputS6xD(4)(3);
  VNStageIntLLRInputS6xD(307)(0) <= CNStageIntLLROutputS6xD(4)(4);
  VNStageIntLLRInputS6xD(371)(0) <= CNStageIntLLROutputS6xD(4)(5);
  VNStageIntLLRInputS6xD(50)(0) <= CNStageIntLLROutputS6xD(5)(0);
  VNStageIntLLRInputS6xD(114)(0) <= CNStageIntLLROutputS6xD(5)(1);
  VNStageIntLLRInputS6xD(178)(0) <= CNStageIntLLROutputS6xD(5)(2);
  VNStageIntLLRInputS6xD(242)(0) <= CNStageIntLLROutputS6xD(5)(3);
  VNStageIntLLRInputS6xD(306)(0) <= CNStageIntLLROutputS6xD(5)(4);
  VNStageIntLLRInputS6xD(370)(0) <= CNStageIntLLROutputS6xD(5)(5);
  VNStageIntLLRInputS6xD(49)(0) <= CNStageIntLLROutputS6xD(6)(0);
  VNStageIntLLRInputS6xD(113)(0) <= CNStageIntLLROutputS6xD(6)(1);
  VNStageIntLLRInputS6xD(177)(0) <= CNStageIntLLROutputS6xD(6)(2);
  VNStageIntLLRInputS6xD(241)(0) <= CNStageIntLLROutputS6xD(6)(3);
  VNStageIntLLRInputS6xD(305)(0) <= CNStageIntLLROutputS6xD(6)(4);
  VNStageIntLLRInputS6xD(369)(0) <= CNStageIntLLROutputS6xD(6)(5);
  VNStageIntLLRInputS6xD(48)(0) <= CNStageIntLLROutputS6xD(7)(0);
  VNStageIntLLRInputS6xD(112)(0) <= CNStageIntLLROutputS6xD(7)(1);
  VNStageIntLLRInputS6xD(176)(0) <= CNStageIntLLROutputS6xD(7)(2);
  VNStageIntLLRInputS6xD(240)(0) <= CNStageIntLLROutputS6xD(7)(3);
  VNStageIntLLRInputS6xD(304)(0) <= CNStageIntLLROutputS6xD(7)(4);
  VNStageIntLLRInputS6xD(368)(0) <= CNStageIntLLROutputS6xD(7)(5);
  VNStageIntLLRInputS6xD(47)(0) <= CNStageIntLLROutputS6xD(8)(0);
  VNStageIntLLRInputS6xD(111)(0) <= CNStageIntLLROutputS6xD(8)(1);
  VNStageIntLLRInputS6xD(175)(0) <= CNStageIntLLROutputS6xD(8)(2);
  VNStageIntLLRInputS6xD(239)(0) <= CNStageIntLLROutputS6xD(8)(3);
  VNStageIntLLRInputS6xD(303)(0) <= CNStageIntLLROutputS6xD(8)(4);
  VNStageIntLLRInputS6xD(367)(0) <= CNStageIntLLROutputS6xD(8)(5);
  VNStageIntLLRInputS6xD(46)(0) <= CNStageIntLLROutputS6xD(9)(0);
  VNStageIntLLRInputS6xD(110)(0) <= CNStageIntLLROutputS6xD(9)(1);
  VNStageIntLLRInputS6xD(174)(0) <= CNStageIntLLROutputS6xD(9)(2);
  VNStageIntLLRInputS6xD(238)(0) <= CNStageIntLLROutputS6xD(9)(3);
  VNStageIntLLRInputS6xD(302)(0) <= CNStageIntLLROutputS6xD(9)(4);
  VNStageIntLLRInputS6xD(366)(0) <= CNStageIntLLROutputS6xD(9)(5);
  VNStageIntLLRInputS6xD(45)(0) <= CNStageIntLLROutputS6xD(10)(0);
  VNStageIntLLRInputS6xD(109)(0) <= CNStageIntLLROutputS6xD(10)(1);
  VNStageIntLLRInputS6xD(173)(0) <= CNStageIntLLROutputS6xD(10)(2);
  VNStageIntLLRInputS6xD(237)(0) <= CNStageIntLLROutputS6xD(10)(3);
  VNStageIntLLRInputS6xD(301)(0) <= CNStageIntLLROutputS6xD(10)(4);
  VNStageIntLLRInputS6xD(365)(0) <= CNStageIntLLROutputS6xD(10)(5);
  VNStageIntLLRInputS6xD(44)(0) <= CNStageIntLLROutputS6xD(11)(0);
  VNStageIntLLRInputS6xD(108)(0) <= CNStageIntLLROutputS6xD(11)(1);
  VNStageIntLLRInputS6xD(172)(0) <= CNStageIntLLROutputS6xD(11)(2);
  VNStageIntLLRInputS6xD(236)(0) <= CNStageIntLLROutputS6xD(11)(3);
  VNStageIntLLRInputS6xD(300)(0) <= CNStageIntLLROutputS6xD(11)(4);
  VNStageIntLLRInputS6xD(364)(0) <= CNStageIntLLROutputS6xD(11)(5);
  VNStageIntLLRInputS6xD(42)(0) <= CNStageIntLLROutputS6xD(12)(0);
  VNStageIntLLRInputS6xD(106)(0) <= CNStageIntLLROutputS6xD(12)(1);
  VNStageIntLLRInputS6xD(170)(0) <= CNStageIntLLROutputS6xD(12)(2);
  VNStageIntLLRInputS6xD(234)(0) <= CNStageIntLLROutputS6xD(12)(3);
  VNStageIntLLRInputS6xD(298)(0) <= CNStageIntLLROutputS6xD(12)(4);
  VNStageIntLLRInputS6xD(362)(0) <= CNStageIntLLROutputS6xD(12)(5);
  VNStageIntLLRInputS6xD(41)(0) <= CNStageIntLLROutputS6xD(13)(0);
  VNStageIntLLRInputS6xD(105)(0) <= CNStageIntLLROutputS6xD(13)(1);
  VNStageIntLLRInputS6xD(169)(0) <= CNStageIntLLROutputS6xD(13)(2);
  VNStageIntLLRInputS6xD(233)(0) <= CNStageIntLLROutputS6xD(13)(3);
  VNStageIntLLRInputS6xD(297)(0) <= CNStageIntLLROutputS6xD(13)(4);
  VNStageIntLLRInputS6xD(361)(0) <= CNStageIntLLROutputS6xD(13)(5);
  VNStageIntLLRInputS6xD(40)(0) <= CNStageIntLLROutputS6xD(14)(0);
  VNStageIntLLRInputS6xD(104)(0) <= CNStageIntLLROutputS6xD(14)(1);
  VNStageIntLLRInputS6xD(168)(0) <= CNStageIntLLROutputS6xD(14)(2);
  VNStageIntLLRInputS6xD(232)(0) <= CNStageIntLLROutputS6xD(14)(3);
  VNStageIntLLRInputS6xD(296)(0) <= CNStageIntLLROutputS6xD(14)(4);
  VNStageIntLLRInputS6xD(360)(0) <= CNStageIntLLROutputS6xD(14)(5);
  VNStageIntLLRInputS6xD(39)(0) <= CNStageIntLLROutputS6xD(15)(0);
  VNStageIntLLRInputS6xD(103)(0) <= CNStageIntLLROutputS6xD(15)(1);
  VNStageIntLLRInputS6xD(167)(0) <= CNStageIntLLROutputS6xD(15)(2);
  VNStageIntLLRInputS6xD(231)(0) <= CNStageIntLLROutputS6xD(15)(3);
  VNStageIntLLRInputS6xD(295)(0) <= CNStageIntLLROutputS6xD(15)(4);
  VNStageIntLLRInputS6xD(359)(0) <= CNStageIntLLROutputS6xD(15)(5);
  VNStageIntLLRInputS6xD(38)(0) <= CNStageIntLLROutputS6xD(16)(0);
  VNStageIntLLRInputS6xD(102)(0) <= CNStageIntLLROutputS6xD(16)(1);
  VNStageIntLLRInputS6xD(166)(0) <= CNStageIntLLROutputS6xD(16)(2);
  VNStageIntLLRInputS6xD(230)(0) <= CNStageIntLLROutputS6xD(16)(3);
  VNStageIntLLRInputS6xD(294)(0) <= CNStageIntLLROutputS6xD(16)(4);
  VNStageIntLLRInputS6xD(358)(0) <= CNStageIntLLROutputS6xD(16)(5);
  VNStageIntLLRInputS6xD(37)(0) <= CNStageIntLLROutputS6xD(17)(0);
  VNStageIntLLRInputS6xD(101)(0) <= CNStageIntLLROutputS6xD(17)(1);
  VNStageIntLLRInputS6xD(165)(0) <= CNStageIntLLROutputS6xD(17)(2);
  VNStageIntLLRInputS6xD(229)(0) <= CNStageIntLLROutputS6xD(17)(3);
  VNStageIntLLRInputS6xD(293)(0) <= CNStageIntLLROutputS6xD(17)(4);
  VNStageIntLLRInputS6xD(357)(0) <= CNStageIntLLROutputS6xD(17)(5);
  VNStageIntLLRInputS6xD(36)(0) <= CNStageIntLLROutputS6xD(18)(0);
  VNStageIntLLRInputS6xD(100)(0) <= CNStageIntLLROutputS6xD(18)(1);
  VNStageIntLLRInputS6xD(164)(0) <= CNStageIntLLROutputS6xD(18)(2);
  VNStageIntLLRInputS6xD(228)(0) <= CNStageIntLLROutputS6xD(18)(3);
  VNStageIntLLRInputS6xD(292)(0) <= CNStageIntLLROutputS6xD(18)(4);
  VNStageIntLLRInputS6xD(356)(0) <= CNStageIntLLROutputS6xD(18)(5);
  VNStageIntLLRInputS6xD(35)(0) <= CNStageIntLLROutputS6xD(19)(0);
  VNStageIntLLRInputS6xD(99)(0) <= CNStageIntLLROutputS6xD(19)(1);
  VNStageIntLLRInputS6xD(163)(0) <= CNStageIntLLROutputS6xD(19)(2);
  VNStageIntLLRInputS6xD(227)(0) <= CNStageIntLLROutputS6xD(19)(3);
  VNStageIntLLRInputS6xD(291)(0) <= CNStageIntLLROutputS6xD(19)(4);
  VNStageIntLLRInputS6xD(355)(0) <= CNStageIntLLROutputS6xD(19)(5);
  VNStageIntLLRInputS6xD(34)(0) <= CNStageIntLLROutputS6xD(20)(0);
  VNStageIntLLRInputS6xD(98)(0) <= CNStageIntLLROutputS6xD(20)(1);
  VNStageIntLLRInputS6xD(162)(0) <= CNStageIntLLROutputS6xD(20)(2);
  VNStageIntLLRInputS6xD(226)(0) <= CNStageIntLLROutputS6xD(20)(3);
  VNStageIntLLRInputS6xD(290)(0) <= CNStageIntLLROutputS6xD(20)(4);
  VNStageIntLLRInputS6xD(354)(0) <= CNStageIntLLROutputS6xD(20)(5);
  VNStageIntLLRInputS6xD(33)(0) <= CNStageIntLLROutputS6xD(21)(0);
  VNStageIntLLRInputS6xD(97)(0) <= CNStageIntLLROutputS6xD(21)(1);
  VNStageIntLLRInputS6xD(161)(0) <= CNStageIntLLROutputS6xD(21)(2);
  VNStageIntLLRInputS6xD(225)(0) <= CNStageIntLLROutputS6xD(21)(3);
  VNStageIntLLRInputS6xD(289)(0) <= CNStageIntLLROutputS6xD(21)(4);
  VNStageIntLLRInputS6xD(353)(0) <= CNStageIntLLROutputS6xD(21)(5);
  VNStageIntLLRInputS6xD(32)(0) <= CNStageIntLLROutputS6xD(22)(0);
  VNStageIntLLRInputS6xD(96)(0) <= CNStageIntLLROutputS6xD(22)(1);
  VNStageIntLLRInputS6xD(160)(0) <= CNStageIntLLROutputS6xD(22)(2);
  VNStageIntLLRInputS6xD(224)(0) <= CNStageIntLLROutputS6xD(22)(3);
  VNStageIntLLRInputS6xD(288)(0) <= CNStageIntLLROutputS6xD(22)(4);
  VNStageIntLLRInputS6xD(352)(0) <= CNStageIntLLROutputS6xD(22)(5);
  VNStageIntLLRInputS6xD(31)(0) <= CNStageIntLLROutputS6xD(23)(0);
  VNStageIntLLRInputS6xD(95)(0) <= CNStageIntLLROutputS6xD(23)(1);
  VNStageIntLLRInputS6xD(159)(0) <= CNStageIntLLROutputS6xD(23)(2);
  VNStageIntLLRInputS6xD(223)(0) <= CNStageIntLLROutputS6xD(23)(3);
  VNStageIntLLRInputS6xD(287)(0) <= CNStageIntLLROutputS6xD(23)(4);
  VNStageIntLLRInputS6xD(351)(0) <= CNStageIntLLROutputS6xD(23)(5);
  VNStageIntLLRInputS6xD(30)(0) <= CNStageIntLLROutputS6xD(24)(0);
  VNStageIntLLRInputS6xD(94)(0) <= CNStageIntLLROutputS6xD(24)(1);
  VNStageIntLLRInputS6xD(158)(0) <= CNStageIntLLROutputS6xD(24)(2);
  VNStageIntLLRInputS6xD(222)(0) <= CNStageIntLLROutputS6xD(24)(3);
  VNStageIntLLRInputS6xD(286)(0) <= CNStageIntLLROutputS6xD(24)(4);
  VNStageIntLLRInputS6xD(350)(0) <= CNStageIntLLROutputS6xD(24)(5);
  VNStageIntLLRInputS6xD(29)(0) <= CNStageIntLLROutputS6xD(25)(0);
  VNStageIntLLRInputS6xD(93)(0) <= CNStageIntLLROutputS6xD(25)(1);
  VNStageIntLLRInputS6xD(157)(0) <= CNStageIntLLROutputS6xD(25)(2);
  VNStageIntLLRInputS6xD(221)(0) <= CNStageIntLLROutputS6xD(25)(3);
  VNStageIntLLRInputS6xD(285)(0) <= CNStageIntLLROutputS6xD(25)(4);
  VNStageIntLLRInputS6xD(349)(0) <= CNStageIntLLROutputS6xD(25)(5);
  VNStageIntLLRInputS6xD(28)(0) <= CNStageIntLLROutputS6xD(26)(0);
  VNStageIntLLRInputS6xD(92)(0) <= CNStageIntLLROutputS6xD(26)(1);
  VNStageIntLLRInputS6xD(156)(0) <= CNStageIntLLROutputS6xD(26)(2);
  VNStageIntLLRInputS6xD(220)(0) <= CNStageIntLLROutputS6xD(26)(3);
  VNStageIntLLRInputS6xD(284)(0) <= CNStageIntLLROutputS6xD(26)(4);
  VNStageIntLLRInputS6xD(348)(0) <= CNStageIntLLROutputS6xD(26)(5);
  VNStageIntLLRInputS6xD(27)(0) <= CNStageIntLLROutputS6xD(27)(0);
  VNStageIntLLRInputS6xD(91)(0) <= CNStageIntLLROutputS6xD(27)(1);
  VNStageIntLLRInputS6xD(155)(0) <= CNStageIntLLROutputS6xD(27)(2);
  VNStageIntLLRInputS6xD(219)(0) <= CNStageIntLLROutputS6xD(27)(3);
  VNStageIntLLRInputS6xD(283)(0) <= CNStageIntLLROutputS6xD(27)(4);
  VNStageIntLLRInputS6xD(347)(0) <= CNStageIntLLROutputS6xD(27)(5);
  VNStageIntLLRInputS6xD(26)(0) <= CNStageIntLLROutputS6xD(28)(0);
  VNStageIntLLRInputS6xD(90)(0) <= CNStageIntLLROutputS6xD(28)(1);
  VNStageIntLLRInputS6xD(154)(0) <= CNStageIntLLROutputS6xD(28)(2);
  VNStageIntLLRInputS6xD(218)(0) <= CNStageIntLLROutputS6xD(28)(3);
  VNStageIntLLRInputS6xD(282)(0) <= CNStageIntLLROutputS6xD(28)(4);
  VNStageIntLLRInputS6xD(346)(0) <= CNStageIntLLROutputS6xD(28)(5);
  VNStageIntLLRInputS6xD(25)(0) <= CNStageIntLLROutputS6xD(29)(0);
  VNStageIntLLRInputS6xD(89)(0) <= CNStageIntLLROutputS6xD(29)(1);
  VNStageIntLLRInputS6xD(153)(0) <= CNStageIntLLROutputS6xD(29)(2);
  VNStageIntLLRInputS6xD(217)(0) <= CNStageIntLLROutputS6xD(29)(3);
  VNStageIntLLRInputS6xD(281)(0) <= CNStageIntLLROutputS6xD(29)(4);
  VNStageIntLLRInputS6xD(345)(0) <= CNStageIntLLROutputS6xD(29)(5);
  VNStageIntLLRInputS6xD(24)(0) <= CNStageIntLLROutputS6xD(30)(0);
  VNStageIntLLRInputS6xD(88)(0) <= CNStageIntLLROutputS6xD(30)(1);
  VNStageIntLLRInputS6xD(152)(0) <= CNStageIntLLROutputS6xD(30)(2);
  VNStageIntLLRInputS6xD(216)(0) <= CNStageIntLLROutputS6xD(30)(3);
  VNStageIntLLRInputS6xD(280)(0) <= CNStageIntLLROutputS6xD(30)(4);
  VNStageIntLLRInputS6xD(344)(0) <= CNStageIntLLROutputS6xD(30)(5);
  VNStageIntLLRInputS6xD(23)(0) <= CNStageIntLLROutputS6xD(31)(0);
  VNStageIntLLRInputS6xD(87)(0) <= CNStageIntLLROutputS6xD(31)(1);
  VNStageIntLLRInputS6xD(151)(0) <= CNStageIntLLROutputS6xD(31)(2);
  VNStageIntLLRInputS6xD(215)(0) <= CNStageIntLLROutputS6xD(31)(3);
  VNStageIntLLRInputS6xD(279)(0) <= CNStageIntLLROutputS6xD(31)(4);
  VNStageIntLLRInputS6xD(343)(0) <= CNStageIntLLROutputS6xD(31)(5);
  VNStageIntLLRInputS6xD(22)(0) <= CNStageIntLLROutputS6xD(32)(0);
  VNStageIntLLRInputS6xD(86)(0) <= CNStageIntLLROutputS6xD(32)(1);
  VNStageIntLLRInputS6xD(150)(0) <= CNStageIntLLROutputS6xD(32)(2);
  VNStageIntLLRInputS6xD(214)(0) <= CNStageIntLLROutputS6xD(32)(3);
  VNStageIntLLRInputS6xD(278)(0) <= CNStageIntLLROutputS6xD(32)(4);
  VNStageIntLLRInputS6xD(342)(0) <= CNStageIntLLROutputS6xD(32)(5);
  VNStageIntLLRInputS6xD(21)(0) <= CNStageIntLLROutputS6xD(33)(0);
  VNStageIntLLRInputS6xD(85)(0) <= CNStageIntLLROutputS6xD(33)(1);
  VNStageIntLLRInputS6xD(149)(0) <= CNStageIntLLROutputS6xD(33)(2);
  VNStageIntLLRInputS6xD(213)(0) <= CNStageIntLLROutputS6xD(33)(3);
  VNStageIntLLRInputS6xD(277)(0) <= CNStageIntLLROutputS6xD(33)(4);
  VNStageIntLLRInputS6xD(341)(0) <= CNStageIntLLROutputS6xD(33)(5);
  VNStageIntLLRInputS6xD(20)(0) <= CNStageIntLLROutputS6xD(34)(0);
  VNStageIntLLRInputS6xD(84)(0) <= CNStageIntLLROutputS6xD(34)(1);
  VNStageIntLLRInputS6xD(148)(0) <= CNStageIntLLROutputS6xD(34)(2);
  VNStageIntLLRInputS6xD(212)(0) <= CNStageIntLLROutputS6xD(34)(3);
  VNStageIntLLRInputS6xD(276)(0) <= CNStageIntLLROutputS6xD(34)(4);
  VNStageIntLLRInputS6xD(340)(0) <= CNStageIntLLROutputS6xD(34)(5);
  VNStageIntLLRInputS6xD(19)(0) <= CNStageIntLLROutputS6xD(35)(0);
  VNStageIntLLRInputS6xD(83)(0) <= CNStageIntLLROutputS6xD(35)(1);
  VNStageIntLLRInputS6xD(147)(0) <= CNStageIntLLROutputS6xD(35)(2);
  VNStageIntLLRInputS6xD(211)(0) <= CNStageIntLLROutputS6xD(35)(3);
  VNStageIntLLRInputS6xD(275)(0) <= CNStageIntLLROutputS6xD(35)(4);
  VNStageIntLLRInputS6xD(339)(0) <= CNStageIntLLROutputS6xD(35)(5);
  VNStageIntLLRInputS6xD(18)(0) <= CNStageIntLLROutputS6xD(36)(0);
  VNStageIntLLRInputS6xD(82)(0) <= CNStageIntLLROutputS6xD(36)(1);
  VNStageIntLLRInputS6xD(146)(0) <= CNStageIntLLROutputS6xD(36)(2);
  VNStageIntLLRInputS6xD(210)(0) <= CNStageIntLLROutputS6xD(36)(3);
  VNStageIntLLRInputS6xD(274)(0) <= CNStageIntLLROutputS6xD(36)(4);
  VNStageIntLLRInputS6xD(338)(0) <= CNStageIntLLROutputS6xD(36)(5);
  VNStageIntLLRInputS6xD(17)(0) <= CNStageIntLLROutputS6xD(37)(0);
  VNStageIntLLRInputS6xD(81)(0) <= CNStageIntLLROutputS6xD(37)(1);
  VNStageIntLLRInputS6xD(145)(0) <= CNStageIntLLROutputS6xD(37)(2);
  VNStageIntLLRInputS6xD(209)(0) <= CNStageIntLLROutputS6xD(37)(3);
  VNStageIntLLRInputS6xD(273)(0) <= CNStageIntLLROutputS6xD(37)(4);
  VNStageIntLLRInputS6xD(337)(0) <= CNStageIntLLROutputS6xD(37)(5);
  VNStageIntLLRInputS6xD(16)(0) <= CNStageIntLLROutputS6xD(38)(0);
  VNStageIntLLRInputS6xD(80)(0) <= CNStageIntLLROutputS6xD(38)(1);
  VNStageIntLLRInputS6xD(144)(0) <= CNStageIntLLROutputS6xD(38)(2);
  VNStageIntLLRInputS6xD(208)(0) <= CNStageIntLLROutputS6xD(38)(3);
  VNStageIntLLRInputS6xD(272)(0) <= CNStageIntLLROutputS6xD(38)(4);
  VNStageIntLLRInputS6xD(336)(0) <= CNStageIntLLROutputS6xD(38)(5);
  VNStageIntLLRInputS6xD(15)(0) <= CNStageIntLLROutputS6xD(39)(0);
  VNStageIntLLRInputS6xD(79)(0) <= CNStageIntLLROutputS6xD(39)(1);
  VNStageIntLLRInputS6xD(143)(0) <= CNStageIntLLROutputS6xD(39)(2);
  VNStageIntLLRInputS6xD(207)(0) <= CNStageIntLLROutputS6xD(39)(3);
  VNStageIntLLRInputS6xD(271)(0) <= CNStageIntLLROutputS6xD(39)(4);
  VNStageIntLLRInputS6xD(335)(0) <= CNStageIntLLROutputS6xD(39)(5);
  VNStageIntLLRInputS6xD(14)(0) <= CNStageIntLLROutputS6xD(40)(0);
  VNStageIntLLRInputS6xD(78)(0) <= CNStageIntLLROutputS6xD(40)(1);
  VNStageIntLLRInputS6xD(142)(0) <= CNStageIntLLROutputS6xD(40)(2);
  VNStageIntLLRInputS6xD(206)(0) <= CNStageIntLLROutputS6xD(40)(3);
  VNStageIntLLRInputS6xD(270)(0) <= CNStageIntLLROutputS6xD(40)(4);
  VNStageIntLLRInputS6xD(334)(0) <= CNStageIntLLROutputS6xD(40)(5);
  VNStageIntLLRInputS6xD(12)(0) <= CNStageIntLLROutputS6xD(41)(0);
  VNStageIntLLRInputS6xD(76)(0) <= CNStageIntLLROutputS6xD(41)(1);
  VNStageIntLLRInputS6xD(140)(0) <= CNStageIntLLROutputS6xD(41)(2);
  VNStageIntLLRInputS6xD(204)(0) <= CNStageIntLLROutputS6xD(41)(3);
  VNStageIntLLRInputS6xD(268)(0) <= CNStageIntLLROutputS6xD(41)(4);
  VNStageIntLLRInputS6xD(332)(0) <= CNStageIntLLROutputS6xD(41)(5);
  VNStageIntLLRInputS6xD(11)(0) <= CNStageIntLLROutputS6xD(42)(0);
  VNStageIntLLRInputS6xD(75)(0) <= CNStageIntLLROutputS6xD(42)(1);
  VNStageIntLLRInputS6xD(139)(0) <= CNStageIntLLROutputS6xD(42)(2);
  VNStageIntLLRInputS6xD(203)(0) <= CNStageIntLLROutputS6xD(42)(3);
  VNStageIntLLRInputS6xD(267)(0) <= CNStageIntLLROutputS6xD(42)(4);
  VNStageIntLLRInputS6xD(331)(0) <= CNStageIntLLROutputS6xD(42)(5);
  VNStageIntLLRInputS6xD(10)(0) <= CNStageIntLLROutputS6xD(43)(0);
  VNStageIntLLRInputS6xD(74)(0) <= CNStageIntLLROutputS6xD(43)(1);
  VNStageIntLLRInputS6xD(138)(0) <= CNStageIntLLROutputS6xD(43)(2);
  VNStageIntLLRInputS6xD(202)(0) <= CNStageIntLLROutputS6xD(43)(3);
  VNStageIntLLRInputS6xD(266)(0) <= CNStageIntLLROutputS6xD(43)(4);
  VNStageIntLLRInputS6xD(330)(0) <= CNStageIntLLROutputS6xD(43)(5);
  VNStageIntLLRInputS6xD(9)(0) <= CNStageIntLLROutputS6xD(44)(0);
  VNStageIntLLRInputS6xD(73)(0) <= CNStageIntLLROutputS6xD(44)(1);
  VNStageIntLLRInputS6xD(137)(0) <= CNStageIntLLROutputS6xD(44)(2);
  VNStageIntLLRInputS6xD(201)(0) <= CNStageIntLLROutputS6xD(44)(3);
  VNStageIntLLRInputS6xD(265)(0) <= CNStageIntLLROutputS6xD(44)(4);
  VNStageIntLLRInputS6xD(329)(0) <= CNStageIntLLROutputS6xD(44)(5);
  VNStageIntLLRInputS6xD(8)(0) <= CNStageIntLLROutputS6xD(45)(0);
  VNStageIntLLRInputS6xD(72)(0) <= CNStageIntLLROutputS6xD(45)(1);
  VNStageIntLLRInputS6xD(136)(0) <= CNStageIntLLROutputS6xD(45)(2);
  VNStageIntLLRInputS6xD(200)(0) <= CNStageIntLLROutputS6xD(45)(3);
  VNStageIntLLRInputS6xD(264)(0) <= CNStageIntLLROutputS6xD(45)(4);
  VNStageIntLLRInputS6xD(328)(0) <= CNStageIntLLROutputS6xD(45)(5);
  VNStageIntLLRInputS6xD(7)(0) <= CNStageIntLLROutputS6xD(46)(0);
  VNStageIntLLRInputS6xD(71)(0) <= CNStageIntLLROutputS6xD(46)(1);
  VNStageIntLLRInputS6xD(135)(0) <= CNStageIntLLROutputS6xD(46)(2);
  VNStageIntLLRInputS6xD(199)(0) <= CNStageIntLLROutputS6xD(46)(3);
  VNStageIntLLRInputS6xD(263)(0) <= CNStageIntLLROutputS6xD(46)(4);
  VNStageIntLLRInputS6xD(327)(0) <= CNStageIntLLROutputS6xD(46)(5);
  VNStageIntLLRInputS6xD(6)(0) <= CNStageIntLLROutputS6xD(47)(0);
  VNStageIntLLRInputS6xD(70)(0) <= CNStageIntLLROutputS6xD(47)(1);
  VNStageIntLLRInputS6xD(134)(0) <= CNStageIntLLROutputS6xD(47)(2);
  VNStageIntLLRInputS6xD(198)(0) <= CNStageIntLLROutputS6xD(47)(3);
  VNStageIntLLRInputS6xD(262)(0) <= CNStageIntLLROutputS6xD(47)(4);
  VNStageIntLLRInputS6xD(326)(0) <= CNStageIntLLROutputS6xD(47)(5);
  VNStageIntLLRInputS6xD(5)(0) <= CNStageIntLLROutputS6xD(48)(0);
  VNStageIntLLRInputS6xD(69)(0) <= CNStageIntLLROutputS6xD(48)(1);
  VNStageIntLLRInputS6xD(133)(0) <= CNStageIntLLROutputS6xD(48)(2);
  VNStageIntLLRInputS6xD(197)(0) <= CNStageIntLLROutputS6xD(48)(3);
  VNStageIntLLRInputS6xD(261)(0) <= CNStageIntLLROutputS6xD(48)(4);
  VNStageIntLLRInputS6xD(325)(0) <= CNStageIntLLROutputS6xD(48)(5);
  VNStageIntLLRInputS6xD(4)(0) <= CNStageIntLLROutputS6xD(49)(0);
  VNStageIntLLRInputS6xD(68)(0) <= CNStageIntLLROutputS6xD(49)(1);
  VNStageIntLLRInputS6xD(132)(0) <= CNStageIntLLROutputS6xD(49)(2);
  VNStageIntLLRInputS6xD(196)(0) <= CNStageIntLLROutputS6xD(49)(3);
  VNStageIntLLRInputS6xD(260)(0) <= CNStageIntLLROutputS6xD(49)(4);
  VNStageIntLLRInputS6xD(324)(0) <= CNStageIntLLROutputS6xD(49)(5);
  VNStageIntLLRInputS6xD(2)(0) <= CNStageIntLLROutputS6xD(50)(0);
  VNStageIntLLRInputS6xD(66)(0) <= CNStageIntLLROutputS6xD(50)(1);
  VNStageIntLLRInputS6xD(130)(0) <= CNStageIntLLROutputS6xD(50)(2);
  VNStageIntLLRInputS6xD(194)(0) <= CNStageIntLLROutputS6xD(50)(3);
  VNStageIntLLRInputS6xD(258)(0) <= CNStageIntLLROutputS6xD(50)(4);
  VNStageIntLLRInputS6xD(322)(0) <= CNStageIntLLROutputS6xD(50)(5);
  VNStageIntLLRInputS6xD(1)(0) <= CNStageIntLLROutputS6xD(51)(0);
  VNStageIntLLRInputS6xD(65)(0) <= CNStageIntLLROutputS6xD(51)(1);
  VNStageIntLLRInputS6xD(129)(0) <= CNStageIntLLROutputS6xD(51)(2);
  VNStageIntLLRInputS6xD(193)(0) <= CNStageIntLLROutputS6xD(51)(3);
  VNStageIntLLRInputS6xD(257)(0) <= CNStageIntLLROutputS6xD(51)(4);
  VNStageIntLLRInputS6xD(321)(0) <= CNStageIntLLROutputS6xD(51)(5);
  VNStageIntLLRInputS6xD(63)(0) <= CNStageIntLLROutputS6xD(52)(0);
  VNStageIntLLRInputS6xD(127)(0) <= CNStageIntLLROutputS6xD(52)(1);
  VNStageIntLLRInputS6xD(191)(0) <= CNStageIntLLROutputS6xD(52)(2);
  VNStageIntLLRInputS6xD(255)(0) <= CNStageIntLLROutputS6xD(52)(3);
  VNStageIntLLRInputS6xD(319)(0) <= CNStageIntLLROutputS6xD(52)(4);
  VNStageIntLLRInputS6xD(383)(0) <= CNStageIntLLROutputS6xD(52)(5);
  VNStageIntLLRInputS6xD(0)(0) <= CNStageIntLLROutputS6xD(53)(0);
  VNStageIntLLRInputS6xD(64)(0) <= CNStageIntLLROutputS6xD(53)(1);
  VNStageIntLLRInputS6xD(128)(0) <= CNStageIntLLROutputS6xD(53)(2);
  VNStageIntLLRInputS6xD(192)(0) <= CNStageIntLLROutputS6xD(53)(3);
  VNStageIntLLRInputS6xD(256)(0) <= CNStageIntLLROutputS6xD(53)(4);
  VNStageIntLLRInputS6xD(320)(0) <= CNStageIntLLROutputS6xD(53)(5);
  VNStageIntLLRInputS6xD(42)(1) <= CNStageIntLLROutputS6xD(54)(0);
  VNStageIntLLRInputS6xD(112)(1) <= CNStageIntLLROutputS6xD(54)(1);
  VNStageIntLLRInputS6xD(182)(1) <= CNStageIntLLROutputS6xD(54)(2);
  VNStageIntLLRInputS6xD(203)(1) <= CNStageIntLLROutputS6xD(54)(3);
  VNStageIntLLRInputS6xD(259)(0) <= CNStageIntLLROutputS6xD(54)(4);
  VNStageIntLLRInputS6xD(361)(1) <= CNStageIntLLROutputS6xD(54)(5);
  VNStageIntLLRInputS6xD(41)(1) <= CNStageIntLLROutputS6xD(55)(0);
  VNStageIntLLRInputS6xD(117)(1) <= CNStageIntLLROutputS6xD(55)(1);
  VNStageIntLLRInputS6xD(138)(1) <= CNStageIntLLROutputS6xD(55)(2);
  VNStageIntLLRInputS6xD(194)(1) <= CNStageIntLLROutputS6xD(55)(3);
  VNStageIntLLRInputS6xD(296)(1) <= CNStageIntLLROutputS6xD(55)(4);
  VNStageIntLLRInputS6xD(362)(1) <= CNStageIntLLROutputS6xD(55)(5);
  VNStageIntLLRInputS6xD(40)(1) <= CNStageIntLLROutputS6xD(56)(0);
  VNStageIntLLRInputS6xD(73)(1) <= CNStageIntLLROutputS6xD(56)(1);
  VNStageIntLLRInputS6xD(129)(1) <= CNStageIntLLROutputS6xD(56)(2);
  VNStageIntLLRInputS6xD(231)(1) <= CNStageIntLLROutputS6xD(56)(3);
  VNStageIntLLRInputS6xD(297)(1) <= CNStageIntLLROutputS6xD(56)(4);
  VNStageIntLLRInputS6xD(323)(0) <= CNStageIntLLROutputS6xD(56)(5);
  VNStageIntLLRInputS6xD(39)(1) <= CNStageIntLLROutputS6xD(57)(0);
  VNStageIntLLRInputS6xD(127)(1) <= CNStageIntLLROutputS6xD(57)(1);
  VNStageIntLLRInputS6xD(166)(1) <= CNStageIntLLROutputS6xD(57)(2);
  VNStageIntLLRInputS6xD(232)(1) <= CNStageIntLLROutputS6xD(57)(3);
  VNStageIntLLRInputS6xD(258)(1) <= CNStageIntLLROutputS6xD(57)(4);
  VNStageIntLLRInputS6xD(344)(1) <= CNStageIntLLROutputS6xD(57)(5);
  VNStageIntLLRInputS6xD(38)(1) <= CNStageIntLLROutputS6xD(58)(0);
  VNStageIntLLRInputS6xD(101)(1) <= CNStageIntLLROutputS6xD(58)(1);
  VNStageIntLLRInputS6xD(167)(1) <= CNStageIntLLROutputS6xD(58)(2);
  VNStageIntLLRInputS6xD(193)(1) <= CNStageIntLLROutputS6xD(58)(3);
  VNStageIntLLRInputS6xD(279)(1) <= CNStageIntLLROutputS6xD(58)(4);
  VNStageIntLLRInputS6xD(340)(1) <= CNStageIntLLROutputS6xD(58)(5);
  VNStageIntLLRInputS6xD(37)(1) <= CNStageIntLLROutputS6xD(59)(0);
  VNStageIntLLRInputS6xD(102)(1) <= CNStageIntLLROutputS6xD(59)(1);
  VNStageIntLLRInputS6xD(191)(1) <= CNStageIntLLROutputS6xD(59)(2);
  VNStageIntLLRInputS6xD(214)(1) <= CNStageIntLLROutputS6xD(59)(3);
  VNStageIntLLRInputS6xD(275)(1) <= CNStageIntLLROutputS6xD(59)(4);
  VNStageIntLLRInputS6xD(355)(1) <= CNStageIntLLROutputS6xD(59)(5);
  VNStageIntLLRInputS6xD(36)(1) <= CNStageIntLLROutputS6xD(60)(0);
  VNStageIntLLRInputS6xD(126)(0) <= CNStageIntLLROutputS6xD(60)(1);
  VNStageIntLLRInputS6xD(149)(1) <= CNStageIntLLROutputS6xD(60)(2);
  VNStageIntLLRInputS6xD(210)(1) <= CNStageIntLLROutputS6xD(60)(3);
  VNStageIntLLRInputS6xD(290)(1) <= CNStageIntLLROutputS6xD(60)(4);
  VNStageIntLLRInputS6xD(381)(0) <= CNStageIntLLROutputS6xD(60)(5);
  VNStageIntLLRInputS6xD(35)(1) <= CNStageIntLLROutputS6xD(61)(0);
  VNStageIntLLRInputS6xD(84)(1) <= CNStageIntLLROutputS6xD(61)(1);
  VNStageIntLLRInputS6xD(145)(1) <= CNStageIntLLROutputS6xD(61)(2);
  VNStageIntLLRInputS6xD(225)(1) <= CNStageIntLLROutputS6xD(61)(3);
  VNStageIntLLRInputS6xD(316)(0) <= CNStageIntLLROutputS6xD(61)(4);
  VNStageIntLLRInputS6xD(357)(1) <= CNStageIntLLROutputS6xD(61)(5);
  VNStageIntLLRInputS6xD(34)(1) <= CNStageIntLLROutputS6xD(62)(0);
  VNStageIntLLRInputS6xD(80)(1) <= CNStageIntLLROutputS6xD(62)(1);
  VNStageIntLLRInputS6xD(160)(1) <= CNStageIntLLROutputS6xD(62)(2);
  VNStageIntLLRInputS6xD(251)(0) <= CNStageIntLLROutputS6xD(62)(3);
  VNStageIntLLRInputS6xD(292)(1) <= CNStageIntLLROutputS6xD(62)(4);
  VNStageIntLLRInputS6xD(326)(1) <= CNStageIntLLROutputS6xD(62)(5);
  VNStageIntLLRInputS6xD(33)(1) <= CNStageIntLLROutputS6xD(63)(0);
  VNStageIntLLRInputS6xD(95)(1) <= CNStageIntLLROutputS6xD(63)(1);
  VNStageIntLLRInputS6xD(186)(0) <= CNStageIntLLROutputS6xD(63)(2);
  VNStageIntLLRInputS6xD(227)(1) <= CNStageIntLLROutputS6xD(63)(3);
  VNStageIntLLRInputS6xD(261)(1) <= CNStageIntLLROutputS6xD(63)(4);
  VNStageIntLLRInputS6xD(342)(1) <= CNStageIntLLROutputS6xD(63)(5);
  VNStageIntLLRInputS6xD(32)(1) <= CNStageIntLLROutputS6xD(64)(0);
  VNStageIntLLRInputS6xD(121)(0) <= CNStageIntLLROutputS6xD(64)(1);
  VNStageIntLLRInputS6xD(162)(1) <= CNStageIntLLROutputS6xD(64)(2);
  VNStageIntLLRInputS6xD(196)(1) <= CNStageIntLLROutputS6xD(64)(3);
  VNStageIntLLRInputS6xD(277)(1) <= CNStageIntLLROutputS6xD(64)(4);
  VNStageIntLLRInputS6xD(375)(1) <= CNStageIntLLROutputS6xD(64)(5);
  VNStageIntLLRInputS6xD(31)(1) <= CNStageIntLLROutputS6xD(65)(0);
  VNStageIntLLRInputS6xD(97)(1) <= CNStageIntLLROutputS6xD(65)(1);
  VNStageIntLLRInputS6xD(131)(0) <= CNStageIntLLROutputS6xD(65)(2);
  VNStageIntLLRInputS6xD(212)(1) <= CNStageIntLLROutputS6xD(65)(3);
  VNStageIntLLRInputS6xD(310)(1) <= CNStageIntLLROutputS6xD(65)(4);
  VNStageIntLLRInputS6xD(321)(1) <= CNStageIntLLROutputS6xD(65)(5);
  VNStageIntLLRInputS6xD(30)(1) <= CNStageIntLLROutputS6xD(66)(0);
  VNStageIntLLRInputS6xD(66)(1) <= CNStageIntLLROutputS6xD(66)(1);
  VNStageIntLLRInputS6xD(147)(1) <= CNStageIntLLROutputS6xD(66)(2);
  VNStageIntLLRInputS6xD(245)(1) <= CNStageIntLLROutputS6xD(66)(3);
  VNStageIntLLRInputS6xD(319)(1) <= CNStageIntLLROutputS6xD(66)(4);
  VNStageIntLLRInputS6xD(334)(1) <= CNStageIntLLROutputS6xD(66)(5);
  VNStageIntLLRInputS6xD(29)(1) <= CNStageIntLLROutputS6xD(67)(0);
  VNStageIntLLRInputS6xD(82)(1) <= CNStageIntLLROutputS6xD(67)(1);
  VNStageIntLLRInputS6xD(180)(0) <= CNStageIntLLROutputS6xD(67)(2);
  VNStageIntLLRInputS6xD(254)(0) <= CNStageIntLLROutputS6xD(67)(3);
  VNStageIntLLRInputS6xD(269)(0) <= CNStageIntLLROutputS6xD(67)(4);
  VNStageIntLLRInputS6xD(376)(1) <= CNStageIntLLROutputS6xD(67)(5);
  VNStageIntLLRInputS6xD(28)(1) <= CNStageIntLLROutputS6xD(68)(0);
  VNStageIntLLRInputS6xD(115)(1) <= CNStageIntLLROutputS6xD(68)(1);
  VNStageIntLLRInputS6xD(189)(0) <= CNStageIntLLROutputS6xD(68)(2);
  VNStageIntLLRInputS6xD(204)(1) <= CNStageIntLLROutputS6xD(68)(3);
  VNStageIntLLRInputS6xD(311)(1) <= CNStageIntLLROutputS6xD(68)(4);
  VNStageIntLLRInputS6xD(341)(1) <= CNStageIntLLROutputS6xD(68)(5);
  VNStageIntLLRInputS6xD(27)(1) <= CNStageIntLLROutputS6xD(69)(0);
  VNStageIntLLRInputS6xD(124)(0) <= CNStageIntLLROutputS6xD(69)(1);
  VNStageIntLLRInputS6xD(139)(1) <= CNStageIntLLROutputS6xD(69)(2);
  VNStageIntLLRInputS6xD(246)(1) <= CNStageIntLLROutputS6xD(69)(3);
  VNStageIntLLRInputS6xD(276)(1) <= CNStageIntLLROutputS6xD(69)(4);
  VNStageIntLLRInputS6xD(343)(1) <= CNStageIntLLROutputS6xD(69)(5);
  VNStageIntLLRInputS6xD(26)(1) <= CNStageIntLLROutputS6xD(70)(0);
  VNStageIntLLRInputS6xD(74)(1) <= CNStageIntLLROutputS6xD(70)(1);
  VNStageIntLLRInputS6xD(181)(1) <= CNStageIntLLROutputS6xD(70)(2);
  VNStageIntLLRInputS6xD(211)(1) <= CNStageIntLLROutputS6xD(70)(3);
  VNStageIntLLRInputS6xD(278)(1) <= CNStageIntLLROutputS6xD(70)(4);
  VNStageIntLLRInputS6xD(325)(1) <= CNStageIntLLROutputS6xD(70)(5);
  VNStageIntLLRInputS6xD(25)(1) <= CNStageIntLLROutputS6xD(71)(0);
  VNStageIntLLRInputS6xD(116)(0) <= CNStageIntLLROutputS6xD(71)(1);
  VNStageIntLLRInputS6xD(146)(1) <= CNStageIntLLROutputS6xD(71)(2);
  VNStageIntLLRInputS6xD(213)(1) <= CNStageIntLLROutputS6xD(71)(3);
  VNStageIntLLRInputS6xD(260)(1) <= CNStageIntLLROutputS6xD(71)(4);
  VNStageIntLLRInputS6xD(332)(1) <= CNStageIntLLROutputS6xD(71)(5);
  VNStageIntLLRInputS6xD(24)(1) <= CNStageIntLLROutputS6xD(72)(0);
  VNStageIntLLRInputS6xD(81)(1) <= CNStageIntLLROutputS6xD(72)(1);
  VNStageIntLLRInputS6xD(148)(1) <= CNStageIntLLROutputS6xD(72)(2);
  VNStageIntLLRInputS6xD(195)(0) <= CNStageIntLLROutputS6xD(72)(3);
  VNStageIntLLRInputS6xD(267)(1) <= CNStageIntLLROutputS6xD(72)(4);
  VNStageIntLLRInputS6xD(359)(1) <= CNStageIntLLROutputS6xD(72)(5);
  VNStageIntLLRInputS6xD(23)(1) <= CNStageIntLLROutputS6xD(73)(0);
  VNStageIntLLRInputS6xD(83)(1) <= CNStageIntLLROutputS6xD(73)(1);
  VNStageIntLLRInputS6xD(130)(1) <= CNStageIntLLROutputS6xD(73)(2);
  VNStageIntLLRInputS6xD(202)(1) <= CNStageIntLLROutputS6xD(73)(3);
  VNStageIntLLRInputS6xD(294)(1) <= CNStageIntLLROutputS6xD(73)(4);
  VNStageIntLLRInputS6xD(347)(1) <= CNStageIntLLROutputS6xD(73)(5);
  VNStageIntLLRInputS6xD(22)(1) <= CNStageIntLLROutputS6xD(74)(0);
  VNStageIntLLRInputS6xD(65)(1) <= CNStageIntLLROutputS6xD(74)(1);
  VNStageIntLLRInputS6xD(137)(1) <= CNStageIntLLROutputS6xD(74)(2);
  VNStageIntLLRInputS6xD(229)(1) <= CNStageIntLLROutputS6xD(74)(3);
  VNStageIntLLRInputS6xD(282)(1) <= CNStageIntLLROutputS6xD(74)(4);
  VNStageIntLLRInputS6xD(353)(1) <= CNStageIntLLROutputS6xD(74)(5);
  VNStageIntLLRInputS6xD(21)(1) <= CNStageIntLLROutputS6xD(75)(0);
  VNStageIntLLRInputS6xD(72)(1) <= CNStageIntLLROutputS6xD(75)(1);
  VNStageIntLLRInputS6xD(164)(1) <= CNStageIntLLROutputS6xD(75)(2);
  VNStageIntLLRInputS6xD(217)(1) <= CNStageIntLLROutputS6xD(75)(3);
  VNStageIntLLRInputS6xD(288)(1) <= CNStageIntLLROutputS6xD(75)(4);
  VNStageIntLLRInputS6xD(348)(1) <= CNStageIntLLROutputS6xD(75)(5);
  VNStageIntLLRInputS6xD(20)(1) <= CNStageIntLLROutputS6xD(76)(0);
  VNStageIntLLRInputS6xD(99)(1) <= CNStageIntLLROutputS6xD(76)(1);
  VNStageIntLLRInputS6xD(152)(1) <= CNStageIntLLROutputS6xD(76)(2);
  VNStageIntLLRInputS6xD(223)(1) <= CNStageIntLLROutputS6xD(76)(3);
  VNStageIntLLRInputS6xD(283)(1) <= CNStageIntLLROutputS6xD(76)(4);
  VNStageIntLLRInputS6xD(358)(1) <= CNStageIntLLROutputS6xD(76)(5);
  VNStageIntLLRInputS6xD(19)(1) <= CNStageIntLLROutputS6xD(77)(0);
  VNStageIntLLRInputS6xD(87)(1) <= CNStageIntLLROutputS6xD(77)(1);
  VNStageIntLLRInputS6xD(158)(1) <= CNStageIntLLROutputS6xD(77)(2);
  VNStageIntLLRInputS6xD(218)(1) <= CNStageIntLLROutputS6xD(77)(3);
  VNStageIntLLRInputS6xD(293)(1) <= CNStageIntLLROutputS6xD(77)(4);
  VNStageIntLLRInputS6xD(380)(0) <= CNStageIntLLROutputS6xD(77)(5);
  VNStageIntLLRInputS6xD(18)(1) <= CNStageIntLLROutputS6xD(78)(0);
  VNStageIntLLRInputS6xD(93)(1) <= CNStageIntLLROutputS6xD(78)(1);
  VNStageIntLLRInputS6xD(153)(1) <= CNStageIntLLROutputS6xD(78)(2);
  VNStageIntLLRInputS6xD(228)(1) <= CNStageIntLLROutputS6xD(78)(3);
  VNStageIntLLRInputS6xD(315)(0) <= CNStageIntLLROutputS6xD(78)(4);
  VNStageIntLLRInputS6xD(335)(1) <= CNStageIntLLROutputS6xD(78)(5);
  VNStageIntLLRInputS6xD(17)(1) <= CNStageIntLLROutputS6xD(79)(0);
  VNStageIntLLRInputS6xD(88)(1) <= CNStageIntLLROutputS6xD(79)(1);
  VNStageIntLLRInputS6xD(163)(1) <= CNStageIntLLROutputS6xD(79)(2);
  VNStageIntLLRInputS6xD(250)(0) <= CNStageIntLLROutputS6xD(79)(3);
  VNStageIntLLRInputS6xD(270)(1) <= CNStageIntLLROutputS6xD(79)(4);
  VNStageIntLLRInputS6xD(383)(1) <= CNStageIntLLROutputS6xD(79)(5);
  VNStageIntLLRInputS6xD(15)(1) <= CNStageIntLLROutputS6xD(80)(0);
  VNStageIntLLRInputS6xD(120)(1) <= CNStageIntLLROutputS6xD(80)(1);
  VNStageIntLLRInputS6xD(140)(1) <= CNStageIntLLROutputS6xD(80)(2);
  VNStageIntLLRInputS6xD(253)(0) <= CNStageIntLLROutputS6xD(80)(3);
  VNStageIntLLRInputS6xD(305)(1) <= CNStageIntLLROutputS6xD(80)(4);
  VNStageIntLLRInputS6xD(338)(1) <= CNStageIntLLROutputS6xD(80)(5);
  VNStageIntLLRInputS6xD(14)(1) <= CNStageIntLLROutputS6xD(81)(0);
  VNStageIntLLRInputS6xD(75)(1) <= CNStageIntLLROutputS6xD(81)(1);
  VNStageIntLLRInputS6xD(188)(0) <= CNStageIntLLROutputS6xD(81)(2);
  VNStageIntLLRInputS6xD(240)(1) <= CNStageIntLLROutputS6xD(81)(3);
  VNStageIntLLRInputS6xD(273)(1) <= CNStageIntLLROutputS6xD(81)(4);
  VNStageIntLLRInputS6xD(350)(1) <= CNStageIntLLROutputS6xD(81)(5);
  VNStageIntLLRInputS6xD(13)(0) <= CNStageIntLLROutputS6xD(82)(0);
  VNStageIntLLRInputS6xD(123)(0) <= CNStageIntLLROutputS6xD(82)(1);
  VNStageIntLLRInputS6xD(175)(1) <= CNStageIntLLROutputS6xD(82)(2);
  VNStageIntLLRInputS6xD(208)(1) <= CNStageIntLLROutputS6xD(82)(3);
  VNStageIntLLRInputS6xD(285)(1) <= CNStageIntLLROutputS6xD(82)(4);
  VNStageIntLLRInputS6xD(364)(1) <= CNStageIntLLROutputS6xD(82)(5);
  VNStageIntLLRInputS6xD(12)(1) <= CNStageIntLLROutputS6xD(83)(0);
  VNStageIntLLRInputS6xD(110)(1) <= CNStageIntLLROutputS6xD(83)(1);
  VNStageIntLLRInputS6xD(143)(1) <= CNStageIntLLROutputS6xD(83)(2);
  VNStageIntLLRInputS6xD(220)(1) <= CNStageIntLLROutputS6xD(83)(3);
  VNStageIntLLRInputS6xD(299)(0) <= CNStageIntLLROutputS6xD(83)(4);
  VNStageIntLLRInputS6xD(345)(1) <= CNStageIntLLROutputS6xD(83)(5);
  VNStageIntLLRInputS6xD(11)(1) <= CNStageIntLLROutputS6xD(84)(0);
  VNStageIntLLRInputS6xD(78)(1) <= CNStageIntLLROutputS6xD(84)(1);
  VNStageIntLLRInputS6xD(155)(1) <= CNStageIntLLROutputS6xD(84)(2);
  VNStageIntLLRInputS6xD(234)(1) <= CNStageIntLLROutputS6xD(84)(3);
  VNStageIntLLRInputS6xD(280)(1) <= CNStageIntLLROutputS6xD(84)(4);
  VNStageIntLLRInputS6xD(322)(1) <= CNStageIntLLROutputS6xD(84)(5);
  VNStageIntLLRInputS6xD(10)(1) <= CNStageIntLLROutputS6xD(85)(0);
  VNStageIntLLRInputS6xD(90)(1) <= CNStageIntLLROutputS6xD(85)(1);
  VNStageIntLLRInputS6xD(169)(1) <= CNStageIntLLROutputS6xD(85)(2);
  VNStageIntLLRInputS6xD(215)(1) <= CNStageIntLLROutputS6xD(85)(3);
  VNStageIntLLRInputS6xD(257)(1) <= CNStageIntLLROutputS6xD(85)(4);
  VNStageIntLLRInputS6xD(374)(1) <= CNStageIntLLROutputS6xD(85)(5);
  VNStageIntLLRInputS6xD(9)(1) <= CNStageIntLLROutputS6xD(86)(0);
  VNStageIntLLRInputS6xD(104)(1) <= CNStageIntLLROutputS6xD(86)(1);
  VNStageIntLLRInputS6xD(150)(1) <= CNStageIntLLROutputS6xD(86)(2);
  VNStageIntLLRInputS6xD(255)(1) <= CNStageIntLLROutputS6xD(86)(3);
  VNStageIntLLRInputS6xD(309)(1) <= CNStageIntLLROutputS6xD(86)(4);
  VNStageIntLLRInputS6xD(378)(0) <= CNStageIntLLROutputS6xD(86)(5);
  VNStageIntLLRInputS6xD(7)(1) <= CNStageIntLLROutputS6xD(87)(0);
  VNStageIntLLRInputS6xD(125)(0) <= CNStageIntLLROutputS6xD(87)(1);
  VNStageIntLLRInputS6xD(179)(1) <= CNStageIntLLROutputS6xD(87)(2);
  VNStageIntLLRInputS6xD(248)(1) <= CNStageIntLLROutputS6xD(87)(3);
  VNStageIntLLRInputS6xD(306)(1) <= CNStageIntLLROutputS6xD(87)(4);
  VNStageIntLLRInputS6xD(382)(0) <= CNStageIntLLROutputS6xD(87)(5);
  VNStageIntLLRInputS6xD(6)(1) <= CNStageIntLLROutputS6xD(88)(0);
  VNStageIntLLRInputS6xD(114)(1) <= CNStageIntLLROutputS6xD(88)(1);
  VNStageIntLLRInputS6xD(183)(1) <= CNStageIntLLROutputS6xD(88)(2);
  VNStageIntLLRInputS6xD(241)(1) <= CNStageIntLLROutputS6xD(88)(3);
  VNStageIntLLRInputS6xD(317)(0) <= CNStageIntLLROutputS6xD(88)(4);
  VNStageIntLLRInputS6xD(354)(1) <= CNStageIntLLROutputS6xD(88)(5);
  VNStageIntLLRInputS6xD(5)(1) <= CNStageIntLLROutputS6xD(89)(0);
  VNStageIntLLRInputS6xD(118)(1) <= CNStageIntLLROutputS6xD(89)(1);
  VNStageIntLLRInputS6xD(176)(1) <= CNStageIntLLROutputS6xD(89)(2);
  VNStageIntLLRInputS6xD(252)(0) <= CNStageIntLLROutputS6xD(89)(3);
  VNStageIntLLRInputS6xD(289)(1) <= CNStageIntLLROutputS6xD(89)(4);
  VNStageIntLLRInputS6xD(346)(1) <= CNStageIntLLROutputS6xD(89)(5);
  VNStageIntLLRInputS6xD(4)(1) <= CNStageIntLLROutputS6xD(90)(0);
  VNStageIntLLRInputS6xD(111)(1) <= CNStageIntLLROutputS6xD(90)(1);
  VNStageIntLLRInputS6xD(187)(0) <= CNStageIntLLROutputS6xD(90)(2);
  VNStageIntLLRInputS6xD(224)(1) <= CNStageIntLLROutputS6xD(90)(3);
  VNStageIntLLRInputS6xD(281)(1) <= CNStageIntLLROutputS6xD(90)(4);
  VNStageIntLLRInputS6xD(363)(0) <= CNStageIntLLROutputS6xD(90)(5);
  VNStageIntLLRInputS6xD(3)(0) <= CNStageIntLLROutputS6xD(91)(0);
  VNStageIntLLRInputS6xD(122)(0) <= CNStageIntLLROutputS6xD(91)(1);
  VNStageIntLLRInputS6xD(159)(1) <= CNStageIntLLROutputS6xD(91)(2);
  VNStageIntLLRInputS6xD(216)(1) <= CNStageIntLLROutputS6xD(91)(3);
  VNStageIntLLRInputS6xD(298)(1) <= CNStageIntLLROutputS6xD(91)(4);
  VNStageIntLLRInputS6xD(360)(1) <= CNStageIntLLROutputS6xD(91)(5);
  VNStageIntLLRInputS6xD(2)(1) <= CNStageIntLLROutputS6xD(92)(0);
  VNStageIntLLRInputS6xD(94)(1) <= CNStageIntLLROutputS6xD(92)(1);
  VNStageIntLLRInputS6xD(151)(1) <= CNStageIntLLROutputS6xD(92)(2);
  VNStageIntLLRInputS6xD(233)(1) <= CNStageIntLLROutputS6xD(92)(3);
  VNStageIntLLRInputS6xD(295)(1) <= CNStageIntLLROutputS6xD(92)(4);
  VNStageIntLLRInputS6xD(331)(1) <= CNStageIntLLROutputS6xD(92)(5);
  VNStageIntLLRInputS6xD(63)(1) <= CNStageIntLLROutputS6xD(93)(0);
  VNStageIntLLRInputS6xD(103)(1) <= CNStageIntLLROutputS6xD(93)(1);
  VNStageIntLLRInputS6xD(165)(1) <= CNStageIntLLROutputS6xD(93)(2);
  VNStageIntLLRInputS6xD(201)(1) <= CNStageIntLLROutputS6xD(93)(3);
  VNStageIntLLRInputS6xD(286)(1) <= CNStageIntLLROutputS6xD(93)(4);
  VNStageIntLLRInputS6xD(337)(1) <= CNStageIntLLROutputS6xD(93)(5);
  VNStageIntLLRInputS6xD(62)(0) <= CNStageIntLLROutputS6xD(94)(0);
  VNStageIntLLRInputS6xD(100)(1) <= CNStageIntLLROutputS6xD(94)(1);
  VNStageIntLLRInputS6xD(136)(1) <= CNStageIntLLROutputS6xD(94)(2);
  VNStageIntLLRInputS6xD(221)(1) <= CNStageIntLLROutputS6xD(94)(3);
  VNStageIntLLRInputS6xD(272)(1) <= CNStageIntLLROutputS6xD(94)(4);
  VNStageIntLLRInputS6xD(327)(1) <= CNStageIntLLROutputS6xD(94)(5);
  VNStageIntLLRInputS6xD(61)(0) <= CNStageIntLLROutputS6xD(95)(0);
  VNStageIntLLRInputS6xD(71)(1) <= CNStageIntLLROutputS6xD(95)(1);
  VNStageIntLLRInputS6xD(156)(1) <= CNStageIntLLROutputS6xD(95)(2);
  VNStageIntLLRInputS6xD(207)(1) <= CNStageIntLLROutputS6xD(95)(3);
  VNStageIntLLRInputS6xD(262)(1) <= CNStageIntLLROutputS6xD(95)(4);
  VNStageIntLLRInputS6xD(356)(1) <= CNStageIntLLROutputS6xD(95)(5);
  VNStageIntLLRInputS6xD(60)(0) <= CNStageIntLLROutputS6xD(96)(0);
  VNStageIntLLRInputS6xD(91)(1) <= CNStageIntLLROutputS6xD(96)(1);
  VNStageIntLLRInputS6xD(142)(1) <= CNStageIntLLROutputS6xD(96)(2);
  VNStageIntLLRInputS6xD(197)(1) <= CNStageIntLLROutputS6xD(96)(3);
  VNStageIntLLRInputS6xD(291)(1) <= CNStageIntLLROutputS6xD(96)(4);
  VNStageIntLLRInputS6xD(339)(1) <= CNStageIntLLROutputS6xD(96)(5);
  VNStageIntLLRInputS6xD(58)(0) <= CNStageIntLLROutputS6xD(97)(0);
  VNStageIntLLRInputS6xD(67)(0) <= CNStageIntLLROutputS6xD(97)(1);
  VNStageIntLLRInputS6xD(161)(1) <= CNStageIntLLROutputS6xD(97)(2);
  VNStageIntLLRInputS6xD(209)(1) <= CNStageIntLLROutputS6xD(97)(3);
  VNStageIntLLRInputS6xD(304)(1) <= CNStageIntLLROutputS6xD(97)(4);
  VNStageIntLLRInputS6xD(329)(1) <= CNStageIntLLROutputS6xD(97)(5);
  VNStageIntLLRInputS6xD(57)(0) <= CNStageIntLLROutputS6xD(98)(0);
  VNStageIntLLRInputS6xD(96)(1) <= CNStageIntLLROutputS6xD(98)(1);
  VNStageIntLLRInputS6xD(144)(1) <= CNStageIntLLROutputS6xD(98)(2);
  VNStageIntLLRInputS6xD(239)(1) <= CNStageIntLLROutputS6xD(98)(3);
  VNStageIntLLRInputS6xD(264)(1) <= CNStageIntLLROutputS6xD(98)(4);
  VNStageIntLLRInputS6xD(365)(1) <= CNStageIntLLROutputS6xD(98)(5);
  VNStageIntLLRInputS6xD(56)(1) <= CNStageIntLLROutputS6xD(99)(0);
  VNStageIntLLRInputS6xD(79)(1) <= CNStageIntLLROutputS6xD(99)(1);
  VNStageIntLLRInputS6xD(174)(1) <= CNStageIntLLROutputS6xD(99)(2);
  VNStageIntLLRInputS6xD(199)(1) <= CNStageIntLLROutputS6xD(99)(3);
  VNStageIntLLRInputS6xD(300)(1) <= CNStageIntLLROutputS6xD(99)(4);
  VNStageIntLLRInputS6xD(349)(1) <= CNStageIntLLROutputS6xD(99)(5);
  VNStageIntLLRInputS6xD(55)(1) <= CNStageIntLLROutputS6xD(100)(0);
  VNStageIntLLRInputS6xD(109)(1) <= CNStageIntLLROutputS6xD(100)(1);
  VNStageIntLLRInputS6xD(134)(1) <= CNStageIntLLROutputS6xD(100)(2);
  VNStageIntLLRInputS6xD(235)(0) <= CNStageIntLLROutputS6xD(100)(3);
  VNStageIntLLRInputS6xD(284)(1) <= CNStageIntLLROutputS6xD(100)(4);
  VNStageIntLLRInputS6xD(352)(1) <= CNStageIntLLROutputS6xD(100)(5);
  VNStageIntLLRInputS6xD(54)(1) <= CNStageIntLLROutputS6xD(101)(0);
  VNStageIntLLRInputS6xD(69)(1) <= CNStageIntLLROutputS6xD(101)(1);
  VNStageIntLLRInputS6xD(170)(1) <= CNStageIntLLROutputS6xD(101)(2);
  VNStageIntLLRInputS6xD(219)(1) <= CNStageIntLLROutputS6xD(101)(3);
  VNStageIntLLRInputS6xD(287)(1) <= CNStageIntLLROutputS6xD(101)(4);
  VNStageIntLLRInputS6xD(330)(1) <= CNStageIntLLROutputS6xD(101)(5);
  VNStageIntLLRInputS6xD(52)(0) <= CNStageIntLLROutputS6xD(102)(0);
  VNStageIntLLRInputS6xD(89)(1) <= CNStageIntLLROutputS6xD(102)(1);
  VNStageIntLLRInputS6xD(157)(1) <= CNStageIntLLROutputS6xD(102)(2);
  VNStageIntLLRInputS6xD(200)(1) <= CNStageIntLLROutputS6xD(102)(3);
  VNStageIntLLRInputS6xD(303)(1) <= CNStageIntLLROutputS6xD(102)(4);
  VNStageIntLLRInputS6xD(366)(1) <= CNStageIntLLROutputS6xD(102)(5);
  VNStageIntLLRInputS6xD(51)(1) <= CNStageIntLLROutputS6xD(103)(0);
  VNStageIntLLRInputS6xD(92)(1) <= CNStageIntLLROutputS6xD(103)(1);
  VNStageIntLLRInputS6xD(135)(1) <= CNStageIntLLROutputS6xD(103)(2);
  VNStageIntLLRInputS6xD(238)(1) <= CNStageIntLLROutputS6xD(103)(3);
  VNStageIntLLRInputS6xD(301)(1) <= CNStageIntLLROutputS6xD(103)(4);
  VNStageIntLLRInputS6xD(328)(1) <= CNStageIntLLROutputS6xD(103)(5);
  VNStageIntLLRInputS6xD(50)(1) <= CNStageIntLLROutputS6xD(104)(0);
  VNStageIntLLRInputS6xD(70)(1) <= CNStageIntLLROutputS6xD(104)(1);
  VNStageIntLLRInputS6xD(173)(1) <= CNStageIntLLROutputS6xD(104)(2);
  VNStageIntLLRInputS6xD(236)(1) <= CNStageIntLLROutputS6xD(104)(3);
  VNStageIntLLRInputS6xD(263)(1) <= CNStageIntLLROutputS6xD(104)(4);
  VNStageIntLLRInputS6xD(336)(1) <= CNStageIntLLROutputS6xD(104)(5);
  VNStageIntLLRInputS6xD(49)(1) <= CNStageIntLLROutputS6xD(105)(0);
  VNStageIntLLRInputS6xD(108)(1) <= CNStageIntLLROutputS6xD(105)(1);
  VNStageIntLLRInputS6xD(171)(0) <= CNStageIntLLROutputS6xD(105)(2);
  VNStageIntLLRInputS6xD(198)(1) <= CNStageIntLLROutputS6xD(105)(3);
  VNStageIntLLRInputS6xD(271)(1) <= CNStageIntLLROutputS6xD(105)(4);
  VNStageIntLLRInputS6xD(379)(0) <= CNStageIntLLROutputS6xD(105)(5);
  VNStageIntLLRInputS6xD(46)(1) <= CNStageIntLLROutputS6xD(106)(0);
  VNStageIntLLRInputS6xD(76)(1) <= CNStageIntLLROutputS6xD(106)(1);
  VNStageIntLLRInputS6xD(184)(1) <= CNStageIntLLROutputS6xD(106)(2);
  VNStageIntLLRInputS6xD(243)(1) <= CNStageIntLLROutputS6xD(106)(3);
  VNStageIntLLRInputS6xD(256)(1) <= CNStageIntLLROutputS6xD(106)(4);
  VNStageIntLLRInputS6xD(372)(0) <= CNStageIntLLROutputS6xD(106)(5);
  VNStageIntLLRInputS6xD(45)(1) <= CNStageIntLLROutputS6xD(107)(0);
  VNStageIntLLRInputS6xD(119)(1) <= CNStageIntLLROutputS6xD(107)(1);
  VNStageIntLLRInputS6xD(178)(1) <= CNStageIntLLROutputS6xD(107)(2);
  VNStageIntLLRInputS6xD(192)(1) <= CNStageIntLLROutputS6xD(107)(3);
  VNStageIntLLRInputS6xD(307)(1) <= CNStageIntLLROutputS6xD(107)(4);
  VNStageIntLLRInputS6xD(377)(0) <= CNStageIntLLROutputS6xD(107)(5);
  VNStageIntLLRInputS6xD(44)(1) <= CNStageIntLLROutputS6xD(108)(0);
  VNStageIntLLRInputS6xD(113)(1) <= CNStageIntLLROutputS6xD(108)(1);
  VNStageIntLLRInputS6xD(128)(1) <= CNStageIntLLROutputS6xD(108)(2);
  VNStageIntLLRInputS6xD(242)(1) <= CNStageIntLLROutputS6xD(108)(3);
  VNStageIntLLRInputS6xD(312)(1) <= CNStageIntLLROutputS6xD(108)(4);
  VNStageIntLLRInputS6xD(333)(0) <= CNStageIntLLROutputS6xD(108)(5);
  VNStageIntLLRInputS6xD(43)(0) <= CNStageIntLLROutputS6xD(109)(0);
  VNStageIntLLRInputS6xD(64)(1) <= CNStageIntLLROutputS6xD(109)(1);
  VNStageIntLLRInputS6xD(177)(1) <= CNStageIntLLROutputS6xD(109)(2);
  VNStageIntLLRInputS6xD(247)(1) <= CNStageIntLLROutputS6xD(109)(3);
  VNStageIntLLRInputS6xD(268)(1) <= CNStageIntLLROutputS6xD(109)(4);
  VNStageIntLLRInputS6xD(324)(1) <= CNStageIntLLROutputS6xD(109)(5);
  VNStageIntLLRInputS6xD(0)(1) <= CNStageIntLLROutputS6xD(110)(0);
  VNStageIntLLRInputS6xD(107)(0) <= CNStageIntLLROutputS6xD(110)(1);
  VNStageIntLLRInputS6xD(172)(1) <= CNStageIntLLROutputS6xD(110)(2);
  VNStageIntLLRInputS6xD(237)(1) <= CNStageIntLLROutputS6xD(110)(3);
  VNStageIntLLRInputS6xD(302)(1) <= CNStageIntLLROutputS6xD(110)(4);
  VNStageIntLLRInputS6xD(367)(1) <= CNStageIntLLROutputS6xD(110)(5);
  VNStageIntLLRInputS6xD(32)(2) <= CNStageIntLLROutputS6xD(111)(0);
  VNStageIntLLRInputS6xD(117)(2) <= CNStageIntLLROutputS6xD(111)(1);
  VNStageIntLLRInputS6xD(136)(2) <= CNStageIntLLROutputS6xD(111)(2);
  VNStageIntLLRInputS6xD(198)(2) <= CNStageIntLLROutputS6xD(111)(3);
  VNStageIntLLRInputS6xD(297)(2) <= CNStageIntLLROutputS6xD(111)(4);
  VNStageIntLLRInputS6xD(382)(1) <= CNStageIntLLROutputS6xD(111)(5);
  VNStageIntLLRInputS6xD(30)(2) <= CNStageIntLLROutputS6xD(112)(0);
  VNStageIntLLRInputS6xD(68)(1) <= CNStageIntLLROutputS6xD(112)(1);
  VNStageIntLLRInputS6xD(167)(2) <= CNStageIntLLROutputS6xD(112)(2);
  VNStageIntLLRInputS6xD(252)(1) <= CNStageIntLLROutputS6xD(112)(3);
  VNStageIntLLRInputS6xD(303)(2) <= CNStageIntLLROutputS6xD(112)(4);
  VNStageIntLLRInputS6xD(358)(2) <= CNStageIntLLROutputS6xD(112)(5);
  VNStageIntLLRInputS6xD(29)(2) <= CNStageIntLLROutputS6xD(113)(0);
  VNStageIntLLRInputS6xD(102)(2) <= CNStageIntLLROutputS6xD(113)(1);
  VNStageIntLLRInputS6xD(187)(1) <= CNStageIntLLROutputS6xD(113)(2);
  VNStageIntLLRInputS6xD(238)(2) <= CNStageIntLLROutputS6xD(113)(3);
  VNStageIntLLRInputS6xD(293)(2) <= CNStageIntLLROutputS6xD(113)(4);
  VNStageIntLLRInputS6xD(324)(2) <= CNStageIntLLROutputS6xD(113)(5);
  VNStageIntLLRInputS6xD(28)(2) <= CNStageIntLLROutputS6xD(114)(0);
  VNStageIntLLRInputS6xD(122)(1) <= CNStageIntLLROutputS6xD(114)(1);
  VNStageIntLLRInputS6xD(173)(2) <= CNStageIntLLROutputS6xD(114)(2);
  VNStageIntLLRInputS6xD(228)(2) <= CNStageIntLLROutputS6xD(114)(3);
  VNStageIntLLRInputS6xD(259)(1) <= CNStageIntLLROutputS6xD(114)(4);
  VNStageIntLLRInputS6xD(370)(1) <= CNStageIntLLROutputS6xD(114)(5);
  VNStageIntLLRInputS6xD(27)(2) <= CNStageIntLLROutputS6xD(115)(0);
  VNStageIntLLRInputS6xD(108)(2) <= CNStageIntLLROutputS6xD(115)(1);
  VNStageIntLLRInputS6xD(163)(2) <= CNStageIntLLROutputS6xD(115)(2);
  VNStageIntLLRInputS6xD(194)(2) <= CNStageIntLLROutputS6xD(115)(3);
  VNStageIntLLRInputS6xD(305)(2) <= CNStageIntLLROutputS6xD(115)(4);
  VNStageIntLLRInputS6xD(337)(2) <= CNStageIntLLROutputS6xD(115)(5);
  VNStageIntLLRInputS6xD(26)(2) <= CNStageIntLLROutputS6xD(116)(0);
  VNStageIntLLRInputS6xD(98)(1) <= CNStageIntLLROutputS6xD(116)(1);
  VNStageIntLLRInputS6xD(129)(2) <= CNStageIntLLROutputS6xD(116)(2);
  VNStageIntLLRInputS6xD(240)(2) <= CNStageIntLLROutputS6xD(116)(3);
  VNStageIntLLRInputS6xD(272)(2) <= CNStageIntLLROutputS6xD(116)(4);
  VNStageIntLLRInputS6xD(360)(2) <= CNStageIntLLROutputS6xD(116)(5);
  VNStageIntLLRInputS6xD(25)(2) <= CNStageIntLLROutputS6xD(117)(0);
  VNStageIntLLRInputS6xD(127)(2) <= CNStageIntLLROutputS6xD(117)(1);
  VNStageIntLLRInputS6xD(175)(2) <= CNStageIntLLROutputS6xD(117)(2);
  VNStageIntLLRInputS6xD(207)(2) <= CNStageIntLLROutputS6xD(117)(3);
  VNStageIntLLRInputS6xD(295)(2) <= CNStageIntLLROutputS6xD(117)(4);
  VNStageIntLLRInputS6xD(333)(1) <= CNStageIntLLROutputS6xD(117)(5);
  VNStageIntLLRInputS6xD(24)(2) <= CNStageIntLLROutputS6xD(118)(0);
  VNStageIntLLRInputS6xD(110)(2) <= CNStageIntLLROutputS6xD(118)(1);
  VNStageIntLLRInputS6xD(142)(2) <= CNStageIntLLROutputS6xD(118)(2);
  VNStageIntLLRInputS6xD(230)(1) <= CNStageIntLLROutputS6xD(118)(3);
  VNStageIntLLRInputS6xD(268)(2) <= CNStageIntLLROutputS6xD(118)(4);
  VNStageIntLLRInputS6xD(380)(1) <= CNStageIntLLROutputS6xD(118)(5);
  VNStageIntLLRInputS6xD(23)(2) <= CNStageIntLLROutputS6xD(119)(0);
  VNStageIntLLRInputS6xD(77)(0) <= CNStageIntLLROutputS6xD(119)(1);
  VNStageIntLLRInputS6xD(165)(2) <= CNStageIntLLROutputS6xD(119)(2);
  VNStageIntLLRInputS6xD(203)(2) <= CNStageIntLLROutputS6xD(119)(3);
  VNStageIntLLRInputS6xD(315)(1) <= CNStageIntLLROutputS6xD(119)(4);
  VNStageIntLLRInputS6xD(383)(2) <= CNStageIntLLROutputS6xD(119)(5);
  VNStageIntLLRInputS6xD(22)(2) <= CNStageIntLLROutputS6xD(120)(0);
  VNStageIntLLRInputS6xD(100)(2) <= CNStageIntLLROutputS6xD(120)(1);
  VNStageIntLLRInputS6xD(138)(2) <= CNStageIntLLROutputS6xD(120)(2);
  VNStageIntLLRInputS6xD(250)(1) <= CNStageIntLLROutputS6xD(120)(3);
  VNStageIntLLRInputS6xD(318)(0) <= CNStageIntLLROutputS6xD(120)(4);
  VNStageIntLLRInputS6xD(361)(2) <= CNStageIntLLROutputS6xD(120)(5);
  VNStageIntLLRInputS6xD(21)(2) <= CNStageIntLLROutputS6xD(121)(0);
  VNStageIntLLRInputS6xD(73)(2) <= CNStageIntLLROutputS6xD(121)(1);
  VNStageIntLLRInputS6xD(185)(0) <= CNStageIntLLROutputS6xD(121)(2);
  VNStageIntLLRInputS6xD(253)(1) <= CNStageIntLLROutputS6xD(121)(3);
  VNStageIntLLRInputS6xD(296)(2) <= CNStageIntLLROutputS6xD(121)(4);
  VNStageIntLLRInputS6xD(336)(2) <= CNStageIntLLROutputS6xD(121)(5);
  VNStageIntLLRInputS6xD(19)(2) <= CNStageIntLLROutputS6xD(122)(0);
  VNStageIntLLRInputS6xD(123)(1) <= CNStageIntLLROutputS6xD(122)(1);
  VNStageIntLLRInputS6xD(166)(2) <= CNStageIntLLROutputS6xD(122)(2);
  VNStageIntLLRInputS6xD(206)(1) <= CNStageIntLLROutputS6xD(122)(3);
  VNStageIntLLRInputS6xD(269)(1) <= CNStageIntLLROutputS6xD(122)(4);
  VNStageIntLLRInputS6xD(359)(2) <= CNStageIntLLROutputS6xD(122)(5);
  VNStageIntLLRInputS6xD(18)(2) <= CNStageIntLLROutputS6xD(123)(0);
  VNStageIntLLRInputS6xD(101)(2) <= CNStageIntLLROutputS6xD(123)(1);
  VNStageIntLLRInputS6xD(141)(0) <= CNStageIntLLROutputS6xD(123)(2);
  VNStageIntLLRInputS6xD(204)(2) <= CNStageIntLLROutputS6xD(123)(3);
  VNStageIntLLRInputS6xD(294)(2) <= CNStageIntLLROutputS6xD(123)(4);
  VNStageIntLLRInputS6xD(367)(2) <= CNStageIntLLROutputS6xD(123)(5);
  VNStageIntLLRInputS6xD(17)(2) <= CNStageIntLLROutputS6xD(124)(0);
  VNStageIntLLRInputS6xD(76)(2) <= CNStageIntLLROutputS6xD(124)(1);
  VNStageIntLLRInputS6xD(139)(2) <= CNStageIntLLROutputS6xD(124)(2);
  VNStageIntLLRInputS6xD(229)(2) <= CNStageIntLLROutputS6xD(124)(3);
  VNStageIntLLRInputS6xD(302)(2) <= CNStageIntLLROutputS6xD(124)(4);
  VNStageIntLLRInputS6xD(347)(2) <= CNStageIntLLROutputS6xD(124)(5);
  VNStageIntLLRInputS6xD(16)(1) <= CNStageIntLLROutputS6xD(125)(0);
  VNStageIntLLRInputS6xD(74)(2) <= CNStageIntLLROutputS6xD(125)(1);
  VNStageIntLLRInputS6xD(164)(2) <= CNStageIntLLROutputS6xD(125)(2);
  VNStageIntLLRInputS6xD(237)(2) <= CNStageIntLLROutputS6xD(125)(3);
  VNStageIntLLRInputS6xD(282)(2) <= CNStageIntLLROutputS6xD(125)(4);
  VNStageIntLLRInputS6xD(341)(2) <= CNStageIntLLROutputS6xD(125)(5);
  VNStageIntLLRInputS6xD(15)(2) <= CNStageIntLLROutputS6xD(126)(0);
  VNStageIntLLRInputS6xD(99)(2) <= CNStageIntLLROutputS6xD(126)(1);
  VNStageIntLLRInputS6xD(172)(2) <= CNStageIntLLROutputS6xD(126)(2);
  VNStageIntLLRInputS6xD(217)(2) <= CNStageIntLLROutputS6xD(126)(3);
  VNStageIntLLRInputS6xD(276)(2) <= CNStageIntLLROutputS6xD(126)(4);
  VNStageIntLLRInputS6xD(320)(1) <= CNStageIntLLROutputS6xD(126)(5);
  VNStageIntLLRInputS6xD(14)(2) <= CNStageIntLLROutputS6xD(127)(0);
  VNStageIntLLRInputS6xD(107)(1) <= CNStageIntLLROutputS6xD(127)(1);
  VNStageIntLLRInputS6xD(152)(2) <= CNStageIntLLROutputS6xD(127)(2);
  VNStageIntLLRInputS6xD(211)(2) <= CNStageIntLLROutputS6xD(127)(3);
  VNStageIntLLRInputS6xD(256)(2) <= CNStageIntLLROutputS6xD(127)(4);
  VNStageIntLLRInputS6xD(340)(2) <= CNStageIntLLROutputS6xD(127)(5);
  VNStageIntLLRInputS6xD(13)(1) <= CNStageIntLLROutputS6xD(128)(0);
  VNStageIntLLRInputS6xD(87)(2) <= CNStageIntLLROutputS6xD(128)(1);
  VNStageIntLLRInputS6xD(146)(2) <= CNStageIntLLROutputS6xD(128)(2);
  VNStageIntLLRInputS6xD(192)(2) <= CNStageIntLLROutputS6xD(128)(3);
  VNStageIntLLRInputS6xD(275)(2) <= CNStageIntLLROutputS6xD(128)(4);
  VNStageIntLLRInputS6xD(345)(2) <= CNStageIntLLROutputS6xD(128)(5);
  VNStageIntLLRInputS6xD(12)(2) <= CNStageIntLLROutputS6xD(129)(0);
  VNStageIntLLRInputS6xD(81)(2) <= CNStageIntLLROutputS6xD(129)(1);
  VNStageIntLLRInputS6xD(128)(2) <= CNStageIntLLROutputS6xD(129)(2);
  VNStageIntLLRInputS6xD(210)(2) <= CNStageIntLLROutputS6xD(129)(3);
  VNStageIntLLRInputS6xD(280)(2) <= CNStageIntLLROutputS6xD(129)(4);
  VNStageIntLLRInputS6xD(364)(2) <= CNStageIntLLROutputS6xD(129)(5);
  VNStageIntLLRInputS6xD(11)(2) <= CNStageIntLLROutputS6xD(130)(0);
  VNStageIntLLRInputS6xD(64)(2) <= CNStageIntLLROutputS6xD(130)(1);
  VNStageIntLLRInputS6xD(145)(2) <= CNStageIntLLROutputS6xD(130)(2);
  VNStageIntLLRInputS6xD(215)(2) <= CNStageIntLLROutputS6xD(130)(3);
  VNStageIntLLRInputS6xD(299)(1) <= CNStageIntLLROutputS6xD(130)(4);
  VNStageIntLLRInputS6xD(355)(2) <= CNStageIntLLROutputS6xD(130)(5);
  VNStageIntLLRInputS6xD(10)(2) <= CNStageIntLLROutputS6xD(131)(0);
  VNStageIntLLRInputS6xD(80)(2) <= CNStageIntLLROutputS6xD(131)(1);
  VNStageIntLLRInputS6xD(150)(2) <= CNStageIntLLROutputS6xD(131)(2);
  VNStageIntLLRInputS6xD(234)(2) <= CNStageIntLLROutputS6xD(131)(3);
  VNStageIntLLRInputS6xD(290)(2) <= CNStageIntLLROutputS6xD(131)(4);
  VNStageIntLLRInputS6xD(329)(2) <= CNStageIntLLROutputS6xD(131)(5);
  VNStageIntLLRInputS6xD(9)(2) <= CNStageIntLLROutputS6xD(132)(0);
  VNStageIntLLRInputS6xD(85)(1) <= CNStageIntLLROutputS6xD(132)(1);
  VNStageIntLLRInputS6xD(169)(2) <= CNStageIntLLROutputS6xD(132)(2);
  VNStageIntLLRInputS6xD(225)(2) <= CNStageIntLLROutputS6xD(132)(3);
  VNStageIntLLRInputS6xD(264)(2) <= CNStageIntLLROutputS6xD(132)(4);
  VNStageIntLLRInputS6xD(330)(2) <= CNStageIntLLROutputS6xD(132)(5);
  VNStageIntLLRInputS6xD(8)(1) <= CNStageIntLLROutputS6xD(133)(0);
  VNStageIntLLRInputS6xD(104)(2) <= CNStageIntLLROutputS6xD(133)(1);
  VNStageIntLLRInputS6xD(160)(2) <= CNStageIntLLROutputS6xD(133)(2);
  VNStageIntLLRInputS6xD(199)(2) <= CNStageIntLLROutputS6xD(133)(3);
  VNStageIntLLRInputS6xD(265)(1) <= CNStageIntLLROutputS6xD(133)(4);
  VNStageIntLLRInputS6xD(354)(2) <= CNStageIntLLROutputS6xD(133)(5);
  VNStageIntLLRInputS6xD(7)(2) <= CNStageIntLLROutputS6xD(134)(0);
  VNStageIntLLRInputS6xD(95)(2) <= CNStageIntLLROutputS6xD(134)(1);
  VNStageIntLLRInputS6xD(134)(2) <= CNStageIntLLROutputS6xD(134)(2);
  VNStageIntLLRInputS6xD(200)(2) <= CNStageIntLLROutputS6xD(134)(3);
  VNStageIntLLRInputS6xD(289)(2) <= CNStageIntLLROutputS6xD(134)(4);
  VNStageIntLLRInputS6xD(375)(2) <= CNStageIntLLROutputS6xD(134)(5);
  VNStageIntLLRInputS6xD(6)(2) <= CNStageIntLLROutputS6xD(135)(0);
  VNStageIntLLRInputS6xD(69)(2) <= CNStageIntLLROutputS6xD(135)(1);
  VNStageIntLLRInputS6xD(135)(2) <= CNStageIntLLROutputS6xD(135)(2);
  VNStageIntLLRInputS6xD(224)(2) <= CNStageIntLLROutputS6xD(135)(3);
  VNStageIntLLRInputS6xD(310)(2) <= CNStageIntLLROutputS6xD(135)(4);
  VNStageIntLLRInputS6xD(371)(1) <= CNStageIntLLROutputS6xD(135)(5);
  VNStageIntLLRInputS6xD(5)(2) <= CNStageIntLLROutputS6xD(136)(0);
  VNStageIntLLRInputS6xD(70)(2) <= CNStageIntLLROutputS6xD(136)(1);
  VNStageIntLLRInputS6xD(159)(2) <= CNStageIntLLROutputS6xD(136)(2);
  VNStageIntLLRInputS6xD(245)(2) <= CNStageIntLLROutputS6xD(136)(3);
  VNStageIntLLRInputS6xD(306)(2) <= CNStageIntLLROutputS6xD(136)(4);
  VNStageIntLLRInputS6xD(323)(1) <= CNStageIntLLROutputS6xD(136)(5);
  VNStageIntLLRInputS6xD(3)(1) <= CNStageIntLLROutputS6xD(137)(0);
  VNStageIntLLRInputS6xD(115)(2) <= CNStageIntLLROutputS6xD(137)(1);
  VNStageIntLLRInputS6xD(176)(2) <= CNStageIntLLROutputS6xD(137)(2);
  VNStageIntLLRInputS6xD(193)(2) <= CNStageIntLLROutputS6xD(137)(3);
  VNStageIntLLRInputS6xD(284)(2) <= CNStageIntLLROutputS6xD(137)(4);
  VNStageIntLLRInputS6xD(325)(2) <= CNStageIntLLROutputS6xD(137)(5);
  VNStageIntLLRInputS6xD(2)(2) <= CNStageIntLLROutputS6xD(138)(0);
  VNStageIntLLRInputS6xD(111)(2) <= CNStageIntLLROutputS6xD(138)(1);
  VNStageIntLLRInputS6xD(191)(2) <= CNStageIntLLROutputS6xD(138)(2);
  VNStageIntLLRInputS6xD(219)(2) <= CNStageIntLLROutputS6xD(138)(3);
  VNStageIntLLRInputS6xD(260)(2) <= CNStageIntLLROutputS6xD(138)(4);
  VNStageIntLLRInputS6xD(357)(2) <= CNStageIntLLROutputS6xD(138)(5);
  VNStageIntLLRInputS6xD(1)(1) <= CNStageIntLLROutputS6xD(139)(0);
  VNStageIntLLRInputS6xD(126)(1) <= CNStageIntLLROutputS6xD(139)(1);
  VNStageIntLLRInputS6xD(154)(1) <= CNStageIntLLROutputS6xD(139)(2);
  VNStageIntLLRInputS6xD(195)(1) <= CNStageIntLLROutputS6xD(139)(3);
  VNStageIntLLRInputS6xD(292)(2) <= CNStageIntLLROutputS6xD(139)(4);
  VNStageIntLLRInputS6xD(373)(1) <= CNStageIntLLROutputS6xD(139)(5);
  VNStageIntLLRInputS6xD(63)(2) <= CNStageIntLLROutputS6xD(140)(0);
  VNStageIntLLRInputS6xD(89)(2) <= CNStageIntLLROutputS6xD(140)(1);
  VNStageIntLLRInputS6xD(130)(2) <= CNStageIntLLROutputS6xD(140)(2);
  VNStageIntLLRInputS6xD(227)(2) <= CNStageIntLLROutputS6xD(140)(3);
  VNStageIntLLRInputS6xD(308)(0) <= CNStageIntLLROutputS6xD(140)(4);
  VNStageIntLLRInputS6xD(343)(2) <= CNStageIntLLROutputS6xD(140)(5);
  VNStageIntLLRInputS6xD(62)(1) <= CNStageIntLLROutputS6xD(141)(0);
  VNStageIntLLRInputS6xD(65)(2) <= CNStageIntLLROutputS6xD(141)(1);
  VNStageIntLLRInputS6xD(162)(2) <= CNStageIntLLROutputS6xD(141)(2);
  VNStageIntLLRInputS6xD(243)(2) <= CNStageIntLLROutputS6xD(141)(3);
  VNStageIntLLRInputS6xD(278)(2) <= CNStageIntLLROutputS6xD(141)(4);
  VNStageIntLLRInputS6xD(352)(2) <= CNStageIntLLROutputS6xD(141)(5);
  VNStageIntLLRInputS6xD(61)(1) <= CNStageIntLLROutputS6xD(142)(0);
  VNStageIntLLRInputS6xD(97)(2) <= CNStageIntLLROutputS6xD(142)(1);
  VNStageIntLLRInputS6xD(178)(2) <= CNStageIntLLROutputS6xD(142)(2);
  VNStageIntLLRInputS6xD(213)(2) <= CNStageIntLLROutputS6xD(142)(3);
  VNStageIntLLRInputS6xD(287)(2) <= CNStageIntLLROutputS6xD(142)(4);
  VNStageIntLLRInputS6xD(365)(2) <= CNStageIntLLROutputS6xD(142)(5);
  VNStageIntLLRInputS6xD(60)(1) <= CNStageIntLLROutputS6xD(143)(0);
  VNStageIntLLRInputS6xD(113)(2) <= CNStageIntLLROutputS6xD(143)(1);
  VNStageIntLLRInputS6xD(148)(2) <= CNStageIntLLROutputS6xD(143)(2);
  VNStageIntLLRInputS6xD(222)(1) <= CNStageIntLLROutputS6xD(143)(3);
  VNStageIntLLRInputS6xD(300)(2) <= CNStageIntLLROutputS6xD(143)(4);
  VNStageIntLLRInputS6xD(344)(2) <= CNStageIntLLROutputS6xD(143)(5);
  VNStageIntLLRInputS6xD(59)(0) <= CNStageIntLLROutputS6xD(144)(0);
  VNStageIntLLRInputS6xD(83)(2) <= CNStageIntLLROutputS6xD(144)(1);
  VNStageIntLLRInputS6xD(157)(2) <= CNStageIntLLROutputS6xD(144)(2);
  VNStageIntLLRInputS6xD(235)(1) <= CNStageIntLLROutputS6xD(144)(3);
  VNStageIntLLRInputS6xD(279)(2) <= CNStageIntLLROutputS6xD(144)(4);
  VNStageIntLLRInputS6xD(372)(1) <= CNStageIntLLROutputS6xD(144)(5);
  VNStageIntLLRInputS6xD(58)(1) <= CNStageIntLLROutputS6xD(145)(0);
  VNStageIntLLRInputS6xD(92)(2) <= CNStageIntLLROutputS6xD(145)(1);
  VNStageIntLLRInputS6xD(170)(2) <= CNStageIntLLROutputS6xD(145)(2);
  VNStageIntLLRInputS6xD(214)(2) <= CNStageIntLLROutputS6xD(145)(3);
  VNStageIntLLRInputS6xD(307)(2) <= CNStageIntLLROutputS6xD(145)(4);
  VNStageIntLLRInputS6xD(374)(2) <= CNStageIntLLROutputS6xD(145)(5);
  VNStageIntLLRInputS6xD(57)(1) <= CNStageIntLLROutputS6xD(146)(0);
  VNStageIntLLRInputS6xD(105)(1) <= CNStageIntLLROutputS6xD(146)(1);
  VNStageIntLLRInputS6xD(149)(2) <= CNStageIntLLROutputS6xD(146)(2);
  VNStageIntLLRInputS6xD(242)(2) <= CNStageIntLLROutputS6xD(146)(3);
  VNStageIntLLRInputS6xD(309)(2) <= CNStageIntLLROutputS6xD(146)(4);
  VNStageIntLLRInputS6xD(356)(2) <= CNStageIntLLROutputS6xD(146)(5);
  VNStageIntLLRInputS6xD(56)(2) <= CNStageIntLLROutputS6xD(147)(0);
  VNStageIntLLRInputS6xD(84)(2) <= CNStageIntLLROutputS6xD(147)(1);
  VNStageIntLLRInputS6xD(177)(2) <= CNStageIntLLROutputS6xD(147)(2);
  VNStageIntLLRInputS6xD(244)(0) <= CNStageIntLLROutputS6xD(147)(3);
  VNStageIntLLRInputS6xD(291)(2) <= CNStageIntLLROutputS6xD(147)(4);
  VNStageIntLLRInputS6xD(363)(1) <= CNStageIntLLROutputS6xD(147)(5);
  VNStageIntLLRInputS6xD(55)(2) <= CNStageIntLLROutputS6xD(148)(0);
  VNStageIntLLRInputS6xD(112)(2) <= CNStageIntLLROutputS6xD(148)(1);
  VNStageIntLLRInputS6xD(179)(2) <= CNStageIntLLROutputS6xD(148)(2);
  VNStageIntLLRInputS6xD(226)(1) <= CNStageIntLLROutputS6xD(148)(3);
  VNStageIntLLRInputS6xD(298)(2) <= CNStageIntLLROutputS6xD(148)(4);
  VNStageIntLLRInputS6xD(327)(2) <= CNStageIntLLROutputS6xD(148)(5);
  VNStageIntLLRInputS6xD(54)(2) <= CNStageIntLLROutputS6xD(149)(0);
  VNStageIntLLRInputS6xD(114)(2) <= CNStageIntLLROutputS6xD(149)(1);
  VNStageIntLLRInputS6xD(161)(2) <= CNStageIntLLROutputS6xD(149)(2);
  VNStageIntLLRInputS6xD(233)(2) <= CNStageIntLLROutputS6xD(149)(3);
  VNStageIntLLRInputS6xD(262)(2) <= CNStageIntLLROutputS6xD(149)(4);
  VNStageIntLLRInputS6xD(378)(1) <= CNStageIntLLROutputS6xD(149)(5);
  VNStageIntLLRInputS6xD(53)(1) <= CNStageIntLLROutputS6xD(150)(0);
  VNStageIntLLRInputS6xD(96)(2) <= CNStageIntLLROutputS6xD(150)(1);
  VNStageIntLLRInputS6xD(168)(1) <= CNStageIntLLROutputS6xD(150)(2);
  VNStageIntLLRInputS6xD(197)(2) <= CNStageIntLLROutputS6xD(150)(3);
  VNStageIntLLRInputS6xD(313)(0) <= CNStageIntLLROutputS6xD(150)(4);
  VNStageIntLLRInputS6xD(321)(2) <= CNStageIntLLROutputS6xD(150)(5);
  VNStageIntLLRInputS6xD(52)(1) <= CNStageIntLLROutputS6xD(151)(0);
  VNStageIntLLRInputS6xD(103)(2) <= CNStageIntLLROutputS6xD(151)(1);
  VNStageIntLLRInputS6xD(132)(1) <= CNStageIntLLROutputS6xD(151)(2);
  VNStageIntLLRInputS6xD(248)(2) <= CNStageIntLLROutputS6xD(151)(3);
  VNStageIntLLRInputS6xD(319)(2) <= CNStageIntLLROutputS6xD(151)(4);
  VNStageIntLLRInputS6xD(379)(1) <= CNStageIntLLROutputS6xD(151)(5);
  VNStageIntLLRInputS6xD(50)(2) <= CNStageIntLLROutputS6xD(152)(0);
  VNStageIntLLRInputS6xD(118)(2) <= CNStageIntLLROutputS6xD(152)(1);
  VNStageIntLLRInputS6xD(189)(1) <= CNStageIntLLROutputS6xD(152)(2);
  VNStageIntLLRInputS6xD(249)(0) <= CNStageIntLLROutputS6xD(152)(3);
  VNStageIntLLRInputS6xD(261)(2) <= CNStageIntLLROutputS6xD(152)(4);
  VNStageIntLLRInputS6xD(348)(2) <= CNStageIntLLROutputS6xD(152)(5);
  VNStageIntLLRInputS6xD(49)(2) <= CNStageIntLLROutputS6xD(153)(0);
  VNStageIntLLRInputS6xD(124)(1) <= CNStageIntLLROutputS6xD(153)(1);
  VNStageIntLLRInputS6xD(184)(2) <= CNStageIntLLROutputS6xD(153)(2);
  VNStageIntLLRInputS6xD(196)(2) <= CNStageIntLLROutputS6xD(153)(3);
  VNStageIntLLRInputS6xD(283)(2) <= CNStageIntLLROutputS6xD(153)(4);
  VNStageIntLLRInputS6xD(366)(2) <= CNStageIntLLROutputS6xD(153)(5);
  VNStageIntLLRInputS6xD(48)(1) <= CNStageIntLLROutputS6xD(154)(0);
  VNStageIntLLRInputS6xD(119)(2) <= CNStageIntLLROutputS6xD(154)(1);
  VNStageIntLLRInputS6xD(131)(1) <= CNStageIntLLROutputS6xD(154)(2);
  VNStageIntLLRInputS6xD(218)(2) <= CNStageIntLLROutputS6xD(154)(3);
  VNStageIntLLRInputS6xD(301)(2) <= CNStageIntLLROutputS6xD(154)(4);
  VNStageIntLLRInputS6xD(351)(1) <= CNStageIntLLROutputS6xD(154)(5);
  VNStageIntLLRInputS6xD(47)(1) <= CNStageIntLLROutputS6xD(155)(0);
  VNStageIntLLRInputS6xD(66)(2) <= CNStageIntLLROutputS6xD(155)(1);
  VNStageIntLLRInputS6xD(153)(2) <= CNStageIntLLROutputS6xD(155)(2);
  VNStageIntLLRInputS6xD(236)(2) <= CNStageIntLLROutputS6xD(155)(3);
  VNStageIntLLRInputS6xD(286)(2) <= CNStageIntLLROutputS6xD(155)(4);
  VNStageIntLLRInputS6xD(338)(2) <= CNStageIntLLROutputS6xD(155)(5);
  VNStageIntLLRInputS6xD(46)(2) <= CNStageIntLLROutputS6xD(156)(0);
  VNStageIntLLRInputS6xD(88)(2) <= CNStageIntLLROutputS6xD(156)(1);
  VNStageIntLLRInputS6xD(171)(1) <= CNStageIntLLROutputS6xD(156)(2);
  VNStageIntLLRInputS6xD(221)(2) <= CNStageIntLLROutputS6xD(156)(3);
  VNStageIntLLRInputS6xD(273)(2) <= CNStageIntLLROutputS6xD(156)(4);
  VNStageIntLLRInputS6xD(369)(1) <= CNStageIntLLROutputS6xD(156)(5);
  VNStageIntLLRInputS6xD(45)(2) <= CNStageIntLLROutputS6xD(157)(0);
  VNStageIntLLRInputS6xD(106)(1) <= CNStageIntLLROutputS6xD(157)(1);
  VNStageIntLLRInputS6xD(156)(2) <= CNStageIntLLROutputS6xD(157)(2);
  VNStageIntLLRInputS6xD(208)(2) <= CNStageIntLLROutputS6xD(157)(3);
  VNStageIntLLRInputS6xD(304)(2) <= CNStageIntLLROutputS6xD(157)(4);
  VNStageIntLLRInputS6xD(381)(1) <= CNStageIntLLROutputS6xD(157)(5);
  VNStageIntLLRInputS6xD(44)(2) <= CNStageIntLLROutputS6xD(158)(0);
  VNStageIntLLRInputS6xD(91)(2) <= CNStageIntLLROutputS6xD(158)(1);
  VNStageIntLLRInputS6xD(143)(2) <= CNStageIntLLROutputS6xD(158)(2);
  VNStageIntLLRInputS6xD(239)(2) <= CNStageIntLLROutputS6xD(158)(3);
  VNStageIntLLRInputS6xD(316)(1) <= CNStageIntLLROutputS6xD(158)(4);
  VNStageIntLLRInputS6xD(332)(2) <= CNStageIntLLROutputS6xD(158)(5);
  VNStageIntLLRInputS6xD(43)(1) <= CNStageIntLLROutputS6xD(159)(0);
  VNStageIntLLRInputS6xD(78)(2) <= CNStageIntLLROutputS6xD(159)(1);
  VNStageIntLLRInputS6xD(174)(2) <= CNStageIntLLROutputS6xD(159)(2);
  VNStageIntLLRInputS6xD(251)(1) <= CNStageIntLLROutputS6xD(159)(3);
  VNStageIntLLRInputS6xD(267)(2) <= CNStageIntLLROutputS6xD(159)(4);
  VNStageIntLLRInputS6xD(376)(2) <= CNStageIntLLROutputS6xD(159)(5);
  VNStageIntLLRInputS6xD(42)(2) <= CNStageIntLLROutputS6xD(160)(0);
  VNStageIntLLRInputS6xD(109)(2) <= CNStageIntLLROutputS6xD(160)(1);
  VNStageIntLLRInputS6xD(186)(1) <= CNStageIntLLROutputS6xD(160)(2);
  VNStageIntLLRInputS6xD(202)(2) <= CNStageIntLLROutputS6xD(160)(3);
  VNStageIntLLRInputS6xD(311)(2) <= CNStageIntLLROutputS6xD(160)(4);
  VNStageIntLLRInputS6xD(353)(2) <= CNStageIntLLROutputS6xD(160)(5);
  VNStageIntLLRInputS6xD(41)(2) <= CNStageIntLLROutputS6xD(161)(0);
  VNStageIntLLRInputS6xD(121)(1) <= CNStageIntLLROutputS6xD(161)(1);
  VNStageIntLLRInputS6xD(137)(2) <= CNStageIntLLROutputS6xD(161)(2);
  VNStageIntLLRInputS6xD(246)(2) <= CNStageIntLLROutputS6xD(161)(3);
  VNStageIntLLRInputS6xD(288)(2) <= CNStageIntLLROutputS6xD(161)(4);
  VNStageIntLLRInputS6xD(342)(2) <= CNStageIntLLROutputS6xD(161)(5);
  VNStageIntLLRInputS6xD(40)(2) <= CNStageIntLLROutputS6xD(162)(0);
  VNStageIntLLRInputS6xD(72)(2) <= CNStageIntLLROutputS6xD(162)(1);
  VNStageIntLLRInputS6xD(181)(2) <= CNStageIntLLROutputS6xD(162)(2);
  VNStageIntLLRInputS6xD(223)(2) <= CNStageIntLLROutputS6xD(162)(3);
  VNStageIntLLRInputS6xD(277)(2) <= CNStageIntLLROutputS6xD(162)(4);
  VNStageIntLLRInputS6xD(346)(2) <= CNStageIntLLROutputS6xD(162)(5);
  VNStageIntLLRInputS6xD(39)(2) <= CNStageIntLLROutputS6xD(163)(0);
  VNStageIntLLRInputS6xD(116)(1) <= CNStageIntLLROutputS6xD(163)(1);
  VNStageIntLLRInputS6xD(158)(2) <= CNStageIntLLROutputS6xD(163)(2);
  VNStageIntLLRInputS6xD(212)(2) <= CNStageIntLLROutputS6xD(163)(3);
  VNStageIntLLRInputS6xD(281)(2) <= CNStageIntLLROutputS6xD(163)(4);
  VNStageIntLLRInputS6xD(339)(2) <= CNStageIntLLROutputS6xD(163)(5);
  VNStageIntLLRInputS6xD(38)(2) <= CNStageIntLLROutputS6xD(164)(0);
  VNStageIntLLRInputS6xD(93)(2) <= CNStageIntLLROutputS6xD(164)(1);
  VNStageIntLLRInputS6xD(147)(2) <= CNStageIntLLROutputS6xD(164)(2);
  VNStageIntLLRInputS6xD(216)(2) <= CNStageIntLLROutputS6xD(164)(3);
  VNStageIntLLRInputS6xD(274)(1) <= CNStageIntLLROutputS6xD(164)(4);
  VNStageIntLLRInputS6xD(350)(2) <= CNStageIntLLROutputS6xD(164)(5);
  VNStageIntLLRInputS6xD(37)(2) <= CNStageIntLLROutputS6xD(165)(0);
  VNStageIntLLRInputS6xD(82)(2) <= CNStageIntLLROutputS6xD(165)(1);
  VNStageIntLLRInputS6xD(151)(2) <= CNStageIntLLROutputS6xD(165)(2);
  VNStageIntLLRInputS6xD(209)(2) <= CNStageIntLLROutputS6xD(165)(3);
  VNStageIntLLRInputS6xD(285)(2) <= CNStageIntLLROutputS6xD(165)(4);
  VNStageIntLLRInputS6xD(322)(2) <= CNStageIntLLROutputS6xD(165)(5);
  VNStageIntLLRInputS6xD(36)(2) <= CNStageIntLLROutputS6xD(166)(0);
  VNStageIntLLRInputS6xD(86)(1) <= CNStageIntLLROutputS6xD(166)(1);
  VNStageIntLLRInputS6xD(144)(2) <= CNStageIntLLROutputS6xD(166)(2);
  VNStageIntLLRInputS6xD(220)(2) <= CNStageIntLLROutputS6xD(166)(3);
  VNStageIntLLRInputS6xD(257)(2) <= CNStageIntLLROutputS6xD(166)(4);
  VNStageIntLLRInputS6xD(377)(1) <= CNStageIntLLROutputS6xD(166)(5);
  VNStageIntLLRInputS6xD(35)(2) <= CNStageIntLLROutputS6xD(167)(0);
  VNStageIntLLRInputS6xD(79)(2) <= CNStageIntLLROutputS6xD(167)(1);
  VNStageIntLLRInputS6xD(155)(2) <= CNStageIntLLROutputS6xD(167)(2);
  VNStageIntLLRInputS6xD(255)(2) <= CNStageIntLLROutputS6xD(167)(3);
  VNStageIntLLRInputS6xD(312)(2) <= CNStageIntLLROutputS6xD(167)(4);
  VNStageIntLLRInputS6xD(331)(2) <= CNStageIntLLROutputS6xD(167)(5);
  VNStageIntLLRInputS6xD(34)(2) <= CNStageIntLLROutputS6xD(168)(0);
  VNStageIntLLRInputS6xD(90)(2) <= CNStageIntLLROutputS6xD(168)(1);
  VNStageIntLLRInputS6xD(190)(0) <= CNStageIntLLROutputS6xD(168)(2);
  VNStageIntLLRInputS6xD(247)(2) <= CNStageIntLLROutputS6xD(168)(3);
  VNStageIntLLRInputS6xD(266)(1) <= CNStageIntLLROutputS6xD(168)(4);
  VNStageIntLLRInputS6xD(328)(2) <= CNStageIntLLROutputS6xD(168)(5);
  VNStageIntLLRInputS6xD(33)(2) <= CNStageIntLLROutputS6xD(169)(0);
  VNStageIntLLRInputS6xD(125)(1) <= CNStageIntLLROutputS6xD(169)(1);
  VNStageIntLLRInputS6xD(182)(2) <= CNStageIntLLROutputS6xD(169)(2);
  VNStageIntLLRInputS6xD(201)(2) <= CNStageIntLLROutputS6xD(169)(3);
  VNStageIntLLRInputS6xD(263)(2) <= CNStageIntLLROutputS6xD(169)(4);
  VNStageIntLLRInputS6xD(362)(2) <= CNStageIntLLROutputS6xD(169)(5);
  VNStageIntLLRInputS6xD(0)(2) <= CNStageIntLLROutputS6xD(170)(0);
  VNStageIntLLRInputS6xD(75)(2) <= CNStageIntLLROutputS6xD(170)(1);
  VNStageIntLLRInputS6xD(140)(2) <= CNStageIntLLROutputS6xD(170)(2);
  VNStageIntLLRInputS6xD(205)(0) <= CNStageIntLLROutputS6xD(170)(3);
  VNStageIntLLRInputS6xD(270)(2) <= CNStageIntLLROutputS6xD(170)(4);
  VNStageIntLLRInputS6xD(335)(2) <= CNStageIntLLROutputS6xD(170)(5);
  VNStageIntLLRInputS6xD(62)(2) <= CNStageIntLLROutputS6xD(171)(0);
  VNStageIntLLRInputS6xD(109)(3) <= CNStageIntLLROutputS6xD(171)(1);
  VNStageIntLLRInputS6xD(161)(3) <= CNStageIntLLROutputS6xD(171)(2);
  VNStageIntLLRInputS6xD(194)(3) <= CNStageIntLLROutputS6xD(171)(3);
  VNStageIntLLRInputS6xD(271)(2) <= CNStageIntLLROutputS6xD(171)(4);
  VNStageIntLLRInputS6xD(350)(3) <= CNStageIntLLROutputS6xD(171)(5);
  VNStageIntLLRInputS6xD(61)(2) <= CNStageIntLLROutputS6xD(172)(0);
  VNStageIntLLRInputS6xD(96)(3) <= CNStageIntLLROutputS6xD(172)(1);
  VNStageIntLLRInputS6xD(129)(3) <= CNStageIntLLROutputS6xD(172)(2);
  VNStageIntLLRInputS6xD(206)(2) <= CNStageIntLLROutputS6xD(172)(3);
  VNStageIntLLRInputS6xD(285)(3) <= CNStageIntLLROutputS6xD(172)(4);
  VNStageIntLLRInputS6xD(331)(3) <= CNStageIntLLROutputS6xD(172)(5);
  VNStageIntLLRInputS6xD(60)(2) <= CNStageIntLLROutputS6xD(173)(0);
  VNStageIntLLRInputS6xD(127)(3) <= CNStageIntLLROutputS6xD(173)(1);
  VNStageIntLLRInputS6xD(141)(1) <= CNStageIntLLROutputS6xD(173)(2);
  VNStageIntLLRInputS6xD(220)(3) <= CNStageIntLLROutputS6xD(173)(3);
  VNStageIntLLRInputS6xD(266)(2) <= CNStageIntLLROutputS6xD(173)(4);
  VNStageIntLLRInputS6xD(371)(2) <= CNStageIntLLROutputS6xD(173)(5);
  VNStageIntLLRInputS6xD(59)(1) <= CNStageIntLLROutputS6xD(174)(0);
  VNStageIntLLRInputS6xD(76)(3) <= CNStageIntLLROutputS6xD(174)(1);
  VNStageIntLLRInputS6xD(155)(3) <= CNStageIntLLROutputS6xD(174)(2);
  VNStageIntLLRInputS6xD(201)(3) <= CNStageIntLLROutputS6xD(174)(3);
  VNStageIntLLRInputS6xD(306)(3) <= CNStageIntLLROutputS6xD(174)(4);
  VNStageIntLLRInputS6xD(360)(3) <= CNStageIntLLROutputS6xD(174)(5);
  VNStageIntLLRInputS6xD(58)(2) <= CNStageIntLLROutputS6xD(175)(0);
  VNStageIntLLRInputS6xD(90)(3) <= CNStageIntLLROutputS6xD(175)(1);
  VNStageIntLLRInputS6xD(136)(3) <= CNStageIntLLROutputS6xD(175)(2);
  VNStageIntLLRInputS6xD(241)(2) <= CNStageIntLLROutputS6xD(175)(3);
  VNStageIntLLRInputS6xD(295)(3) <= CNStageIntLLROutputS6xD(175)(4);
  VNStageIntLLRInputS6xD(364)(3) <= CNStageIntLLROutputS6xD(175)(5);
  VNStageIntLLRInputS6xD(57)(2) <= CNStageIntLLROutputS6xD(176)(0);
  VNStageIntLLRInputS6xD(71)(2) <= CNStageIntLLROutputS6xD(176)(1);
  VNStageIntLLRInputS6xD(176)(3) <= CNStageIntLLROutputS6xD(176)(2);
  VNStageIntLLRInputS6xD(230)(2) <= CNStageIntLLROutputS6xD(176)(3);
  VNStageIntLLRInputS6xD(299)(2) <= CNStageIntLLROutputS6xD(176)(4);
  VNStageIntLLRInputS6xD(357)(3) <= CNStageIntLLROutputS6xD(176)(5);
  VNStageIntLLRInputS6xD(56)(3) <= CNStageIntLLROutputS6xD(177)(0);
  VNStageIntLLRInputS6xD(111)(3) <= CNStageIntLLROutputS6xD(177)(1);
  VNStageIntLLRInputS6xD(165)(3) <= CNStageIntLLROutputS6xD(177)(2);
  VNStageIntLLRInputS6xD(234)(3) <= CNStageIntLLROutputS6xD(177)(3);
  VNStageIntLLRInputS6xD(292)(3) <= CNStageIntLLROutputS6xD(177)(4);
  VNStageIntLLRInputS6xD(368)(1) <= CNStageIntLLROutputS6xD(177)(5);
  VNStageIntLLRInputS6xD(55)(3) <= CNStageIntLLROutputS6xD(178)(0);
  VNStageIntLLRInputS6xD(100)(3) <= CNStageIntLLROutputS6xD(178)(1);
  VNStageIntLLRInputS6xD(169)(3) <= CNStageIntLLROutputS6xD(178)(2);
  VNStageIntLLRInputS6xD(227)(3) <= CNStageIntLLROutputS6xD(178)(3);
  VNStageIntLLRInputS6xD(303)(3) <= CNStageIntLLROutputS6xD(178)(4);
  VNStageIntLLRInputS6xD(340)(3) <= CNStageIntLLROutputS6xD(178)(5);
  VNStageIntLLRInputS6xD(54)(3) <= CNStageIntLLROutputS6xD(179)(0);
  VNStageIntLLRInputS6xD(104)(3) <= CNStageIntLLROutputS6xD(179)(1);
  VNStageIntLLRInputS6xD(162)(3) <= CNStageIntLLROutputS6xD(179)(2);
  VNStageIntLLRInputS6xD(238)(3) <= CNStageIntLLROutputS6xD(179)(3);
  VNStageIntLLRInputS6xD(275)(3) <= CNStageIntLLROutputS6xD(179)(4);
  VNStageIntLLRInputS6xD(332)(3) <= CNStageIntLLROutputS6xD(179)(5);
  VNStageIntLLRInputS6xD(53)(2) <= CNStageIntLLROutputS6xD(180)(0);
  VNStageIntLLRInputS6xD(97)(3) <= CNStageIntLLROutputS6xD(180)(1);
  VNStageIntLLRInputS6xD(173)(3) <= CNStageIntLLROutputS6xD(180)(2);
  VNStageIntLLRInputS6xD(210)(3) <= CNStageIntLLROutputS6xD(180)(3);
  VNStageIntLLRInputS6xD(267)(3) <= CNStageIntLLROutputS6xD(180)(4);
  VNStageIntLLRInputS6xD(349)(2) <= CNStageIntLLROutputS6xD(180)(5);
  VNStageIntLLRInputS6xD(52)(2) <= CNStageIntLLROutputS6xD(181)(0);
  VNStageIntLLRInputS6xD(108)(3) <= CNStageIntLLROutputS6xD(181)(1);
  VNStageIntLLRInputS6xD(145)(3) <= CNStageIntLLROutputS6xD(181)(2);
  VNStageIntLLRInputS6xD(202)(3) <= CNStageIntLLROutputS6xD(181)(3);
  VNStageIntLLRInputS6xD(284)(3) <= CNStageIntLLROutputS6xD(181)(4);
  VNStageIntLLRInputS6xD(346)(3) <= CNStageIntLLROutputS6xD(181)(5);
  VNStageIntLLRInputS6xD(51)(2) <= CNStageIntLLROutputS6xD(182)(0);
  VNStageIntLLRInputS6xD(80)(3) <= CNStageIntLLROutputS6xD(182)(1);
  VNStageIntLLRInputS6xD(137)(3) <= CNStageIntLLROutputS6xD(182)(2);
  VNStageIntLLRInputS6xD(219)(3) <= CNStageIntLLROutputS6xD(182)(3);
  VNStageIntLLRInputS6xD(281)(3) <= CNStageIntLLROutputS6xD(182)(4);
  VNStageIntLLRInputS6xD(380)(2) <= CNStageIntLLROutputS6xD(182)(5);
  VNStageIntLLRInputS6xD(50)(3) <= CNStageIntLLROutputS6xD(183)(0);
  VNStageIntLLRInputS6xD(72)(3) <= CNStageIntLLROutputS6xD(183)(1);
  VNStageIntLLRInputS6xD(154)(2) <= CNStageIntLLROutputS6xD(183)(2);
  VNStageIntLLRInputS6xD(216)(3) <= CNStageIntLLROutputS6xD(183)(3);
  VNStageIntLLRInputS6xD(315)(2) <= CNStageIntLLROutputS6xD(183)(4);
  VNStageIntLLRInputS6xD(337)(3) <= CNStageIntLLROutputS6xD(183)(5);
  VNStageIntLLRInputS6xD(49)(3) <= CNStageIntLLROutputS6xD(184)(0);
  VNStageIntLLRInputS6xD(89)(3) <= CNStageIntLLROutputS6xD(184)(1);
  VNStageIntLLRInputS6xD(151)(3) <= CNStageIntLLROutputS6xD(184)(2);
  VNStageIntLLRInputS6xD(250)(2) <= CNStageIntLLROutputS6xD(184)(3);
  VNStageIntLLRInputS6xD(272)(3) <= CNStageIntLLROutputS6xD(184)(4);
  VNStageIntLLRInputS6xD(323)(2) <= CNStageIntLLROutputS6xD(184)(5);
  VNStageIntLLRInputS6xD(46)(3) <= CNStageIntLLROutputS6xD(185)(0);
  VNStageIntLLRInputS6xD(77)(1) <= CNStageIntLLROutputS6xD(185)(1);
  VNStageIntLLRInputS6xD(191)(3) <= CNStageIntLLROutputS6xD(185)(2);
  VNStageIntLLRInputS6xD(246)(3) <= CNStageIntLLROutputS6xD(185)(3);
  VNStageIntLLRInputS6xD(277)(3) <= CNStageIntLLROutputS6xD(185)(4);
  VNStageIntLLRInputS6xD(325)(3) <= CNStageIntLLROutputS6xD(185)(5);
  VNStageIntLLRInputS6xD(45)(3) <= CNStageIntLLROutputS6xD(186)(0);
  VNStageIntLLRInputS6xD(126)(2) <= CNStageIntLLROutputS6xD(186)(1);
  VNStageIntLLRInputS6xD(181)(3) <= CNStageIntLLROutputS6xD(186)(2);
  VNStageIntLLRInputS6xD(212)(3) <= CNStageIntLLROutputS6xD(186)(3);
  VNStageIntLLRInputS6xD(260)(3) <= CNStageIntLLROutputS6xD(186)(4);
  VNStageIntLLRInputS6xD(355)(3) <= CNStageIntLLROutputS6xD(186)(5);
  VNStageIntLLRInputS6xD(44)(3) <= CNStageIntLLROutputS6xD(187)(0);
  VNStageIntLLRInputS6xD(116)(2) <= CNStageIntLLROutputS6xD(187)(1);
  VNStageIntLLRInputS6xD(147)(3) <= CNStageIntLLROutputS6xD(187)(2);
  VNStageIntLLRInputS6xD(195)(2) <= CNStageIntLLROutputS6xD(187)(3);
  VNStageIntLLRInputS6xD(290)(3) <= CNStageIntLLROutputS6xD(187)(4);
  VNStageIntLLRInputS6xD(378)(2) <= CNStageIntLLROutputS6xD(187)(5);
  VNStageIntLLRInputS6xD(43)(2) <= CNStageIntLLROutputS6xD(188)(0);
  VNStageIntLLRInputS6xD(82)(3) <= CNStageIntLLROutputS6xD(188)(1);
  VNStageIntLLRInputS6xD(130)(3) <= CNStageIntLLROutputS6xD(188)(2);
  VNStageIntLLRInputS6xD(225)(3) <= CNStageIntLLROutputS6xD(188)(3);
  VNStageIntLLRInputS6xD(313)(1) <= CNStageIntLLROutputS6xD(188)(4);
  VNStageIntLLRInputS6xD(351)(2) <= CNStageIntLLROutputS6xD(188)(5);
  VNStageIntLLRInputS6xD(42)(3) <= CNStageIntLLROutputS6xD(189)(0);
  VNStageIntLLRInputS6xD(65)(3) <= CNStageIntLLROutputS6xD(189)(1);
  VNStageIntLLRInputS6xD(160)(3) <= CNStageIntLLROutputS6xD(189)(2);
  VNStageIntLLRInputS6xD(248)(3) <= CNStageIntLLROutputS6xD(189)(3);
  VNStageIntLLRInputS6xD(286)(3) <= CNStageIntLLROutputS6xD(189)(4);
  VNStageIntLLRInputS6xD(335)(3) <= CNStageIntLLROutputS6xD(189)(5);
  VNStageIntLLRInputS6xD(41)(3) <= CNStageIntLLROutputS6xD(190)(0);
  VNStageIntLLRInputS6xD(95)(3) <= CNStageIntLLROutputS6xD(190)(1);
  VNStageIntLLRInputS6xD(183)(2) <= CNStageIntLLROutputS6xD(190)(2);
  VNStageIntLLRInputS6xD(221)(3) <= CNStageIntLLROutputS6xD(190)(3);
  VNStageIntLLRInputS6xD(270)(3) <= CNStageIntLLROutputS6xD(190)(4);
  VNStageIntLLRInputS6xD(338)(3) <= CNStageIntLLROutputS6xD(190)(5);
  VNStageIntLLRInputS6xD(39)(3) <= CNStageIntLLROutputS6xD(191)(0);
  VNStageIntLLRInputS6xD(91)(3) <= CNStageIntLLROutputS6xD(191)(1);
  VNStageIntLLRInputS6xD(140)(3) <= CNStageIntLLROutputS6xD(191)(2);
  VNStageIntLLRInputS6xD(208)(3) <= CNStageIntLLROutputS6xD(191)(3);
  VNStageIntLLRInputS6xD(314)(0) <= CNStageIntLLROutputS6xD(191)(4);
  VNStageIntLLRInputS6xD(354)(3) <= CNStageIntLLROutputS6xD(191)(5);
  VNStageIntLLRInputS6xD(38)(3) <= CNStageIntLLROutputS6xD(192)(0);
  VNStageIntLLRInputS6xD(75)(3) <= CNStageIntLLROutputS6xD(192)(1);
  VNStageIntLLRInputS6xD(143)(3) <= CNStageIntLLROutputS6xD(192)(2);
  VNStageIntLLRInputS6xD(249)(1) <= CNStageIntLLROutputS6xD(192)(3);
  VNStageIntLLRInputS6xD(289)(3) <= CNStageIntLLROutputS6xD(192)(4);
  VNStageIntLLRInputS6xD(352)(3) <= CNStageIntLLROutputS6xD(192)(5);
  VNStageIntLLRInputS6xD(37)(3) <= CNStageIntLLROutputS6xD(193)(0);
  VNStageIntLLRInputS6xD(78)(3) <= CNStageIntLLROutputS6xD(193)(1);
  VNStageIntLLRInputS6xD(184)(3) <= CNStageIntLLROutputS6xD(193)(2);
  VNStageIntLLRInputS6xD(224)(3) <= CNStageIntLLROutputS6xD(193)(3);
  VNStageIntLLRInputS6xD(287)(3) <= CNStageIntLLROutputS6xD(193)(4);
  VNStageIntLLRInputS6xD(377)(2) <= CNStageIntLLROutputS6xD(193)(5);
  VNStageIntLLRInputS6xD(35)(3) <= CNStageIntLLROutputS6xD(194)(0);
  VNStageIntLLRInputS6xD(94)(2) <= CNStageIntLLROutputS6xD(194)(1);
  VNStageIntLLRInputS6xD(157)(3) <= CNStageIntLLROutputS6xD(194)(2);
  VNStageIntLLRInputS6xD(247)(3) <= CNStageIntLLROutputS6xD(194)(3);
  VNStageIntLLRInputS6xD(257)(3) <= CNStageIntLLROutputS6xD(194)(4);
  VNStageIntLLRInputS6xD(365)(3) <= CNStageIntLLROutputS6xD(194)(5);
  VNStageIntLLRInputS6xD(34)(3) <= CNStageIntLLROutputS6xD(195)(0);
  VNStageIntLLRInputS6xD(92)(3) <= CNStageIntLLROutputS6xD(195)(1);
  VNStageIntLLRInputS6xD(182)(3) <= CNStageIntLLROutputS6xD(195)(2);
  VNStageIntLLRInputS6xD(255)(3) <= CNStageIntLLROutputS6xD(195)(3);
  VNStageIntLLRInputS6xD(300)(3) <= CNStageIntLLROutputS6xD(195)(4);
  VNStageIntLLRInputS6xD(359)(3) <= CNStageIntLLROutputS6xD(195)(5);
  VNStageIntLLRInputS6xD(33)(3) <= CNStageIntLLROutputS6xD(196)(0);
  VNStageIntLLRInputS6xD(117)(3) <= CNStageIntLLROutputS6xD(196)(1);
  VNStageIntLLRInputS6xD(190)(1) <= CNStageIntLLROutputS6xD(196)(2);
  VNStageIntLLRInputS6xD(235)(2) <= CNStageIntLLROutputS6xD(196)(3);
  VNStageIntLLRInputS6xD(294)(3) <= CNStageIntLLROutputS6xD(196)(4);
  VNStageIntLLRInputS6xD(320)(2) <= CNStageIntLLROutputS6xD(196)(5);
  VNStageIntLLRInputS6xD(31)(2) <= CNStageIntLLROutputS6xD(197)(0);
  VNStageIntLLRInputS6xD(105)(2) <= CNStageIntLLROutputS6xD(197)(1);
  VNStageIntLLRInputS6xD(164)(3) <= CNStageIntLLROutputS6xD(197)(2);
  VNStageIntLLRInputS6xD(192)(3) <= CNStageIntLLROutputS6xD(197)(3);
  VNStageIntLLRInputS6xD(293)(3) <= CNStageIntLLROutputS6xD(197)(4);
  VNStageIntLLRInputS6xD(363)(2) <= CNStageIntLLROutputS6xD(197)(5);
  VNStageIntLLRInputS6xD(30)(3) <= CNStageIntLLROutputS6xD(198)(0);
  VNStageIntLLRInputS6xD(99)(3) <= CNStageIntLLROutputS6xD(198)(1);
  VNStageIntLLRInputS6xD(128)(3) <= CNStageIntLLROutputS6xD(198)(2);
  VNStageIntLLRInputS6xD(228)(3) <= CNStageIntLLROutputS6xD(198)(3);
  VNStageIntLLRInputS6xD(298)(3) <= CNStageIntLLROutputS6xD(198)(4);
  VNStageIntLLRInputS6xD(382)(2) <= CNStageIntLLROutputS6xD(198)(5);
  VNStageIntLLRInputS6xD(28)(3) <= CNStageIntLLROutputS6xD(199)(0);
  VNStageIntLLRInputS6xD(98)(2) <= CNStageIntLLROutputS6xD(199)(1);
  VNStageIntLLRInputS6xD(168)(2) <= CNStageIntLLROutputS6xD(199)(2);
  VNStageIntLLRInputS6xD(252)(2) <= CNStageIntLLROutputS6xD(199)(3);
  VNStageIntLLRInputS6xD(308)(1) <= CNStageIntLLROutputS6xD(199)(4);
  VNStageIntLLRInputS6xD(347)(3) <= CNStageIntLLROutputS6xD(199)(5);
  VNStageIntLLRInputS6xD(27)(3) <= CNStageIntLLROutputS6xD(200)(0);
  VNStageIntLLRInputS6xD(103)(3) <= CNStageIntLLROutputS6xD(200)(1);
  VNStageIntLLRInputS6xD(187)(2) <= CNStageIntLLROutputS6xD(200)(2);
  VNStageIntLLRInputS6xD(243)(3) <= CNStageIntLLROutputS6xD(200)(3);
  VNStageIntLLRInputS6xD(282)(3) <= CNStageIntLLROutputS6xD(200)(4);
  VNStageIntLLRInputS6xD(348)(3) <= CNStageIntLLROutputS6xD(200)(5);
  VNStageIntLLRInputS6xD(26)(3) <= CNStageIntLLROutputS6xD(201)(0);
  VNStageIntLLRInputS6xD(122)(2) <= CNStageIntLLROutputS6xD(201)(1);
  VNStageIntLLRInputS6xD(178)(3) <= CNStageIntLLROutputS6xD(201)(2);
  VNStageIntLLRInputS6xD(217)(3) <= CNStageIntLLROutputS6xD(201)(3);
  VNStageIntLLRInputS6xD(283)(3) <= CNStageIntLLROutputS6xD(201)(4);
  VNStageIntLLRInputS6xD(372)(2) <= CNStageIntLLROutputS6xD(201)(5);
  VNStageIntLLRInputS6xD(25)(3) <= CNStageIntLLROutputS6xD(202)(0);
  VNStageIntLLRInputS6xD(113)(3) <= CNStageIntLLROutputS6xD(202)(1);
  VNStageIntLLRInputS6xD(152)(3) <= CNStageIntLLROutputS6xD(202)(2);
  VNStageIntLLRInputS6xD(218)(3) <= CNStageIntLLROutputS6xD(202)(3);
  VNStageIntLLRInputS6xD(307)(3) <= CNStageIntLLROutputS6xD(202)(4);
  VNStageIntLLRInputS6xD(330)(3) <= CNStageIntLLROutputS6xD(202)(5);
  VNStageIntLLRInputS6xD(24)(3) <= CNStageIntLLROutputS6xD(203)(0);
  VNStageIntLLRInputS6xD(87)(3) <= CNStageIntLLROutputS6xD(203)(1);
  VNStageIntLLRInputS6xD(153)(3) <= CNStageIntLLROutputS6xD(203)(2);
  VNStageIntLLRInputS6xD(242)(3) <= CNStageIntLLROutputS6xD(203)(3);
  VNStageIntLLRInputS6xD(265)(2) <= CNStageIntLLROutputS6xD(203)(4);
  VNStageIntLLRInputS6xD(326)(2) <= CNStageIntLLROutputS6xD(203)(5);
  VNStageIntLLRInputS6xD(23)(3) <= CNStageIntLLROutputS6xD(204)(0);
  VNStageIntLLRInputS6xD(88)(3) <= CNStageIntLLROutputS6xD(204)(1);
  VNStageIntLLRInputS6xD(177)(3) <= CNStageIntLLROutputS6xD(204)(2);
  VNStageIntLLRInputS6xD(200)(3) <= CNStageIntLLROutputS6xD(204)(3);
  VNStageIntLLRInputS6xD(261)(3) <= CNStageIntLLROutputS6xD(204)(4);
  VNStageIntLLRInputS6xD(341)(3) <= CNStageIntLLROutputS6xD(204)(5);
  VNStageIntLLRInputS6xD(22)(3) <= CNStageIntLLROutputS6xD(205)(0);
  VNStageIntLLRInputS6xD(112)(3) <= CNStageIntLLROutputS6xD(205)(1);
  VNStageIntLLRInputS6xD(135)(3) <= CNStageIntLLROutputS6xD(205)(2);
  VNStageIntLLRInputS6xD(196)(3) <= CNStageIntLLROutputS6xD(205)(3);
  VNStageIntLLRInputS6xD(276)(3) <= CNStageIntLLROutputS6xD(205)(4);
  VNStageIntLLRInputS6xD(367)(3) <= CNStageIntLLROutputS6xD(205)(5);
  VNStageIntLLRInputS6xD(21)(3) <= CNStageIntLLROutputS6xD(206)(0);
  VNStageIntLLRInputS6xD(70)(3) <= CNStageIntLLROutputS6xD(206)(1);
  VNStageIntLLRInputS6xD(131)(2) <= CNStageIntLLROutputS6xD(206)(2);
  VNStageIntLLRInputS6xD(211)(3) <= CNStageIntLLROutputS6xD(206)(3);
  VNStageIntLLRInputS6xD(302)(3) <= CNStageIntLLROutputS6xD(206)(4);
  VNStageIntLLRInputS6xD(343)(3) <= CNStageIntLLROutputS6xD(206)(5);
  VNStageIntLLRInputS6xD(18)(3) <= CNStageIntLLROutputS6xD(207)(0);
  VNStageIntLLRInputS6xD(107)(2) <= CNStageIntLLROutputS6xD(207)(1);
  VNStageIntLLRInputS6xD(148)(3) <= CNStageIntLLROutputS6xD(207)(2);
  VNStageIntLLRInputS6xD(245)(3) <= CNStageIntLLROutputS6xD(207)(3);
  VNStageIntLLRInputS6xD(263)(3) <= CNStageIntLLROutputS6xD(207)(4);
  VNStageIntLLRInputS6xD(361)(3) <= CNStageIntLLROutputS6xD(207)(5);
  VNStageIntLLRInputS6xD(17)(3) <= CNStageIntLLROutputS6xD(208)(0);
  VNStageIntLLRInputS6xD(83)(3) <= CNStageIntLLROutputS6xD(208)(1);
  VNStageIntLLRInputS6xD(180)(1) <= CNStageIntLLROutputS6xD(208)(2);
  VNStageIntLLRInputS6xD(198)(3) <= CNStageIntLLROutputS6xD(208)(3);
  VNStageIntLLRInputS6xD(296)(3) <= CNStageIntLLROutputS6xD(208)(4);
  VNStageIntLLRInputS6xD(370)(2) <= CNStageIntLLROutputS6xD(208)(5);
  VNStageIntLLRInputS6xD(16)(2) <= CNStageIntLLROutputS6xD(209)(0);
  VNStageIntLLRInputS6xD(115)(3) <= CNStageIntLLROutputS6xD(209)(1);
  VNStageIntLLRInputS6xD(133)(1) <= CNStageIntLLROutputS6xD(209)(2);
  VNStageIntLLRInputS6xD(231)(2) <= CNStageIntLLROutputS6xD(209)(3);
  VNStageIntLLRInputS6xD(305)(3) <= CNStageIntLLROutputS6xD(209)(4);
  VNStageIntLLRInputS6xD(383)(3) <= CNStageIntLLROutputS6xD(209)(5);
  VNStageIntLLRInputS6xD(15)(3) <= CNStageIntLLROutputS6xD(210)(0);
  VNStageIntLLRInputS6xD(68)(2) <= CNStageIntLLROutputS6xD(210)(1);
  VNStageIntLLRInputS6xD(166)(3) <= CNStageIntLLROutputS6xD(210)(2);
  VNStageIntLLRInputS6xD(240)(3) <= CNStageIntLLROutputS6xD(210)(3);
  VNStageIntLLRInputS6xD(318)(1) <= CNStageIntLLROutputS6xD(210)(4);
  VNStageIntLLRInputS6xD(362)(3) <= CNStageIntLLROutputS6xD(210)(5);
  VNStageIntLLRInputS6xD(14)(3) <= CNStageIntLLROutputS6xD(211)(0);
  VNStageIntLLRInputS6xD(101)(3) <= CNStageIntLLROutputS6xD(211)(1);
  VNStageIntLLRInputS6xD(175)(3) <= CNStageIntLLROutputS6xD(211)(2);
  VNStageIntLLRInputS6xD(253)(2) <= CNStageIntLLROutputS6xD(211)(3);
  VNStageIntLLRInputS6xD(297)(3) <= CNStageIntLLROutputS6xD(211)(4);
  VNStageIntLLRInputS6xD(327)(3) <= CNStageIntLLROutputS6xD(211)(5);
  VNStageIntLLRInputS6xD(13)(2) <= CNStageIntLLROutputS6xD(212)(0);
  VNStageIntLLRInputS6xD(110)(3) <= CNStageIntLLROutputS6xD(212)(1);
  VNStageIntLLRInputS6xD(188)(1) <= CNStageIntLLROutputS6xD(212)(2);
  VNStageIntLLRInputS6xD(232)(2) <= CNStageIntLLROutputS6xD(212)(3);
  VNStageIntLLRInputS6xD(262)(3) <= CNStageIntLLROutputS6xD(212)(4);
  VNStageIntLLRInputS6xD(329)(3) <= CNStageIntLLROutputS6xD(212)(5);
  VNStageIntLLRInputS6xD(12)(3) <= CNStageIntLLROutputS6xD(213)(0);
  VNStageIntLLRInputS6xD(123)(2) <= CNStageIntLLROutputS6xD(213)(1);
  VNStageIntLLRInputS6xD(167)(3) <= CNStageIntLLROutputS6xD(213)(2);
  VNStageIntLLRInputS6xD(197)(3) <= CNStageIntLLROutputS6xD(213)(3);
  VNStageIntLLRInputS6xD(264)(3) <= CNStageIntLLROutputS6xD(213)(4);
  VNStageIntLLRInputS6xD(374)(3) <= CNStageIntLLROutputS6xD(213)(5);
  VNStageIntLLRInputS6xD(11)(3) <= CNStageIntLLROutputS6xD(214)(0);
  VNStageIntLLRInputS6xD(102)(3) <= CNStageIntLLROutputS6xD(214)(1);
  VNStageIntLLRInputS6xD(132)(2) <= CNStageIntLLROutputS6xD(214)(2);
  VNStageIntLLRInputS6xD(199)(3) <= CNStageIntLLROutputS6xD(214)(3);
  VNStageIntLLRInputS6xD(309)(3) <= CNStageIntLLROutputS6xD(214)(4);
  VNStageIntLLRInputS6xD(381)(2) <= CNStageIntLLROutputS6xD(214)(5);
  VNStageIntLLRInputS6xD(9)(3) <= CNStageIntLLROutputS6xD(215)(0);
  VNStageIntLLRInputS6xD(69)(3) <= CNStageIntLLROutputS6xD(215)(1);
  VNStageIntLLRInputS6xD(179)(3) <= CNStageIntLLROutputS6xD(215)(2);
  VNStageIntLLRInputS6xD(251)(2) <= CNStageIntLLROutputS6xD(215)(3);
  VNStageIntLLRInputS6xD(280)(3) <= CNStageIntLLROutputS6xD(215)(4);
  VNStageIntLLRInputS6xD(333)(2) <= CNStageIntLLROutputS6xD(215)(5);
  VNStageIntLLRInputS6xD(8)(2) <= CNStageIntLLROutputS6xD(216)(0);
  VNStageIntLLRInputS6xD(114)(3) <= CNStageIntLLROutputS6xD(216)(1);
  VNStageIntLLRInputS6xD(186)(2) <= CNStageIntLLROutputS6xD(216)(2);
  VNStageIntLLRInputS6xD(215)(3) <= CNStageIntLLROutputS6xD(216)(3);
  VNStageIntLLRInputS6xD(268)(3) <= CNStageIntLLROutputS6xD(216)(4);
  VNStageIntLLRInputS6xD(339)(3) <= CNStageIntLLROutputS6xD(216)(5);
  VNStageIntLLRInputS6xD(7)(3) <= CNStageIntLLROutputS6xD(217)(0);
  VNStageIntLLRInputS6xD(121)(2) <= CNStageIntLLROutputS6xD(217)(1);
  VNStageIntLLRInputS6xD(150)(3) <= CNStageIntLLROutputS6xD(217)(2);
  VNStageIntLLRInputS6xD(203)(3) <= CNStageIntLLROutputS6xD(217)(3);
  VNStageIntLLRInputS6xD(274)(2) <= CNStageIntLLROutputS6xD(217)(4);
  VNStageIntLLRInputS6xD(334)(2) <= CNStageIntLLROutputS6xD(217)(5);
  VNStageIntLLRInputS6xD(6)(3) <= CNStageIntLLROutputS6xD(218)(0);
  VNStageIntLLRInputS6xD(85)(2) <= CNStageIntLLROutputS6xD(218)(1);
  VNStageIntLLRInputS6xD(138)(3) <= CNStageIntLLROutputS6xD(218)(2);
  VNStageIntLLRInputS6xD(209)(3) <= CNStageIntLLROutputS6xD(218)(3);
  VNStageIntLLRInputS6xD(269)(2) <= CNStageIntLLROutputS6xD(218)(4);
  VNStageIntLLRInputS6xD(344)(3) <= CNStageIntLLROutputS6xD(218)(5);
  VNStageIntLLRInputS6xD(5)(3) <= CNStageIntLLROutputS6xD(219)(0);
  VNStageIntLLRInputS6xD(73)(3) <= CNStageIntLLROutputS6xD(219)(1);
  VNStageIntLLRInputS6xD(144)(3) <= CNStageIntLLROutputS6xD(219)(2);
  VNStageIntLLRInputS6xD(204)(3) <= CNStageIntLLROutputS6xD(219)(3);
  VNStageIntLLRInputS6xD(279)(3) <= CNStageIntLLROutputS6xD(219)(4);
  VNStageIntLLRInputS6xD(366)(3) <= CNStageIntLLROutputS6xD(219)(5);
  VNStageIntLLRInputS6xD(4)(2) <= CNStageIntLLROutputS6xD(220)(0);
  VNStageIntLLRInputS6xD(79)(3) <= CNStageIntLLROutputS6xD(220)(1);
  VNStageIntLLRInputS6xD(139)(3) <= CNStageIntLLROutputS6xD(220)(2);
  VNStageIntLLRInputS6xD(214)(3) <= CNStageIntLLROutputS6xD(220)(3);
  VNStageIntLLRInputS6xD(301)(3) <= CNStageIntLLROutputS6xD(220)(4);
  VNStageIntLLRInputS6xD(321)(3) <= CNStageIntLLROutputS6xD(220)(5);
  VNStageIntLLRInputS6xD(3)(2) <= CNStageIntLLROutputS6xD(221)(0);
  VNStageIntLLRInputS6xD(74)(3) <= CNStageIntLLROutputS6xD(221)(1);
  VNStageIntLLRInputS6xD(149)(3) <= CNStageIntLLROutputS6xD(221)(2);
  VNStageIntLLRInputS6xD(236)(3) <= CNStageIntLLROutputS6xD(221)(3);
  VNStageIntLLRInputS6xD(319)(3) <= CNStageIntLLROutputS6xD(221)(4);
  VNStageIntLLRInputS6xD(369)(2) <= CNStageIntLLROutputS6xD(221)(5);
  VNStageIntLLRInputS6xD(2)(3) <= CNStageIntLLROutputS6xD(222)(0);
  VNStageIntLLRInputS6xD(84)(3) <= CNStageIntLLROutputS6xD(222)(1);
  VNStageIntLLRInputS6xD(171)(2) <= CNStageIntLLROutputS6xD(222)(2);
  VNStageIntLLRInputS6xD(254)(1) <= CNStageIntLLROutputS6xD(222)(3);
  VNStageIntLLRInputS6xD(304)(3) <= CNStageIntLLROutputS6xD(222)(4);
  VNStageIntLLRInputS6xD(356)(3) <= CNStageIntLLROutputS6xD(222)(5);
  VNStageIntLLRInputS6xD(1)(2) <= CNStageIntLLROutputS6xD(223)(0);
  VNStageIntLLRInputS6xD(106)(2) <= CNStageIntLLROutputS6xD(223)(1);
  VNStageIntLLRInputS6xD(189)(2) <= CNStageIntLLROutputS6xD(223)(2);
  VNStageIntLLRInputS6xD(239)(3) <= CNStageIntLLROutputS6xD(223)(3);
  VNStageIntLLRInputS6xD(291)(3) <= CNStageIntLLROutputS6xD(223)(4);
  VNStageIntLLRInputS6xD(324)(3) <= CNStageIntLLROutputS6xD(223)(5);
  VNStageIntLLRInputS6xD(0)(3) <= CNStageIntLLROutputS6xD(224)(0);
  VNStageIntLLRInputS6xD(93)(3) <= CNStageIntLLROutputS6xD(224)(1);
  VNStageIntLLRInputS6xD(158)(3) <= CNStageIntLLROutputS6xD(224)(2);
  VNStageIntLLRInputS6xD(223)(3) <= CNStageIntLLROutputS6xD(224)(3);
  VNStageIntLLRInputS6xD(288)(3) <= CNStageIntLLROutputS6xD(224)(4);
  VNStageIntLLRInputS6xD(353)(3) <= CNStageIntLLROutputS6xD(224)(5);
  VNStageIntLLRInputS6xD(18)(4) <= CNStageIntLLROutputS6xD(225)(0);
  VNStageIntLLRInputS6xD(110)(4) <= CNStageIntLLROutputS6xD(225)(1);
  VNStageIntLLRInputS6xD(167)(4) <= CNStageIntLLROutputS6xD(225)(2);
  VNStageIntLLRInputS6xD(249)(2) <= CNStageIntLLROutputS6xD(225)(3);
  VNStageIntLLRInputS6xD(311)(3) <= CNStageIntLLROutputS6xD(225)(4);
  VNStageIntLLRInputS6xD(347)(4) <= CNStageIntLLROutputS6xD(225)(5);
  VNStageIntLLRInputS6xD(17)(4) <= CNStageIntLLROutputS6xD(226)(0);
  VNStageIntLLRInputS6xD(102)(4) <= CNStageIntLLROutputS6xD(226)(1);
  VNStageIntLLRInputS6xD(184)(4) <= CNStageIntLLROutputS6xD(226)(2);
  VNStageIntLLRInputS6xD(246)(4) <= CNStageIntLLROutputS6xD(226)(3);
  VNStageIntLLRInputS6xD(282)(4) <= CNStageIntLLROutputS6xD(226)(4);
  VNStageIntLLRInputS6xD(367)(4) <= CNStageIntLLROutputS6xD(226)(5);
  VNStageIntLLRInputS6xD(16)(3) <= CNStageIntLLROutputS6xD(227)(0);
  VNStageIntLLRInputS6xD(119)(3) <= CNStageIntLLROutputS6xD(227)(1);
  VNStageIntLLRInputS6xD(181)(4) <= CNStageIntLLROutputS6xD(227)(2);
  VNStageIntLLRInputS6xD(217)(4) <= CNStageIntLLROutputS6xD(227)(3);
  VNStageIntLLRInputS6xD(302)(4) <= CNStageIntLLROutputS6xD(227)(4);
  VNStageIntLLRInputS6xD(353)(4) <= CNStageIntLLROutputS6xD(227)(5);
  VNStageIntLLRInputS6xD(15)(4) <= CNStageIntLLROutputS6xD(228)(0);
  VNStageIntLLRInputS6xD(116)(3) <= CNStageIntLLROutputS6xD(228)(1);
  VNStageIntLLRInputS6xD(152)(4) <= CNStageIntLLROutputS6xD(228)(2);
  VNStageIntLLRInputS6xD(237)(3) <= CNStageIntLLROutputS6xD(228)(3);
  VNStageIntLLRInputS6xD(288)(4) <= CNStageIntLLROutputS6xD(228)(4);
  VNStageIntLLRInputS6xD(343)(4) <= CNStageIntLLROutputS6xD(228)(5);
  VNStageIntLLRInputS6xD(14)(4) <= CNStageIntLLROutputS6xD(229)(0);
  VNStageIntLLRInputS6xD(87)(4) <= CNStageIntLLROutputS6xD(229)(1);
  VNStageIntLLRInputS6xD(172)(3) <= CNStageIntLLROutputS6xD(229)(2);
  VNStageIntLLRInputS6xD(223)(4) <= CNStageIntLLROutputS6xD(229)(3);
  VNStageIntLLRInputS6xD(278)(3) <= CNStageIntLLROutputS6xD(229)(4);
  VNStageIntLLRInputS6xD(372)(3) <= CNStageIntLLROutputS6xD(229)(5);
  VNStageIntLLRInputS6xD(13)(3) <= CNStageIntLLROutputS6xD(230)(0);
  VNStageIntLLRInputS6xD(107)(3) <= CNStageIntLLROutputS6xD(230)(1);
  VNStageIntLLRInputS6xD(158)(4) <= CNStageIntLLROutputS6xD(230)(2);
  VNStageIntLLRInputS6xD(213)(3) <= CNStageIntLLROutputS6xD(230)(3);
  VNStageIntLLRInputS6xD(307)(4) <= CNStageIntLLROutputS6xD(230)(4);
  VNStageIntLLRInputS6xD(355)(4) <= CNStageIntLLROutputS6xD(230)(5);
  VNStageIntLLRInputS6xD(12)(4) <= CNStageIntLLROutputS6xD(231)(0);
  VNStageIntLLRInputS6xD(93)(4) <= CNStageIntLLROutputS6xD(231)(1);
  VNStageIntLLRInputS6xD(148)(4) <= CNStageIntLLROutputS6xD(231)(2);
  VNStageIntLLRInputS6xD(242)(4) <= CNStageIntLLROutputS6xD(231)(3);
  VNStageIntLLRInputS6xD(290)(4) <= CNStageIntLLROutputS6xD(231)(4);
  VNStageIntLLRInputS6xD(322)(3) <= CNStageIntLLROutputS6xD(231)(5);
  VNStageIntLLRInputS6xD(11)(4) <= CNStageIntLLROutputS6xD(232)(0);
  VNStageIntLLRInputS6xD(83)(4) <= CNStageIntLLROutputS6xD(232)(1);
  VNStageIntLLRInputS6xD(177)(4) <= CNStageIntLLROutputS6xD(232)(2);
  VNStageIntLLRInputS6xD(225)(4) <= CNStageIntLLROutputS6xD(232)(3);
  VNStageIntLLRInputS6xD(257)(4) <= CNStageIntLLROutputS6xD(232)(4);
  VNStageIntLLRInputS6xD(345)(3) <= CNStageIntLLROutputS6xD(232)(5);
  VNStageIntLLRInputS6xD(10)(3) <= CNStageIntLLROutputS6xD(233)(0);
  VNStageIntLLRInputS6xD(112)(4) <= CNStageIntLLROutputS6xD(233)(1);
  VNStageIntLLRInputS6xD(160)(4) <= CNStageIntLLROutputS6xD(233)(2);
  VNStageIntLLRInputS6xD(255)(4) <= CNStageIntLLROutputS6xD(233)(3);
  VNStageIntLLRInputS6xD(280)(4) <= CNStageIntLLROutputS6xD(233)(4);
  VNStageIntLLRInputS6xD(381)(3) <= CNStageIntLLROutputS6xD(233)(5);
  VNStageIntLLRInputS6xD(9)(4) <= CNStageIntLLROutputS6xD(234)(0);
  VNStageIntLLRInputS6xD(95)(4) <= CNStageIntLLROutputS6xD(234)(1);
  VNStageIntLLRInputS6xD(190)(2) <= CNStageIntLLROutputS6xD(234)(2);
  VNStageIntLLRInputS6xD(215)(4) <= CNStageIntLLROutputS6xD(234)(3);
  VNStageIntLLRInputS6xD(316)(2) <= CNStageIntLLROutputS6xD(234)(4);
  VNStageIntLLRInputS6xD(365)(4) <= CNStageIntLLROutputS6xD(234)(5);
  VNStageIntLLRInputS6xD(7)(4) <= CNStageIntLLROutputS6xD(235)(0);
  VNStageIntLLRInputS6xD(85)(3) <= CNStageIntLLROutputS6xD(235)(1);
  VNStageIntLLRInputS6xD(186)(3) <= CNStageIntLLROutputS6xD(235)(2);
  VNStageIntLLRInputS6xD(235)(3) <= CNStageIntLLROutputS6xD(235)(3);
  VNStageIntLLRInputS6xD(303)(4) <= CNStageIntLLROutputS6xD(235)(4);
  VNStageIntLLRInputS6xD(346)(4) <= CNStageIntLLROutputS6xD(235)(5);
  VNStageIntLLRInputS6xD(6)(4) <= CNStageIntLLROutputS6xD(236)(0);
  VNStageIntLLRInputS6xD(121)(3) <= CNStageIntLLROutputS6xD(236)(1);
  VNStageIntLLRInputS6xD(170)(3) <= CNStageIntLLROutputS6xD(236)(2);
  VNStageIntLLRInputS6xD(238)(4) <= CNStageIntLLROutputS6xD(236)(3);
  VNStageIntLLRInputS6xD(281)(4) <= CNStageIntLLROutputS6xD(236)(4);
  VNStageIntLLRInputS6xD(321)(4) <= CNStageIntLLROutputS6xD(236)(5);
  VNStageIntLLRInputS6xD(5)(4) <= CNStageIntLLROutputS6xD(237)(0);
  VNStageIntLLRInputS6xD(105)(3) <= CNStageIntLLROutputS6xD(237)(1);
  VNStageIntLLRInputS6xD(173)(4) <= CNStageIntLLROutputS6xD(237)(2);
  VNStageIntLLRInputS6xD(216)(4) <= CNStageIntLLROutputS6xD(237)(3);
  VNStageIntLLRInputS6xD(319)(4) <= CNStageIntLLROutputS6xD(237)(4);
  VNStageIntLLRInputS6xD(382)(3) <= CNStageIntLLROutputS6xD(237)(5);
  VNStageIntLLRInputS6xD(4)(3) <= CNStageIntLLROutputS6xD(238)(0);
  VNStageIntLLRInputS6xD(108)(4) <= CNStageIntLLROutputS6xD(238)(1);
  VNStageIntLLRInputS6xD(151)(4) <= CNStageIntLLROutputS6xD(238)(2);
  VNStageIntLLRInputS6xD(254)(2) <= CNStageIntLLROutputS6xD(238)(3);
  VNStageIntLLRInputS6xD(317)(1) <= CNStageIntLLROutputS6xD(238)(4);
  VNStageIntLLRInputS6xD(344)(4) <= CNStageIntLLROutputS6xD(238)(5);
  VNStageIntLLRInputS6xD(3)(3) <= CNStageIntLLROutputS6xD(239)(0);
  VNStageIntLLRInputS6xD(86)(2) <= CNStageIntLLROutputS6xD(239)(1);
  VNStageIntLLRInputS6xD(189)(3) <= CNStageIntLLROutputS6xD(239)(2);
  VNStageIntLLRInputS6xD(252)(3) <= CNStageIntLLROutputS6xD(239)(3);
  VNStageIntLLRInputS6xD(279)(4) <= CNStageIntLLROutputS6xD(239)(4);
  VNStageIntLLRInputS6xD(352)(4) <= CNStageIntLLROutputS6xD(239)(5);
  VNStageIntLLRInputS6xD(2)(4) <= CNStageIntLLROutputS6xD(240)(0);
  VNStageIntLLRInputS6xD(124)(2) <= CNStageIntLLROutputS6xD(240)(1);
  VNStageIntLLRInputS6xD(187)(3) <= CNStageIntLLROutputS6xD(240)(2);
  VNStageIntLLRInputS6xD(214)(4) <= CNStageIntLLROutputS6xD(240)(3);
  VNStageIntLLRInputS6xD(287)(4) <= CNStageIntLLROutputS6xD(240)(4);
  VNStageIntLLRInputS6xD(332)(4) <= CNStageIntLLROutputS6xD(240)(5);
  VNStageIntLLRInputS6xD(1)(3) <= CNStageIntLLROutputS6xD(241)(0);
  VNStageIntLLRInputS6xD(122)(3) <= CNStageIntLLROutputS6xD(241)(1);
  VNStageIntLLRInputS6xD(149)(4) <= CNStageIntLLROutputS6xD(241)(2);
  VNStageIntLLRInputS6xD(222)(2) <= CNStageIntLLROutputS6xD(241)(3);
  VNStageIntLLRInputS6xD(267)(4) <= CNStageIntLLROutputS6xD(241)(4);
  VNStageIntLLRInputS6xD(326)(3) <= CNStageIntLLROutputS6xD(241)(5);
  VNStageIntLLRInputS6xD(62)(3) <= CNStageIntLLROutputS6xD(242)(0);
  VNStageIntLLRInputS6xD(92)(4) <= CNStageIntLLROutputS6xD(242)(1);
  VNStageIntLLRInputS6xD(137)(4) <= CNStageIntLLROutputS6xD(242)(2);
  VNStageIntLLRInputS6xD(196)(4) <= CNStageIntLLROutputS6xD(242)(3);
  VNStageIntLLRInputS6xD(256)(3) <= CNStageIntLLROutputS6xD(242)(4);
  VNStageIntLLRInputS6xD(325)(4) <= CNStageIntLLROutputS6xD(242)(5);
  VNStageIntLLRInputS6xD(61)(3) <= CNStageIntLLROutputS6xD(243)(0);
  VNStageIntLLRInputS6xD(72)(4) <= CNStageIntLLROutputS6xD(243)(1);
  VNStageIntLLRInputS6xD(131)(3) <= CNStageIntLLROutputS6xD(243)(2);
  VNStageIntLLRInputS6xD(192)(4) <= CNStageIntLLROutputS6xD(243)(3);
  VNStageIntLLRInputS6xD(260)(4) <= CNStageIntLLROutputS6xD(243)(4);
  VNStageIntLLRInputS6xD(330)(4) <= CNStageIntLLROutputS6xD(243)(5);
  VNStageIntLLRInputS6xD(60)(3) <= CNStageIntLLROutputS6xD(244)(0);
  VNStageIntLLRInputS6xD(66)(3) <= CNStageIntLLROutputS6xD(244)(1);
  VNStageIntLLRInputS6xD(128)(4) <= CNStageIntLLROutputS6xD(244)(2);
  VNStageIntLLRInputS6xD(195)(3) <= CNStageIntLLROutputS6xD(244)(3);
  VNStageIntLLRInputS6xD(265)(3) <= CNStageIntLLROutputS6xD(244)(4);
  VNStageIntLLRInputS6xD(349)(3) <= CNStageIntLLROutputS6xD(244)(5);
  VNStageIntLLRInputS6xD(59)(2) <= CNStageIntLLROutputS6xD(245)(0);
  VNStageIntLLRInputS6xD(64)(3) <= CNStageIntLLROutputS6xD(245)(1);
  VNStageIntLLRInputS6xD(130)(4) <= CNStageIntLLROutputS6xD(245)(2);
  VNStageIntLLRInputS6xD(200)(4) <= CNStageIntLLROutputS6xD(245)(3);
  VNStageIntLLRInputS6xD(284)(4) <= CNStageIntLLROutputS6xD(245)(4);
  VNStageIntLLRInputS6xD(340)(4) <= CNStageIntLLROutputS6xD(245)(5);
  VNStageIntLLRInputS6xD(57)(3) <= CNStageIntLLROutputS6xD(246)(0);
  VNStageIntLLRInputS6xD(70)(4) <= CNStageIntLLROutputS6xD(246)(1);
  VNStageIntLLRInputS6xD(154)(3) <= CNStageIntLLROutputS6xD(246)(2);
  VNStageIntLLRInputS6xD(210)(4) <= CNStageIntLLROutputS6xD(246)(3);
  VNStageIntLLRInputS6xD(312)(3) <= CNStageIntLLROutputS6xD(246)(4);
  VNStageIntLLRInputS6xD(378)(3) <= CNStageIntLLROutputS6xD(246)(5);
  VNStageIntLLRInputS6xD(56)(4) <= CNStageIntLLROutputS6xD(247)(0);
  VNStageIntLLRInputS6xD(89)(4) <= CNStageIntLLROutputS6xD(247)(1);
  VNStageIntLLRInputS6xD(145)(4) <= CNStageIntLLROutputS6xD(247)(2);
  VNStageIntLLRInputS6xD(247)(4) <= CNStageIntLLROutputS6xD(247)(3);
  VNStageIntLLRInputS6xD(313)(2) <= CNStageIntLLROutputS6xD(247)(4);
  VNStageIntLLRInputS6xD(339)(4) <= CNStageIntLLROutputS6xD(247)(5);
  VNStageIntLLRInputS6xD(55)(4) <= CNStageIntLLROutputS6xD(248)(0);
  VNStageIntLLRInputS6xD(80)(4) <= CNStageIntLLROutputS6xD(248)(1);
  VNStageIntLLRInputS6xD(182)(4) <= CNStageIntLLROutputS6xD(248)(2);
  VNStageIntLLRInputS6xD(248)(4) <= CNStageIntLLROutputS6xD(248)(3);
  VNStageIntLLRInputS6xD(274)(3) <= CNStageIntLLROutputS6xD(248)(4);
  VNStageIntLLRInputS6xD(360)(4) <= CNStageIntLLROutputS6xD(248)(5);
  VNStageIntLLRInputS6xD(53)(3) <= CNStageIntLLROutputS6xD(249)(0);
  VNStageIntLLRInputS6xD(118)(3) <= CNStageIntLLROutputS6xD(249)(1);
  VNStageIntLLRInputS6xD(144)(4) <= CNStageIntLLROutputS6xD(249)(2);
  VNStageIntLLRInputS6xD(230)(3) <= CNStageIntLLROutputS6xD(249)(3);
  VNStageIntLLRInputS6xD(291)(4) <= CNStageIntLLROutputS6xD(249)(4);
  VNStageIntLLRInputS6xD(371)(3) <= CNStageIntLLROutputS6xD(249)(5);
  VNStageIntLLRInputS6xD(51)(3) <= CNStageIntLLROutputS6xD(250)(0);
  VNStageIntLLRInputS6xD(100)(4) <= CNStageIntLLROutputS6xD(250)(1);
  VNStageIntLLRInputS6xD(161)(4) <= CNStageIntLLROutputS6xD(250)(2);
  VNStageIntLLRInputS6xD(241)(3) <= CNStageIntLLROutputS6xD(250)(3);
  VNStageIntLLRInputS6xD(269)(3) <= CNStageIntLLROutputS6xD(250)(4);
  VNStageIntLLRInputS6xD(373)(2) <= CNStageIntLLROutputS6xD(250)(5);
  VNStageIntLLRInputS6xD(50)(4) <= CNStageIntLLROutputS6xD(251)(0);
  VNStageIntLLRInputS6xD(96)(4) <= CNStageIntLLROutputS6xD(251)(1);
  VNStageIntLLRInputS6xD(176)(4) <= CNStageIntLLROutputS6xD(251)(2);
  VNStageIntLLRInputS6xD(204)(4) <= CNStageIntLLROutputS6xD(251)(3);
  VNStageIntLLRInputS6xD(308)(2) <= CNStageIntLLROutputS6xD(251)(4);
  VNStageIntLLRInputS6xD(342)(3) <= CNStageIntLLROutputS6xD(251)(5);
  VNStageIntLLRInputS6xD(49)(4) <= CNStageIntLLROutputS6xD(252)(0);
  VNStageIntLLRInputS6xD(111)(4) <= CNStageIntLLROutputS6xD(252)(1);
  VNStageIntLLRInputS6xD(139)(4) <= CNStageIntLLROutputS6xD(252)(2);
  VNStageIntLLRInputS6xD(243)(4) <= CNStageIntLLROutputS6xD(252)(3);
  VNStageIntLLRInputS6xD(277)(4) <= CNStageIntLLROutputS6xD(252)(4);
  VNStageIntLLRInputS6xD(358)(3) <= CNStageIntLLROutputS6xD(252)(5);
  VNStageIntLLRInputS6xD(47)(2) <= CNStageIntLLROutputS6xD(253)(0);
  VNStageIntLLRInputS6xD(113)(4) <= CNStageIntLLROutputS6xD(253)(1);
  VNStageIntLLRInputS6xD(147)(4) <= CNStageIntLLROutputS6xD(253)(2);
  VNStageIntLLRInputS6xD(228)(4) <= CNStageIntLLROutputS6xD(253)(3);
  VNStageIntLLRInputS6xD(263)(4) <= CNStageIntLLROutputS6xD(253)(4);
  VNStageIntLLRInputS6xD(337)(4) <= CNStageIntLLROutputS6xD(253)(5);
  VNStageIntLLRInputS6xD(46)(4) <= CNStageIntLLROutputS6xD(254)(0);
  VNStageIntLLRInputS6xD(82)(4) <= CNStageIntLLROutputS6xD(254)(1);
  VNStageIntLLRInputS6xD(163)(3) <= CNStageIntLLROutputS6xD(254)(2);
  VNStageIntLLRInputS6xD(198)(4) <= CNStageIntLLROutputS6xD(254)(3);
  VNStageIntLLRInputS6xD(272)(4) <= CNStageIntLLROutputS6xD(254)(4);
  VNStageIntLLRInputS6xD(350)(4) <= CNStageIntLLROutputS6xD(254)(5);
  VNStageIntLLRInputS6xD(45)(4) <= CNStageIntLLROutputS6xD(255)(0);
  VNStageIntLLRInputS6xD(98)(3) <= CNStageIntLLROutputS6xD(255)(1);
  VNStageIntLLRInputS6xD(133)(2) <= CNStageIntLLROutputS6xD(255)(2);
  VNStageIntLLRInputS6xD(207)(3) <= CNStageIntLLROutputS6xD(255)(3);
  VNStageIntLLRInputS6xD(285)(4) <= CNStageIntLLROutputS6xD(255)(4);
  VNStageIntLLRInputS6xD(329)(4) <= CNStageIntLLROutputS6xD(255)(5);
  VNStageIntLLRInputS6xD(44)(4) <= CNStageIntLLROutputS6xD(256)(0);
  VNStageIntLLRInputS6xD(68)(3) <= CNStageIntLLROutputS6xD(256)(1);
  VNStageIntLLRInputS6xD(142)(3) <= CNStageIntLLROutputS6xD(256)(2);
  VNStageIntLLRInputS6xD(220)(4) <= CNStageIntLLROutputS6xD(256)(3);
  VNStageIntLLRInputS6xD(264)(4) <= CNStageIntLLROutputS6xD(256)(4);
  VNStageIntLLRInputS6xD(357)(4) <= CNStageIntLLROutputS6xD(256)(5);
  VNStageIntLLRInputS6xD(43)(3) <= CNStageIntLLROutputS6xD(257)(0);
  VNStageIntLLRInputS6xD(77)(2) <= CNStageIntLLROutputS6xD(257)(1);
  VNStageIntLLRInputS6xD(155)(4) <= CNStageIntLLROutputS6xD(257)(2);
  VNStageIntLLRInputS6xD(199)(4) <= CNStageIntLLROutputS6xD(257)(3);
  VNStageIntLLRInputS6xD(292)(4) <= CNStageIntLLROutputS6xD(257)(4);
  VNStageIntLLRInputS6xD(359)(4) <= CNStageIntLLROutputS6xD(257)(5);
  VNStageIntLLRInputS6xD(42)(4) <= CNStageIntLLROutputS6xD(258)(0);
  VNStageIntLLRInputS6xD(90)(4) <= CNStageIntLLROutputS6xD(258)(1);
  VNStageIntLLRInputS6xD(134)(3) <= CNStageIntLLROutputS6xD(258)(2);
  VNStageIntLLRInputS6xD(227)(4) <= CNStageIntLLROutputS6xD(258)(3);
  VNStageIntLLRInputS6xD(294)(4) <= CNStageIntLLROutputS6xD(258)(4);
  VNStageIntLLRInputS6xD(341)(4) <= CNStageIntLLROutputS6xD(258)(5);
  VNStageIntLLRInputS6xD(41)(4) <= CNStageIntLLROutputS6xD(259)(0);
  VNStageIntLLRInputS6xD(69)(4) <= CNStageIntLLROutputS6xD(259)(1);
  VNStageIntLLRInputS6xD(162)(4) <= CNStageIntLLROutputS6xD(259)(2);
  VNStageIntLLRInputS6xD(229)(3) <= CNStageIntLLROutputS6xD(259)(3);
  VNStageIntLLRInputS6xD(276)(4) <= CNStageIntLLROutputS6xD(259)(4);
  VNStageIntLLRInputS6xD(348)(4) <= CNStageIntLLROutputS6xD(259)(5);
  VNStageIntLLRInputS6xD(40)(3) <= CNStageIntLLROutputS6xD(260)(0);
  VNStageIntLLRInputS6xD(97)(4) <= CNStageIntLLROutputS6xD(260)(1);
  VNStageIntLLRInputS6xD(164)(4) <= CNStageIntLLROutputS6xD(260)(2);
  VNStageIntLLRInputS6xD(211)(4) <= CNStageIntLLROutputS6xD(260)(3);
  VNStageIntLLRInputS6xD(283)(4) <= CNStageIntLLROutputS6xD(260)(4);
  VNStageIntLLRInputS6xD(375)(3) <= CNStageIntLLROutputS6xD(260)(5);
  VNStageIntLLRInputS6xD(39)(4) <= CNStageIntLLROutputS6xD(261)(0);
  VNStageIntLLRInputS6xD(99)(4) <= CNStageIntLLROutputS6xD(261)(1);
  VNStageIntLLRInputS6xD(146)(3) <= CNStageIntLLROutputS6xD(261)(2);
  VNStageIntLLRInputS6xD(218)(4) <= CNStageIntLLROutputS6xD(261)(3);
  VNStageIntLLRInputS6xD(310)(3) <= CNStageIntLLROutputS6xD(261)(4);
  VNStageIntLLRInputS6xD(363)(3) <= CNStageIntLLROutputS6xD(261)(5);
  VNStageIntLLRInputS6xD(38)(4) <= CNStageIntLLROutputS6xD(262)(0);
  VNStageIntLLRInputS6xD(81)(3) <= CNStageIntLLROutputS6xD(262)(1);
  VNStageIntLLRInputS6xD(153)(4) <= CNStageIntLLROutputS6xD(262)(2);
  VNStageIntLLRInputS6xD(245)(4) <= CNStageIntLLROutputS6xD(262)(3);
  VNStageIntLLRInputS6xD(298)(4) <= CNStageIntLLROutputS6xD(262)(4);
  VNStageIntLLRInputS6xD(369)(3) <= CNStageIntLLROutputS6xD(262)(5);
  VNStageIntLLRInputS6xD(37)(4) <= CNStageIntLLROutputS6xD(263)(0);
  VNStageIntLLRInputS6xD(88)(4) <= CNStageIntLLROutputS6xD(263)(1);
  VNStageIntLLRInputS6xD(180)(2) <= CNStageIntLLROutputS6xD(263)(2);
  VNStageIntLLRInputS6xD(233)(3) <= CNStageIntLLROutputS6xD(263)(3);
  VNStageIntLLRInputS6xD(304)(4) <= CNStageIntLLROutputS6xD(263)(4);
  VNStageIntLLRInputS6xD(364)(4) <= CNStageIntLLROutputS6xD(263)(5);
  VNStageIntLLRInputS6xD(36)(3) <= CNStageIntLLROutputS6xD(264)(0);
  VNStageIntLLRInputS6xD(115)(4) <= CNStageIntLLROutputS6xD(264)(1);
  VNStageIntLLRInputS6xD(168)(3) <= CNStageIntLLROutputS6xD(264)(2);
  VNStageIntLLRInputS6xD(239)(4) <= CNStageIntLLROutputS6xD(264)(3);
  VNStageIntLLRInputS6xD(299)(3) <= CNStageIntLLROutputS6xD(264)(4);
  VNStageIntLLRInputS6xD(374)(4) <= CNStageIntLLROutputS6xD(264)(5);
  VNStageIntLLRInputS6xD(35)(4) <= CNStageIntLLROutputS6xD(265)(0);
  VNStageIntLLRInputS6xD(103)(4) <= CNStageIntLLROutputS6xD(265)(1);
  VNStageIntLLRInputS6xD(174)(3) <= CNStageIntLLROutputS6xD(265)(2);
  VNStageIntLLRInputS6xD(234)(4) <= CNStageIntLLROutputS6xD(265)(3);
  VNStageIntLLRInputS6xD(309)(4) <= CNStageIntLLROutputS6xD(265)(4);
  VNStageIntLLRInputS6xD(333)(3) <= CNStageIntLLROutputS6xD(265)(5);
  VNStageIntLLRInputS6xD(34)(4) <= CNStageIntLLROutputS6xD(266)(0);
  VNStageIntLLRInputS6xD(109)(4) <= CNStageIntLLROutputS6xD(266)(1);
  VNStageIntLLRInputS6xD(169)(4) <= CNStageIntLLROutputS6xD(266)(2);
  VNStageIntLLRInputS6xD(244)(1) <= CNStageIntLLROutputS6xD(266)(3);
  VNStageIntLLRInputS6xD(268)(4) <= CNStageIntLLROutputS6xD(266)(4);
  VNStageIntLLRInputS6xD(351)(3) <= CNStageIntLLROutputS6xD(266)(5);
  VNStageIntLLRInputS6xD(33)(4) <= CNStageIntLLROutputS6xD(267)(0);
  VNStageIntLLRInputS6xD(104)(4) <= CNStageIntLLROutputS6xD(267)(1);
  VNStageIntLLRInputS6xD(179)(4) <= CNStageIntLLROutputS6xD(267)(2);
  VNStageIntLLRInputS6xD(203)(4) <= CNStageIntLLROutputS6xD(267)(3);
  VNStageIntLLRInputS6xD(286)(4) <= CNStageIntLLROutputS6xD(267)(4);
  VNStageIntLLRInputS6xD(336)(3) <= CNStageIntLLROutputS6xD(267)(5);
  VNStageIntLLRInputS6xD(32)(3) <= CNStageIntLLROutputS6xD(268)(0);
  VNStageIntLLRInputS6xD(114)(4) <= CNStageIntLLROutputS6xD(268)(1);
  VNStageIntLLRInputS6xD(138)(4) <= CNStageIntLLROutputS6xD(268)(2);
  VNStageIntLLRInputS6xD(221)(4) <= CNStageIntLLROutputS6xD(268)(3);
  VNStageIntLLRInputS6xD(271)(3) <= CNStageIntLLROutputS6xD(268)(4);
  VNStageIntLLRInputS6xD(323)(3) <= CNStageIntLLROutputS6xD(268)(5);
  VNStageIntLLRInputS6xD(30)(4) <= CNStageIntLLROutputS6xD(269)(0);
  VNStageIntLLRInputS6xD(91)(4) <= CNStageIntLLROutputS6xD(269)(1);
  VNStageIntLLRInputS6xD(141)(2) <= CNStageIntLLROutputS6xD(269)(2);
  VNStageIntLLRInputS6xD(193)(3) <= CNStageIntLLROutputS6xD(269)(3);
  VNStageIntLLRInputS6xD(289)(4) <= CNStageIntLLROutputS6xD(269)(4);
  VNStageIntLLRInputS6xD(366)(4) <= CNStageIntLLROutputS6xD(269)(5);
  VNStageIntLLRInputS6xD(29)(3) <= CNStageIntLLROutputS6xD(270)(0);
  VNStageIntLLRInputS6xD(76)(4) <= CNStageIntLLROutputS6xD(270)(1);
  VNStageIntLLRInputS6xD(191)(4) <= CNStageIntLLROutputS6xD(270)(2);
  VNStageIntLLRInputS6xD(224)(4) <= CNStageIntLLROutputS6xD(270)(3);
  VNStageIntLLRInputS6xD(301)(4) <= CNStageIntLLROutputS6xD(270)(4);
  VNStageIntLLRInputS6xD(380)(3) <= CNStageIntLLROutputS6xD(270)(5);
  VNStageIntLLRInputS6xD(28)(4) <= CNStageIntLLROutputS6xD(271)(0);
  VNStageIntLLRInputS6xD(126)(3) <= CNStageIntLLROutputS6xD(271)(1);
  VNStageIntLLRInputS6xD(159)(3) <= CNStageIntLLROutputS6xD(271)(2);
  VNStageIntLLRInputS6xD(236)(4) <= CNStageIntLLROutputS6xD(271)(3);
  VNStageIntLLRInputS6xD(315)(3) <= CNStageIntLLROutputS6xD(271)(4);
  VNStageIntLLRInputS6xD(361)(4) <= CNStageIntLLROutputS6xD(271)(5);
  VNStageIntLLRInputS6xD(26)(4) <= CNStageIntLLROutputS6xD(272)(0);
  VNStageIntLLRInputS6xD(106)(3) <= CNStageIntLLROutputS6xD(272)(1);
  VNStageIntLLRInputS6xD(185)(1) <= CNStageIntLLROutputS6xD(272)(2);
  VNStageIntLLRInputS6xD(231)(3) <= CNStageIntLLROutputS6xD(272)(3);
  VNStageIntLLRInputS6xD(273)(3) <= CNStageIntLLROutputS6xD(272)(4);
  VNStageIntLLRInputS6xD(327)(4) <= CNStageIntLLROutputS6xD(272)(5);
  VNStageIntLLRInputS6xD(24)(4) <= CNStageIntLLROutputS6xD(273)(0);
  VNStageIntLLRInputS6xD(101)(4) <= CNStageIntLLROutputS6xD(273)(1);
  VNStageIntLLRInputS6xD(143)(4) <= CNStageIntLLROutputS6xD(273)(2);
  VNStageIntLLRInputS6xD(197)(4) <= CNStageIntLLROutputS6xD(273)(3);
  VNStageIntLLRInputS6xD(266)(3) <= CNStageIntLLROutputS6xD(273)(4);
  VNStageIntLLRInputS6xD(324)(4) <= CNStageIntLLROutputS6xD(273)(5);
  VNStageIntLLRInputS6xD(23)(4) <= CNStageIntLLROutputS6xD(274)(0);
  VNStageIntLLRInputS6xD(78)(4) <= CNStageIntLLROutputS6xD(274)(1);
  VNStageIntLLRInputS6xD(132)(3) <= CNStageIntLLROutputS6xD(274)(2);
  VNStageIntLLRInputS6xD(201)(4) <= CNStageIntLLROutputS6xD(274)(3);
  VNStageIntLLRInputS6xD(259)(2) <= CNStageIntLLROutputS6xD(274)(4);
  VNStageIntLLRInputS6xD(335)(4) <= CNStageIntLLROutputS6xD(274)(5);
  VNStageIntLLRInputS6xD(22)(4) <= CNStageIntLLROutputS6xD(275)(0);
  VNStageIntLLRInputS6xD(67)(1) <= CNStageIntLLROutputS6xD(275)(1);
  VNStageIntLLRInputS6xD(136)(4) <= CNStageIntLLROutputS6xD(275)(2);
  VNStageIntLLRInputS6xD(194)(4) <= CNStageIntLLROutputS6xD(275)(3);
  VNStageIntLLRInputS6xD(270)(4) <= CNStageIntLLROutputS6xD(275)(4);
  VNStageIntLLRInputS6xD(370)(3) <= CNStageIntLLROutputS6xD(275)(5);
  VNStageIntLLRInputS6xD(21)(4) <= CNStageIntLLROutputS6xD(276)(0);
  VNStageIntLLRInputS6xD(71)(3) <= CNStageIntLLROutputS6xD(276)(1);
  VNStageIntLLRInputS6xD(129)(4) <= CNStageIntLLROutputS6xD(276)(2);
  VNStageIntLLRInputS6xD(205)(1) <= CNStageIntLLROutputS6xD(276)(3);
  VNStageIntLLRInputS6xD(305)(4) <= CNStageIntLLROutputS6xD(276)(4);
  VNStageIntLLRInputS6xD(362)(4) <= CNStageIntLLROutputS6xD(276)(5);
  VNStageIntLLRInputS6xD(20)(2) <= CNStageIntLLROutputS6xD(277)(0);
  VNStageIntLLRInputS6xD(127)(4) <= CNStageIntLLROutputS6xD(277)(1);
  VNStageIntLLRInputS6xD(140)(4) <= CNStageIntLLROutputS6xD(277)(2);
  VNStageIntLLRInputS6xD(240)(4) <= CNStageIntLLROutputS6xD(277)(3);
  VNStageIntLLRInputS6xD(297)(4) <= CNStageIntLLROutputS6xD(277)(4);
  VNStageIntLLRInputS6xD(379)(2) <= CNStageIntLLROutputS6xD(277)(5);
  VNStageIntLLRInputS6xD(19)(3) <= CNStageIntLLROutputS6xD(278)(0);
  VNStageIntLLRInputS6xD(75)(4) <= CNStageIntLLROutputS6xD(278)(1);
  VNStageIntLLRInputS6xD(175)(4) <= CNStageIntLLROutputS6xD(278)(2);
  VNStageIntLLRInputS6xD(232)(3) <= CNStageIntLLROutputS6xD(278)(3);
  VNStageIntLLRInputS6xD(314)(1) <= CNStageIntLLROutputS6xD(278)(4);
  VNStageIntLLRInputS6xD(376)(3) <= CNStageIntLLROutputS6xD(278)(5);
  VNStageIntLLRInputS6xD(0)(4) <= CNStageIntLLROutputS6xD(279)(0);
  VNStageIntLLRInputS6xD(123)(3) <= CNStageIntLLROutputS6xD(279)(1);
  VNStageIntLLRInputS6xD(188)(2) <= CNStageIntLLROutputS6xD(279)(2);
  VNStageIntLLRInputS6xD(253)(3) <= CNStageIntLLROutputS6xD(279)(3);
  VNStageIntLLRInputS6xD(318)(2) <= CNStageIntLLROutputS6xD(279)(4);
  VNStageIntLLRInputS6xD(383)(4) <= CNStageIntLLROutputS6xD(279)(5);
  VNStageIntLLRInputS6xD(35)(5) <= CNStageIntLLROutputS6xD(280)(0);
  VNStageIntLLRInputS6xD(91)(5) <= CNStageIntLLROutputS6xD(280)(1);
  VNStageIntLLRInputS6xD(191)(5) <= CNStageIntLLROutputS6xD(280)(2);
  VNStageIntLLRInputS6xD(248)(5) <= CNStageIntLLROutputS6xD(280)(3);
  VNStageIntLLRInputS6xD(267)(5) <= CNStageIntLLROutputS6xD(280)(4);
  VNStageIntLLRInputS6xD(329)(5) <= CNStageIntLLROutputS6xD(280)(5);
  VNStageIntLLRInputS6xD(34)(5) <= CNStageIntLLROutputS6xD(281)(0);
  VNStageIntLLRInputS6xD(126)(4) <= CNStageIntLLROutputS6xD(281)(1);
  VNStageIntLLRInputS6xD(183)(3) <= CNStageIntLLROutputS6xD(281)(2);
  VNStageIntLLRInputS6xD(202)(4) <= CNStageIntLLROutputS6xD(281)(3);
  VNStageIntLLRInputS6xD(264)(5) <= CNStageIntLLROutputS6xD(281)(4);
  VNStageIntLLRInputS6xD(363)(4) <= CNStageIntLLROutputS6xD(281)(5);
  VNStageIntLLRInputS6xD(33)(5) <= CNStageIntLLROutputS6xD(282)(0);
  VNStageIntLLRInputS6xD(118)(4) <= CNStageIntLLROutputS6xD(282)(1);
  VNStageIntLLRInputS6xD(137)(5) <= CNStageIntLLROutputS6xD(282)(2);
  VNStageIntLLRInputS6xD(199)(5) <= CNStageIntLLROutputS6xD(282)(3);
  VNStageIntLLRInputS6xD(298)(5) <= CNStageIntLLROutputS6xD(282)(4);
  VNStageIntLLRInputS6xD(383)(5) <= CNStageIntLLROutputS6xD(282)(5);
  VNStageIntLLRInputS6xD(31)(3) <= CNStageIntLLROutputS6xD(283)(0);
  VNStageIntLLRInputS6xD(69)(5) <= CNStageIntLLROutputS6xD(283)(1);
  VNStageIntLLRInputS6xD(168)(4) <= CNStageIntLLROutputS6xD(283)(2);
  VNStageIntLLRInputS6xD(253)(4) <= CNStageIntLLROutputS6xD(283)(3);
  VNStageIntLLRInputS6xD(304)(5) <= CNStageIntLLROutputS6xD(283)(4);
  VNStageIntLLRInputS6xD(359)(5) <= CNStageIntLLROutputS6xD(283)(5);
  VNStageIntLLRInputS6xD(30)(5) <= CNStageIntLLROutputS6xD(284)(0);
  VNStageIntLLRInputS6xD(103)(5) <= CNStageIntLLROutputS6xD(284)(1);
  VNStageIntLLRInputS6xD(188)(3) <= CNStageIntLLROutputS6xD(284)(2);
  VNStageIntLLRInputS6xD(239)(5) <= CNStageIntLLROutputS6xD(284)(3);
  VNStageIntLLRInputS6xD(294)(5) <= CNStageIntLLROutputS6xD(284)(4);
  VNStageIntLLRInputS6xD(325)(5) <= CNStageIntLLROutputS6xD(284)(5);
  VNStageIntLLRInputS6xD(27)(4) <= CNStageIntLLROutputS6xD(285)(0);
  VNStageIntLLRInputS6xD(99)(5) <= CNStageIntLLROutputS6xD(285)(1);
  VNStageIntLLRInputS6xD(130)(5) <= CNStageIntLLROutputS6xD(285)(2);
  VNStageIntLLRInputS6xD(241)(4) <= CNStageIntLLROutputS6xD(285)(3);
  VNStageIntLLRInputS6xD(273)(4) <= CNStageIntLLROutputS6xD(285)(4);
  VNStageIntLLRInputS6xD(361)(5) <= CNStageIntLLROutputS6xD(285)(5);
  VNStageIntLLRInputS6xD(26)(5) <= CNStageIntLLROutputS6xD(286)(0);
  VNStageIntLLRInputS6xD(65)(4) <= CNStageIntLLROutputS6xD(286)(1);
  VNStageIntLLRInputS6xD(176)(5) <= CNStageIntLLROutputS6xD(286)(2);
  VNStageIntLLRInputS6xD(208)(4) <= CNStageIntLLROutputS6xD(286)(3);
  VNStageIntLLRInputS6xD(296)(4) <= CNStageIntLLROutputS6xD(286)(4);
  VNStageIntLLRInputS6xD(334)(3) <= CNStageIntLLROutputS6xD(286)(5);
  VNStageIntLLRInputS6xD(25)(4) <= CNStageIntLLROutputS6xD(287)(0);
  VNStageIntLLRInputS6xD(111)(5) <= CNStageIntLLROutputS6xD(287)(1);
  VNStageIntLLRInputS6xD(143)(5) <= CNStageIntLLROutputS6xD(287)(2);
  VNStageIntLLRInputS6xD(231)(4) <= CNStageIntLLROutputS6xD(287)(3);
  VNStageIntLLRInputS6xD(269)(4) <= CNStageIntLLROutputS6xD(287)(4);
  VNStageIntLLRInputS6xD(381)(4) <= CNStageIntLLROutputS6xD(287)(5);
  VNStageIntLLRInputS6xD(24)(5) <= CNStageIntLLROutputS6xD(288)(0);
  VNStageIntLLRInputS6xD(78)(5) <= CNStageIntLLROutputS6xD(288)(1);
  VNStageIntLLRInputS6xD(166)(4) <= CNStageIntLLROutputS6xD(288)(2);
  VNStageIntLLRInputS6xD(204)(5) <= CNStageIntLLROutputS6xD(288)(3);
  VNStageIntLLRInputS6xD(316)(3) <= CNStageIntLLROutputS6xD(288)(4);
  VNStageIntLLRInputS6xD(321)(5) <= CNStageIntLLROutputS6xD(288)(5);
  VNStageIntLLRInputS6xD(23)(5) <= CNStageIntLLROutputS6xD(289)(0);
  VNStageIntLLRInputS6xD(101)(5) <= CNStageIntLLROutputS6xD(289)(1);
  VNStageIntLLRInputS6xD(139)(5) <= CNStageIntLLROutputS6xD(289)(2);
  VNStageIntLLRInputS6xD(251)(3) <= CNStageIntLLROutputS6xD(289)(3);
  VNStageIntLLRInputS6xD(319)(5) <= CNStageIntLLROutputS6xD(289)(4);
  VNStageIntLLRInputS6xD(362)(5) <= CNStageIntLLROutputS6xD(289)(5);
  VNStageIntLLRInputS6xD(22)(5) <= CNStageIntLLROutputS6xD(290)(0);
  VNStageIntLLRInputS6xD(74)(4) <= CNStageIntLLROutputS6xD(290)(1);
  VNStageIntLLRInputS6xD(186)(4) <= CNStageIntLLROutputS6xD(290)(2);
  VNStageIntLLRInputS6xD(254)(3) <= CNStageIntLLROutputS6xD(290)(3);
  VNStageIntLLRInputS6xD(297)(5) <= CNStageIntLLROutputS6xD(290)(4);
  VNStageIntLLRInputS6xD(337)(5) <= CNStageIntLLROutputS6xD(290)(5);
  VNStageIntLLRInputS6xD(21)(5) <= CNStageIntLLROutputS6xD(291)(0);
  VNStageIntLLRInputS6xD(121)(4) <= CNStageIntLLROutputS6xD(291)(1);
  VNStageIntLLRInputS6xD(189)(4) <= CNStageIntLLROutputS6xD(291)(2);
  VNStageIntLLRInputS6xD(232)(4) <= CNStageIntLLROutputS6xD(291)(3);
  VNStageIntLLRInputS6xD(272)(5) <= CNStageIntLLROutputS6xD(291)(4);
  VNStageIntLLRInputS6xD(335)(5) <= CNStageIntLLROutputS6xD(291)(5);
  VNStageIntLLRInputS6xD(20)(3) <= CNStageIntLLROutputS6xD(292)(0);
  VNStageIntLLRInputS6xD(124)(3) <= CNStageIntLLROutputS6xD(292)(1);
  VNStageIntLLRInputS6xD(167)(5) <= CNStageIntLLROutputS6xD(292)(2);
  VNStageIntLLRInputS6xD(207)(4) <= CNStageIntLLROutputS6xD(292)(3);
  VNStageIntLLRInputS6xD(270)(5) <= CNStageIntLLROutputS6xD(292)(4);
  VNStageIntLLRInputS6xD(360)(5) <= CNStageIntLLROutputS6xD(292)(5);
  VNStageIntLLRInputS6xD(18)(5) <= CNStageIntLLROutputS6xD(293)(0);
  VNStageIntLLRInputS6xD(77)(3) <= CNStageIntLLROutputS6xD(293)(1);
  VNStageIntLLRInputS6xD(140)(5) <= CNStageIntLLROutputS6xD(293)(2);
  VNStageIntLLRInputS6xD(230)(4) <= CNStageIntLLROutputS6xD(293)(3);
  VNStageIntLLRInputS6xD(303)(5) <= CNStageIntLLROutputS6xD(293)(4);
  VNStageIntLLRInputS6xD(348)(5) <= CNStageIntLLROutputS6xD(293)(5);
  VNStageIntLLRInputS6xD(17)(5) <= CNStageIntLLROutputS6xD(294)(0);
  VNStageIntLLRInputS6xD(75)(5) <= CNStageIntLLROutputS6xD(294)(1);
  VNStageIntLLRInputS6xD(165)(4) <= CNStageIntLLROutputS6xD(294)(2);
  VNStageIntLLRInputS6xD(238)(5) <= CNStageIntLLROutputS6xD(294)(3);
  VNStageIntLLRInputS6xD(283)(5) <= CNStageIntLLROutputS6xD(294)(4);
  VNStageIntLLRInputS6xD(342)(4) <= CNStageIntLLROutputS6xD(294)(5);
  VNStageIntLLRInputS6xD(16)(4) <= CNStageIntLLROutputS6xD(295)(0);
  VNStageIntLLRInputS6xD(100)(5) <= CNStageIntLLROutputS6xD(295)(1);
  VNStageIntLLRInputS6xD(173)(5) <= CNStageIntLLROutputS6xD(295)(2);
  VNStageIntLLRInputS6xD(218)(5) <= CNStageIntLLROutputS6xD(295)(3);
  VNStageIntLLRInputS6xD(277)(5) <= CNStageIntLLROutputS6xD(295)(4);
  VNStageIntLLRInputS6xD(320)(3) <= CNStageIntLLROutputS6xD(295)(5);
  VNStageIntLLRInputS6xD(15)(5) <= CNStageIntLLROutputS6xD(296)(0);
  VNStageIntLLRInputS6xD(108)(5) <= CNStageIntLLROutputS6xD(296)(1);
  VNStageIntLLRInputS6xD(153)(5) <= CNStageIntLLROutputS6xD(296)(2);
  VNStageIntLLRInputS6xD(212)(4) <= CNStageIntLLROutputS6xD(296)(3);
  VNStageIntLLRInputS6xD(256)(4) <= CNStageIntLLROutputS6xD(296)(4);
  VNStageIntLLRInputS6xD(341)(5) <= CNStageIntLLROutputS6xD(296)(5);
  VNStageIntLLRInputS6xD(14)(5) <= CNStageIntLLROutputS6xD(297)(0);
  VNStageIntLLRInputS6xD(88)(5) <= CNStageIntLLROutputS6xD(297)(1);
  VNStageIntLLRInputS6xD(147)(5) <= CNStageIntLLROutputS6xD(297)(2);
  VNStageIntLLRInputS6xD(192)(5) <= CNStageIntLLROutputS6xD(297)(3);
  VNStageIntLLRInputS6xD(276)(5) <= CNStageIntLLROutputS6xD(297)(4);
  VNStageIntLLRInputS6xD(346)(5) <= CNStageIntLLROutputS6xD(297)(5);
  VNStageIntLLRInputS6xD(13)(4) <= CNStageIntLLROutputS6xD(298)(0);
  VNStageIntLLRInputS6xD(82)(5) <= CNStageIntLLROutputS6xD(298)(1);
  VNStageIntLLRInputS6xD(128)(5) <= CNStageIntLLROutputS6xD(298)(2);
  VNStageIntLLRInputS6xD(211)(5) <= CNStageIntLLROutputS6xD(298)(3);
  VNStageIntLLRInputS6xD(281)(5) <= CNStageIntLLROutputS6xD(298)(4);
  VNStageIntLLRInputS6xD(365)(5) <= CNStageIntLLROutputS6xD(298)(5);
  VNStageIntLLRInputS6xD(12)(5) <= CNStageIntLLROutputS6xD(299)(0);
  VNStageIntLLRInputS6xD(64)(4) <= CNStageIntLLROutputS6xD(299)(1);
  VNStageIntLLRInputS6xD(146)(4) <= CNStageIntLLROutputS6xD(299)(2);
  VNStageIntLLRInputS6xD(216)(5) <= CNStageIntLLROutputS6xD(299)(3);
  VNStageIntLLRInputS6xD(300)(4) <= CNStageIntLLROutputS6xD(299)(4);
  VNStageIntLLRInputS6xD(356)(4) <= CNStageIntLLROutputS6xD(299)(5);
  VNStageIntLLRInputS6xD(9)(5) <= CNStageIntLLROutputS6xD(300)(0);
  VNStageIntLLRInputS6xD(105)(4) <= CNStageIntLLROutputS6xD(300)(1);
  VNStageIntLLRInputS6xD(161)(5) <= CNStageIntLLROutputS6xD(300)(2);
  VNStageIntLLRInputS6xD(200)(5) <= CNStageIntLLROutputS6xD(300)(3);
  VNStageIntLLRInputS6xD(266)(4) <= CNStageIntLLROutputS6xD(300)(4);
  VNStageIntLLRInputS6xD(355)(5) <= CNStageIntLLROutputS6xD(300)(5);
  VNStageIntLLRInputS6xD(7)(5) <= CNStageIntLLROutputS6xD(301)(0);
  VNStageIntLLRInputS6xD(70)(5) <= CNStageIntLLROutputS6xD(301)(1);
  VNStageIntLLRInputS6xD(136)(5) <= CNStageIntLLROutputS6xD(301)(2);
  VNStageIntLLRInputS6xD(225)(5) <= CNStageIntLLROutputS6xD(301)(3);
  VNStageIntLLRInputS6xD(311)(4) <= CNStageIntLLROutputS6xD(301)(4);
  VNStageIntLLRInputS6xD(372)(4) <= CNStageIntLLROutputS6xD(301)(5);
  VNStageIntLLRInputS6xD(6)(5) <= CNStageIntLLROutputS6xD(302)(0);
  VNStageIntLLRInputS6xD(71)(4) <= CNStageIntLLROutputS6xD(302)(1);
  VNStageIntLLRInputS6xD(160)(5) <= CNStageIntLLROutputS6xD(302)(2);
  VNStageIntLLRInputS6xD(246)(5) <= CNStageIntLLROutputS6xD(302)(3);
  VNStageIntLLRInputS6xD(307)(5) <= CNStageIntLLROutputS6xD(302)(4);
  VNStageIntLLRInputS6xD(324)(5) <= CNStageIntLLROutputS6xD(302)(5);
  VNStageIntLLRInputS6xD(5)(5) <= CNStageIntLLROutputS6xD(303)(0);
  VNStageIntLLRInputS6xD(95)(5) <= CNStageIntLLROutputS6xD(303)(1);
  VNStageIntLLRInputS6xD(181)(5) <= CNStageIntLLROutputS6xD(303)(2);
  VNStageIntLLRInputS6xD(242)(5) <= CNStageIntLLROutputS6xD(303)(3);
  VNStageIntLLRInputS6xD(259)(3) <= CNStageIntLLROutputS6xD(303)(4);
  VNStageIntLLRInputS6xD(350)(5) <= CNStageIntLLROutputS6xD(303)(5);
  VNStageIntLLRInputS6xD(4)(4) <= CNStageIntLLROutputS6xD(304)(0);
  VNStageIntLLRInputS6xD(116)(4) <= CNStageIntLLROutputS6xD(304)(1);
  VNStageIntLLRInputS6xD(177)(5) <= CNStageIntLLROutputS6xD(304)(2);
  VNStageIntLLRInputS6xD(194)(5) <= CNStageIntLLROutputS6xD(304)(3);
  VNStageIntLLRInputS6xD(285)(5) <= CNStageIntLLROutputS6xD(304)(4);
  VNStageIntLLRInputS6xD(326)(4) <= CNStageIntLLROutputS6xD(304)(5);
  VNStageIntLLRInputS6xD(3)(4) <= CNStageIntLLROutputS6xD(305)(0);
  VNStageIntLLRInputS6xD(112)(5) <= CNStageIntLLROutputS6xD(305)(1);
  VNStageIntLLRInputS6xD(129)(5) <= CNStageIntLLROutputS6xD(305)(2);
  VNStageIntLLRInputS6xD(220)(5) <= CNStageIntLLROutputS6xD(305)(3);
  VNStageIntLLRInputS6xD(261)(4) <= CNStageIntLLROutputS6xD(305)(4);
  VNStageIntLLRInputS6xD(358)(4) <= CNStageIntLLROutputS6xD(305)(5);
  VNStageIntLLRInputS6xD(2)(5) <= CNStageIntLLROutputS6xD(306)(0);
  VNStageIntLLRInputS6xD(127)(5) <= CNStageIntLLROutputS6xD(306)(1);
  VNStageIntLLRInputS6xD(155)(5) <= CNStageIntLLROutputS6xD(306)(2);
  VNStageIntLLRInputS6xD(196)(5) <= CNStageIntLLROutputS6xD(306)(3);
  VNStageIntLLRInputS6xD(293)(4) <= CNStageIntLLROutputS6xD(306)(4);
  VNStageIntLLRInputS6xD(374)(5) <= CNStageIntLLROutputS6xD(306)(5);
  VNStageIntLLRInputS6xD(1)(4) <= CNStageIntLLROutputS6xD(307)(0);
  VNStageIntLLRInputS6xD(90)(5) <= CNStageIntLLROutputS6xD(307)(1);
  VNStageIntLLRInputS6xD(131)(4) <= CNStageIntLLROutputS6xD(307)(2);
  VNStageIntLLRInputS6xD(228)(5) <= CNStageIntLLROutputS6xD(307)(3);
  VNStageIntLLRInputS6xD(309)(5) <= CNStageIntLLROutputS6xD(307)(4);
  VNStageIntLLRInputS6xD(344)(5) <= CNStageIntLLROutputS6xD(307)(5);
  VNStageIntLLRInputS6xD(62)(4) <= CNStageIntLLROutputS6xD(308)(0);
  VNStageIntLLRInputS6xD(98)(4) <= CNStageIntLLROutputS6xD(308)(1);
  VNStageIntLLRInputS6xD(179)(5) <= CNStageIntLLROutputS6xD(308)(2);
  VNStageIntLLRInputS6xD(214)(5) <= CNStageIntLLROutputS6xD(308)(3);
  VNStageIntLLRInputS6xD(288)(5) <= CNStageIntLLROutputS6xD(308)(4);
  VNStageIntLLRInputS6xD(366)(5) <= CNStageIntLLROutputS6xD(308)(5);
  VNStageIntLLRInputS6xD(61)(4) <= CNStageIntLLROutputS6xD(309)(0);
  VNStageIntLLRInputS6xD(114)(5) <= CNStageIntLLROutputS6xD(309)(1);
  VNStageIntLLRInputS6xD(149)(5) <= CNStageIntLLROutputS6xD(309)(2);
  VNStageIntLLRInputS6xD(223)(5) <= CNStageIntLLROutputS6xD(309)(3);
  VNStageIntLLRInputS6xD(301)(5) <= CNStageIntLLROutputS6xD(309)(4);
  VNStageIntLLRInputS6xD(345)(4) <= CNStageIntLLROutputS6xD(309)(5);
  VNStageIntLLRInputS6xD(60)(4) <= CNStageIntLLROutputS6xD(310)(0);
  VNStageIntLLRInputS6xD(84)(4) <= CNStageIntLLROutputS6xD(310)(1);
  VNStageIntLLRInputS6xD(158)(5) <= CNStageIntLLROutputS6xD(310)(2);
  VNStageIntLLRInputS6xD(236)(5) <= CNStageIntLLROutputS6xD(310)(3);
  VNStageIntLLRInputS6xD(280)(5) <= CNStageIntLLROutputS6xD(310)(4);
  VNStageIntLLRInputS6xD(373)(3) <= CNStageIntLLROutputS6xD(310)(5);
  VNStageIntLLRInputS6xD(59)(3) <= CNStageIntLLROutputS6xD(311)(0);
  VNStageIntLLRInputS6xD(93)(5) <= CNStageIntLLROutputS6xD(311)(1);
  VNStageIntLLRInputS6xD(171)(3) <= CNStageIntLLROutputS6xD(311)(2);
  VNStageIntLLRInputS6xD(215)(5) <= CNStageIntLLROutputS6xD(311)(3);
  VNStageIntLLRInputS6xD(308)(3) <= CNStageIntLLROutputS6xD(311)(4);
  VNStageIntLLRInputS6xD(375)(4) <= CNStageIntLLROutputS6xD(311)(5);
  VNStageIntLLRInputS6xD(58)(3) <= CNStageIntLLROutputS6xD(312)(0);
  VNStageIntLLRInputS6xD(106)(4) <= CNStageIntLLROutputS6xD(312)(1);
  VNStageIntLLRInputS6xD(150)(4) <= CNStageIntLLROutputS6xD(312)(2);
  VNStageIntLLRInputS6xD(243)(5) <= CNStageIntLLROutputS6xD(312)(3);
  VNStageIntLLRInputS6xD(310)(4) <= CNStageIntLLROutputS6xD(312)(4);
  VNStageIntLLRInputS6xD(357)(5) <= CNStageIntLLROutputS6xD(312)(5);
  VNStageIntLLRInputS6xD(57)(4) <= CNStageIntLLROutputS6xD(313)(0);
  VNStageIntLLRInputS6xD(85)(4) <= CNStageIntLLROutputS6xD(313)(1);
  VNStageIntLLRInputS6xD(178)(4) <= CNStageIntLLROutputS6xD(313)(2);
  VNStageIntLLRInputS6xD(245)(5) <= CNStageIntLLROutputS6xD(313)(3);
  VNStageIntLLRInputS6xD(292)(5) <= CNStageIntLLROutputS6xD(313)(4);
  VNStageIntLLRInputS6xD(364)(5) <= CNStageIntLLROutputS6xD(313)(5);
  VNStageIntLLRInputS6xD(56)(5) <= CNStageIntLLROutputS6xD(314)(0);
  VNStageIntLLRInputS6xD(113)(5) <= CNStageIntLLROutputS6xD(314)(1);
  VNStageIntLLRInputS6xD(180)(3) <= CNStageIntLLROutputS6xD(314)(2);
  VNStageIntLLRInputS6xD(227)(5) <= CNStageIntLLROutputS6xD(314)(3);
  VNStageIntLLRInputS6xD(299)(4) <= CNStageIntLLROutputS6xD(314)(4);
  VNStageIntLLRInputS6xD(328)(3) <= CNStageIntLLROutputS6xD(314)(5);
  VNStageIntLLRInputS6xD(55)(5) <= CNStageIntLLROutputS6xD(315)(0);
  VNStageIntLLRInputS6xD(115)(5) <= CNStageIntLLROutputS6xD(315)(1);
  VNStageIntLLRInputS6xD(162)(5) <= CNStageIntLLROutputS6xD(315)(2);
  VNStageIntLLRInputS6xD(234)(5) <= CNStageIntLLROutputS6xD(315)(3);
  VNStageIntLLRInputS6xD(263)(5) <= CNStageIntLLROutputS6xD(315)(4);
  VNStageIntLLRInputS6xD(379)(3) <= CNStageIntLLROutputS6xD(315)(5);
  VNStageIntLLRInputS6xD(54)(4) <= CNStageIntLLROutputS6xD(316)(0);
  VNStageIntLLRInputS6xD(97)(5) <= CNStageIntLLROutputS6xD(316)(1);
  VNStageIntLLRInputS6xD(169)(5) <= CNStageIntLLROutputS6xD(316)(2);
  VNStageIntLLRInputS6xD(198)(5) <= CNStageIntLLROutputS6xD(316)(3);
  VNStageIntLLRInputS6xD(314)(2) <= CNStageIntLLROutputS6xD(316)(4);
  VNStageIntLLRInputS6xD(322)(4) <= CNStageIntLLROutputS6xD(316)(5);
  VNStageIntLLRInputS6xD(53)(4) <= CNStageIntLLROutputS6xD(317)(0);
  VNStageIntLLRInputS6xD(104)(5) <= CNStageIntLLROutputS6xD(317)(1);
  VNStageIntLLRInputS6xD(133)(3) <= CNStageIntLLROutputS6xD(317)(2);
  VNStageIntLLRInputS6xD(249)(3) <= CNStageIntLLROutputS6xD(317)(3);
  VNStageIntLLRInputS6xD(257)(5) <= CNStageIntLLROutputS6xD(317)(4);
  VNStageIntLLRInputS6xD(380)(4) <= CNStageIntLLROutputS6xD(317)(5);
  VNStageIntLLRInputS6xD(52)(3) <= CNStageIntLLROutputS6xD(318)(0);
  VNStageIntLLRInputS6xD(68)(4) <= CNStageIntLLROutputS6xD(318)(1);
  VNStageIntLLRInputS6xD(184)(5) <= CNStageIntLLROutputS6xD(318)(2);
  VNStageIntLLRInputS6xD(255)(5) <= CNStageIntLLROutputS6xD(318)(3);
  VNStageIntLLRInputS6xD(315)(4) <= CNStageIntLLROutputS6xD(318)(4);
  VNStageIntLLRInputS6xD(327)(5) <= CNStageIntLLROutputS6xD(318)(5);
  VNStageIntLLRInputS6xD(51)(4) <= CNStageIntLLROutputS6xD(319)(0);
  VNStageIntLLRInputS6xD(119)(4) <= CNStageIntLLROutputS6xD(319)(1);
  VNStageIntLLRInputS6xD(190)(3) <= CNStageIntLLROutputS6xD(319)(2);
  VNStageIntLLRInputS6xD(250)(3) <= CNStageIntLLROutputS6xD(319)(3);
  VNStageIntLLRInputS6xD(262)(4) <= CNStageIntLLROutputS6xD(319)(4);
  VNStageIntLLRInputS6xD(349)(4) <= CNStageIntLLROutputS6xD(319)(5);
  VNStageIntLLRInputS6xD(50)(5) <= CNStageIntLLROutputS6xD(320)(0);
  VNStageIntLLRInputS6xD(125)(2) <= CNStageIntLLROutputS6xD(320)(1);
  VNStageIntLLRInputS6xD(185)(2) <= CNStageIntLLROutputS6xD(320)(2);
  VNStageIntLLRInputS6xD(197)(5) <= CNStageIntLLROutputS6xD(320)(3);
  VNStageIntLLRInputS6xD(284)(5) <= CNStageIntLLROutputS6xD(320)(4);
  VNStageIntLLRInputS6xD(367)(5) <= CNStageIntLLROutputS6xD(320)(5);
  VNStageIntLLRInputS6xD(49)(5) <= CNStageIntLLROutputS6xD(321)(0);
  VNStageIntLLRInputS6xD(120)(2) <= CNStageIntLLROutputS6xD(321)(1);
  VNStageIntLLRInputS6xD(132)(4) <= CNStageIntLLROutputS6xD(321)(2);
  VNStageIntLLRInputS6xD(219)(4) <= CNStageIntLLROutputS6xD(321)(3);
  VNStageIntLLRInputS6xD(302)(5) <= CNStageIntLLROutputS6xD(321)(4);
  VNStageIntLLRInputS6xD(352)(5) <= CNStageIntLLROutputS6xD(321)(5);
  VNStageIntLLRInputS6xD(48)(2) <= CNStageIntLLROutputS6xD(322)(0);
  VNStageIntLLRInputS6xD(67)(2) <= CNStageIntLLROutputS6xD(322)(1);
  VNStageIntLLRInputS6xD(154)(4) <= CNStageIntLLROutputS6xD(322)(2);
  VNStageIntLLRInputS6xD(237)(4) <= CNStageIntLLROutputS6xD(322)(3);
  VNStageIntLLRInputS6xD(287)(5) <= CNStageIntLLROutputS6xD(322)(4);
  VNStageIntLLRInputS6xD(339)(5) <= CNStageIntLLROutputS6xD(322)(5);
  VNStageIntLLRInputS6xD(46)(5) <= CNStageIntLLROutputS6xD(323)(0);
  VNStageIntLLRInputS6xD(107)(4) <= CNStageIntLLROutputS6xD(323)(1);
  VNStageIntLLRInputS6xD(157)(4) <= CNStageIntLLROutputS6xD(323)(2);
  VNStageIntLLRInputS6xD(209)(4) <= CNStageIntLLROutputS6xD(323)(3);
  VNStageIntLLRInputS6xD(305)(5) <= CNStageIntLLROutputS6xD(323)(4);
  VNStageIntLLRInputS6xD(382)(4) <= CNStageIntLLROutputS6xD(323)(5);
  VNStageIntLLRInputS6xD(45)(5) <= CNStageIntLLROutputS6xD(324)(0);
  VNStageIntLLRInputS6xD(92)(5) <= CNStageIntLLROutputS6xD(324)(1);
  VNStageIntLLRInputS6xD(144)(5) <= CNStageIntLLROutputS6xD(324)(2);
  VNStageIntLLRInputS6xD(240)(5) <= CNStageIntLLROutputS6xD(324)(3);
  VNStageIntLLRInputS6xD(317)(2) <= CNStageIntLLROutputS6xD(324)(4);
  VNStageIntLLRInputS6xD(333)(4) <= CNStageIntLLROutputS6xD(324)(5);
  VNStageIntLLRInputS6xD(44)(5) <= CNStageIntLLROutputS6xD(325)(0);
  VNStageIntLLRInputS6xD(79)(4) <= CNStageIntLLROutputS6xD(325)(1);
  VNStageIntLLRInputS6xD(175)(5) <= CNStageIntLLROutputS6xD(325)(2);
  VNStageIntLLRInputS6xD(252)(4) <= CNStageIntLLROutputS6xD(325)(3);
  VNStageIntLLRInputS6xD(268)(5) <= CNStageIntLLROutputS6xD(325)(4);
  VNStageIntLLRInputS6xD(377)(3) <= CNStageIntLLROutputS6xD(325)(5);
  VNStageIntLLRInputS6xD(43)(4) <= CNStageIntLLROutputS6xD(326)(0);
  VNStageIntLLRInputS6xD(110)(5) <= CNStageIntLLROutputS6xD(326)(1);
  VNStageIntLLRInputS6xD(187)(4) <= CNStageIntLLROutputS6xD(326)(2);
  VNStageIntLLRInputS6xD(203)(5) <= CNStageIntLLROutputS6xD(326)(3);
  VNStageIntLLRInputS6xD(312)(4) <= CNStageIntLLROutputS6xD(326)(4);
  VNStageIntLLRInputS6xD(354)(4) <= CNStageIntLLROutputS6xD(326)(5);
  VNStageIntLLRInputS6xD(42)(5) <= CNStageIntLLROutputS6xD(327)(0);
  VNStageIntLLRInputS6xD(122)(4) <= CNStageIntLLROutputS6xD(327)(1);
  VNStageIntLLRInputS6xD(138)(5) <= CNStageIntLLROutputS6xD(327)(2);
  VNStageIntLLRInputS6xD(247)(5) <= CNStageIntLLROutputS6xD(327)(3);
  VNStageIntLLRInputS6xD(289)(5) <= CNStageIntLLROutputS6xD(327)(4);
  VNStageIntLLRInputS6xD(343)(5) <= CNStageIntLLROutputS6xD(327)(5);
  VNStageIntLLRInputS6xD(41)(5) <= CNStageIntLLROutputS6xD(328)(0);
  VNStageIntLLRInputS6xD(73)(4) <= CNStageIntLLROutputS6xD(328)(1);
  VNStageIntLLRInputS6xD(182)(5) <= CNStageIntLLROutputS6xD(328)(2);
  VNStageIntLLRInputS6xD(224)(5) <= CNStageIntLLROutputS6xD(328)(3);
  VNStageIntLLRInputS6xD(278)(4) <= CNStageIntLLROutputS6xD(328)(4);
  VNStageIntLLRInputS6xD(347)(5) <= CNStageIntLLROutputS6xD(328)(5);
  VNStageIntLLRInputS6xD(39)(5) <= CNStageIntLLROutputS6xD(329)(0);
  VNStageIntLLRInputS6xD(94)(3) <= CNStageIntLLROutputS6xD(329)(1);
  VNStageIntLLRInputS6xD(148)(5) <= CNStageIntLLROutputS6xD(329)(2);
  VNStageIntLLRInputS6xD(217)(5) <= CNStageIntLLROutputS6xD(329)(3);
  VNStageIntLLRInputS6xD(275)(4) <= CNStageIntLLROutputS6xD(329)(4);
  VNStageIntLLRInputS6xD(351)(4) <= CNStageIntLLROutputS6xD(329)(5);
  VNStageIntLLRInputS6xD(38)(5) <= CNStageIntLLROutputS6xD(330)(0);
  VNStageIntLLRInputS6xD(83)(5) <= CNStageIntLLROutputS6xD(330)(1);
  VNStageIntLLRInputS6xD(152)(5) <= CNStageIntLLROutputS6xD(330)(2);
  VNStageIntLLRInputS6xD(210)(5) <= CNStageIntLLROutputS6xD(330)(3);
  VNStageIntLLRInputS6xD(286)(5) <= CNStageIntLLROutputS6xD(330)(4);
  VNStageIntLLRInputS6xD(323)(4) <= CNStageIntLLROutputS6xD(330)(5);
  VNStageIntLLRInputS6xD(37)(5) <= CNStageIntLLROutputS6xD(331)(0);
  VNStageIntLLRInputS6xD(87)(5) <= CNStageIntLLROutputS6xD(331)(1);
  VNStageIntLLRInputS6xD(145)(5) <= CNStageIntLLROutputS6xD(331)(2);
  VNStageIntLLRInputS6xD(221)(5) <= CNStageIntLLROutputS6xD(331)(3);
  VNStageIntLLRInputS6xD(258)(2) <= CNStageIntLLROutputS6xD(331)(4);
  VNStageIntLLRInputS6xD(378)(4) <= CNStageIntLLROutputS6xD(331)(5);
  VNStageIntLLRInputS6xD(0)(5) <= CNStageIntLLROutputS6xD(332)(0);
  VNStageIntLLRInputS6xD(76)(5) <= CNStageIntLLROutputS6xD(332)(1);
  VNStageIntLLRInputS6xD(141)(3) <= CNStageIntLLROutputS6xD(332)(2);
  VNStageIntLLRInputS6xD(206)(3) <= CNStageIntLLROutputS6xD(332)(3);
  VNStageIntLLRInputS6xD(271)(4) <= CNStageIntLLROutputS6xD(332)(4);
  VNStageIntLLRInputS6xD(336)(4) <= CNStageIntLLROutputS6xD(332)(5);
  VNStageIntLLRInputS6xD(28)(5) <= CNStageIntLLROutputS6xD(333)(0);
  VNStageIntLLRInputS6xD(106)(5) <= CNStageIntLLROutputS6xD(333)(1);
  VNStageIntLLRInputS6xD(144)(6) <= CNStageIntLLROutputS6xD(333)(2);
  VNStageIntLLRInputS6xD(193)(4) <= CNStageIntLLROutputS6xD(333)(3);
  VNStageIntLLRInputS6xD(261)(5) <= CNStageIntLLROutputS6xD(333)(4);
  VNStageIntLLRInputS6xD(367)(6) <= CNStageIntLLROutputS6xD(333)(5);
  VNStageIntLLRInputS6xD(26)(6) <= CNStageIntLLROutputS6xD(334)(0);
  VNStageIntLLRInputS6xD(126)(5) <= CNStageIntLLROutputS6xD(334)(1);
  VNStageIntLLRInputS6xD(131)(5) <= CNStageIntLLROutputS6xD(334)(2);
  VNStageIntLLRInputS6xD(237)(5) <= CNStageIntLLROutputS6xD(334)(3);
  VNStageIntLLRInputS6xD(277)(6) <= CNStageIntLLROutputS6xD(334)(4);
  VNStageIntLLRInputS6xD(340)(5) <= CNStageIntLLROutputS6xD(334)(5);
  VNStageIntLLRInputS6xD(24)(6) <= CNStageIntLLROutputS6xD(335)(0);
  VNStageIntLLRInputS6xD(107)(5) <= CNStageIntLLROutputS6xD(335)(1);
  VNStageIntLLRInputS6xD(147)(6) <= CNStageIntLLROutputS6xD(335)(2);
  VNStageIntLLRInputS6xD(210)(6) <= CNStageIntLLROutputS6xD(335)(3);
  VNStageIntLLRInputS6xD(300)(5) <= CNStageIntLLROutputS6xD(335)(4);
  VNStageIntLLRInputS6xD(373)(4) <= CNStageIntLLROutputS6xD(335)(5);
  VNStageIntLLRInputS6xD(23)(6) <= CNStageIntLLROutputS6xD(336)(0);
  VNStageIntLLRInputS6xD(82)(6) <= CNStageIntLLROutputS6xD(336)(1);
  VNStageIntLLRInputS6xD(145)(6) <= CNStageIntLLROutputS6xD(336)(2);
  VNStageIntLLRInputS6xD(235)(4) <= CNStageIntLLROutputS6xD(336)(3);
  VNStageIntLLRInputS6xD(308)(4) <= CNStageIntLLROutputS6xD(336)(4);
  VNStageIntLLRInputS6xD(353)(5) <= CNStageIntLLROutputS6xD(336)(5);
  VNStageIntLLRInputS6xD(22)(6) <= CNStageIntLLROutputS6xD(337)(0);
  VNStageIntLLRInputS6xD(80)(5) <= CNStageIntLLROutputS6xD(337)(1);
  VNStageIntLLRInputS6xD(170)(4) <= CNStageIntLLROutputS6xD(337)(2);
  VNStageIntLLRInputS6xD(243)(6) <= CNStageIntLLROutputS6xD(337)(3);
  VNStageIntLLRInputS6xD(288)(6) <= CNStageIntLLROutputS6xD(337)(4);
  VNStageIntLLRInputS6xD(347)(6) <= CNStageIntLLROutputS6xD(337)(5);
  VNStageIntLLRInputS6xD(21)(6) <= CNStageIntLLROutputS6xD(338)(0);
  VNStageIntLLRInputS6xD(105)(5) <= CNStageIntLLROutputS6xD(338)(1);
  VNStageIntLLRInputS6xD(178)(5) <= CNStageIntLLROutputS6xD(338)(2);
  VNStageIntLLRInputS6xD(223)(6) <= CNStageIntLLROutputS6xD(338)(3);
  VNStageIntLLRInputS6xD(282)(5) <= CNStageIntLLROutputS6xD(338)(4);
  VNStageIntLLRInputS6xD(320)(4) <= CNStageIntLLROutputS6xD(338)(5);
  VNStageIntLLRInputS6xD(20)(4) <= CNStageIntLLROutputS6xD(339)(0);
  VNStageIntLLRInputS6xD(113)(6) <= CNStageIntLLROutputS6xD(339)(1);
  VNStageIntLLRInputS6xD(158)(6) <= CNStageIntLLROutputS6xD(339)(2);
  VNStageIntLLRInputS6xD(217)(6) <= CNStageIntLLROutputS6xD(339)(3);
  VNStageIntLLRInputS6xD(256)(5) <= CNStageIntLLROutputS6xD(339)(4);
  VNStageIntLLRInputS6xD(346)(6) <= CNStageIntLLROutputS6xD(339)(5);
  VNStageIntLLRInputS6xD(19)(4) <= CNStageIntLLROutputS6xD(340)(0);
  VNStageIntLLRInputS6xD(93)(6) <= CNStageIntLLROutputS6xD(340)(1);
  VNStageIntLLRInputS6xD(152)(6) <= CNStageIntLLROutputS6xD(340)(2);
  VNStageIntLLRInputS6xD(192)(6) <= CNStageIntLLROutputS6xD(340)(3);
  VNStageIntLLRInputS6xD(281)(6) <= CNStageIntLLROutputS6xD(340)(4);
  VNStageIntLLRInputS6xD(351)(5) <= CNStageIntLLROutputS6xD(340)(5);
  VNStageIntLLRInputS6xD(18)(6) <= CNStageIntLLROutputS6xD(341)(0);
  VNStageIntLLRInputS6xD(87)(6) <= CNStageIntLLROutputS6xD(341)(1);
  VNStageIntLLRInputS6xD(128)(6) <= CNStageIntLLROutputS6xD(341)(2);
  VNStageIntLLRInputS6xD(216)(6) <= CNStageIntLLROutputS6xD(341)(3);
  VNStageIntLLRInputS6xD(286)(6) <= CNStageIntLLROutputS6xD(341)(4);
  VNStageIntLLRInputS6xD(370)(4) <= CNStageIntLLROutputS6xD(341)(5);
  VNStageIntLLRInputS6xD(17)(6) <= CNStageIntLLROutputS6xD(342)(0);
  VNStageIntLLRInputS6xD(64)(5) <= CNStageIntLLROutputS6xD(342)(1);
  VNStageIntLLRInputS6xD(151)(5) <= CNStageIntLLROutputS6xD(342)(2);
  VNStageIntLLRInputS6xD(221)(6) <= CNStageIntLLROutputS6xD(342)(3);
  VNStageIntLLRInputS6xD(305)(6) <= CNStageIntLLROutputS6xD(342)(4);
  VNStageIntLLRInputS6xD(361)(6) <= CNStageIntLLROutputS6xD(342)(5);
  VNStageIntLLRInputS6xD(16)(5) <= CNStageIntLLROutputS6xD(343)(0);
  VNStageIntLLRInputS6xD(86)(3) <= CNStageIntLLROutputS6xD(343)(1);
  VNStageIntLLRInputS6xD(156)(3) <= CNStageIntLLROutputS6xD(343)(2);
  VNStageIntLLRInputS6xD(240)(6) <= CNStageIntLLROutputS6xD(343)(3);
  VNStageIntLLRInputS6xD(296)(5) <= CNStageIntLLROutputS6xD(343)(4);
  VNStageIntLLRInputS6xD(335)(6) <= CNStageIntLLROutputS6xD(343)(5);
  VNStageIntLLRInputS6xD(15)(6) <= CNStageIntLLROutputS6xD(344)(0);
  VNStageIntLLRInputS6xD(91)(6) <= CNStageIntLLROutputS6xD(344)(1);
  VNStageIntLLRInputS6xD(175)(6) <= CNStageIntLLROutputS6xD(344)(2);
  VNStageIntLLRInputS6xD(231)(5) <= CNStageIntLLROutputS6xD(344)(3);
  VNStageIntLLRInputS6xD(270)(6) <= CNStageIntLLROutputS6xD(344)(4);
  VNStageIntLLRInputS6xD(336)(5) <= CNStageIntLLROutputS6xD(344)(5);
  VNStageIntLLRInputS6xD(14)(6) <= CNStageIntLLROutputS6xD(345)(0);
  VNStageIntLLRInputS6xD(110)(6) <= CNStageIntLLROutputS6xD(345)(1);
  VNStageIntLLRInputS6xD(166)(5) <= CNStageIntLLROutputS6xD(345)(2);
  VNStageIntLLRInputS6xD(205)(2) <= CNStageIntLLROutputS6xD(345)(3);
  VNStageIntLLRInputS6xD(271)(5) <= CNStageIntLLROutputS6xD(345)(4);
  VNStageIntLLRInputS6xD(360)(6) <= CNStageIntLLROutputS6xD(345)(5);
  VNStageIntLLRInputS6xD(13)(5) <= CNStageIntLLROutputS6xD(346)(0);
  VNStageIntLLRInputS6xD(101)(6) <= CNStageIntLLROutputS6xD(346)(1);
  VNStageIntLLRInputS6xD(140)(6) <= CNStageIntLLROutputS6xD(346)(2);
  VNStageIntLLRInputS6xD(206)(4) <= CNStageIntLLROutputS6xD(346)(3);
  VNStageIntLLRInputS6xD(295)(4) <= CNStageIntLLROutputS6xD(346)(4);
  VNStageIntLLRInputS6xD(381)(5) <= CNStageIntLLROutputS6xD(346)(5);
  VNStageIntLLRInputS6xD(12)(6) <= CNStageIntLLROutputS6xD(347)(0);
  VNStageIntLLRInputS6xD(75)(6) <= CNStageIntLLROutputS6xD(347)(1);
  VNStageIntLLRInputS6xD(141)(4) <= CNStageIntLLROutputS6xD(347)(2);
  VNStageIntLLRInputS6xD(230)(5) <= CNStageIntLLROutputS6xD(347)(3);
  VNStageIntLLRInputS6xD(316)(4) <= CNStageIntLLROutputS6xD(347)(4);
  VNStageIntLLRInputS6xD(377)(4) <= CNStageIntLLROutputS6xD(347)(5);
  VNStageIntLLRInputS6xD(11)(5) <= CNStageIntLLROutputS6xD(348)(0);
  VNStageIntLLRInputS6xD(76)(6) <= CNStageIntLLROutputS6xD(348)(1);
  VNStageIntLLRInputS6xD(165)(5) <= CNStageIntLLROutputS6xD(348)(2);
  VNStageIntLLRInputS6xD(251)(4) <= CNStageIntLLROutputS6xD(348)(3);
  VNStageIntLLRInputS6xD(312)(5) <= CNStageIntLLROutputS6xD(348)(4);
  VNStageIntLLRInputS6xD(329)(6) <= CNStageIntLLROutputS6xD(348)(5);
  VNStageIntLLRInputS6xD(10)(4) <= CNStageIntLLROutputS6xD(349)(0);
  VNStageIntLLRInputS6xD(100)(6) <= CNStageIntLLROutputS6xD(349)(1);
  VNStageIntLLRInputS6xD(186)(5) <= CNStageIntLLROutputS6xD(349)(2);
  VNStageIntLLRInputS6xD(247)(6) <= CNStageIntLLROutputS6xD(349)(3);
  VNStageIntLLRInputS6xD(264)(6) <= CNStageIntLLROutputS6xD(349)(4);
  VNStageIntLLRInputS6xD(355)(6) <= CNStageIntLLROutputS6xD(349)(5);
  VNStageIntLLRInputS6xD(9)(6) <= CNStageIntLLROutputS6xD(350)(0);
  VNStageIntLLRInputS6xD(121)(5) <= CNStageIntLLROutputS6xD(350)(1);
  VNStageIntLLRInputS6xD(182)(6) <= CNStageIntLLROutputS6xD(350)(2);
  VNStageIntLLRInputS6xD(199)(6) <= CNStageIntLLROutputS6xD(350)(3);
  VNStageIntLLRInputS6xD(290)(5) <= CNStageIntLLROutputS6xD(350)(4);
  VNStageIntLLRInputS6xD(331)(4) <= CNStageIntLLROutputS6xD(350)(5);
  VNStageIntLLRInputS6xD(7)(6) <= CNStageIntLLROutputS6xD(351)(0);
  VNStageIntLLRInputS6xD(69)(6) <= CNStageIntLLROutputS6xD(351)(1);
  VNStageIntLLRInputS6xD(160)(6) <= CNStageIntLLROutputS6xD(351)(2);
  VNStageIntLLRInputS6xD(201)(5) <= CNStageIntLLROutputS6xD(351)(3);
  VNStageIntLLRInputS6xD(298)(6) <= CNStageIntLLROutputS6xD(351)(4);
  VNStageIntLLRInputS6xD(379)(4) <= CNStageIntLLROutputS6xD(351)(5);
  VNStageIntLLRInputS6xD(6)(6) <= CNStageIntLLROutputS6xD(352)(0);
  VNStageIntLLRInputS6xD(95)(6) <= CNStageIntLLROutputS6xD(352)(1);
  VNStageIntLLRInputS6xD(136)(6) <= CNStageIntLLROutputS6xD(352)(2);
  VNStageIntLLRInputS6xD(233)(4) <= CNStageIntLLROutputS6xD(352)(3);
  VNStageIntLLRInputS6xD(314)(3) <= CNStageIntLLROutputS6xD(352)(4);
  VNStageIntLLRInputS6xD(349)(5) <= CNStageIntLLROutputS6xD(352)(5);
  VNStageIntLLRInputS6xD(5)(6) <= CNStageIntLLROutputS6xD(353)(0);
  VNStageIntLLRInputS6xD(71)(5) <= CNStageIntLLROutputS6xD(353)(1);
  VNStageIntLLRInputS6xD(168)(5) <= CNStageIntLLROutputS6xD(353)(2);
  VNStageIntLLRInputS6xD(249)(4) <= CNStageIntLLROutputS6xD(353)(3);
  VNStageIntLLRInputS6xD(284)(6) <= CNStageIntLLROutputS6xD(353)(4);
  VNStageIntLLRInputS6xD(358)(5) <= CNStageIntLLROutputS6xD(353)(5);
  VNStageIntLLRInputS6xD(4)(5) <= CNStageIntLLROutputS6xD(354)(0);
  VNStageIntLLRInputS6xD(103)(6) <= CNStageIntLLROutputS6xD(354)(1);
  VNStageIntLLRInputS6xD(184)(6) <= CNStageIntLLROutputS6xD(354)(2);
  VNStageIntLLRInputS6xD(219)(5) <= CNStageIntLLROutputS6xD(354)(3);
  VNStageIntLLRInputS6xD(293)(5) <= CNStageIntLLROutputS6xD(354)(4);
  VNStageIntLLRInputS6xD(371)(4) <= CNStageIntLLROutputS6xD(354)(5);
  VNStageIntLLRInputS6xD(2)(6) <= CNStageIntLLROutputS6xD(355)(0);
  VNStageIntLLRInputS6xD(89)(5) <= CNStageIntLLROutputS6xD(355)(1);
  VNStageIntLLRInputS6xD(163)(4) <= CNStageIntLLROutputS6xD(355)(2);
  VNStageIntLLRInputS6xD(241)(5) <= CNStageIntLLROutputS6xD(355)(3);
  VNStageIntLLRInputS6xD(285)(6) <= CNStageIntLLROutputS6xD(355)(4);
  VNStageIntLLRInputS6xD(378)(5) <= CNStageIntLLROutputS6xD(355)(5);
  VNStageIntLLRInputS6xD(1)(5) <= CNStageIntLLROutputS6xD(356)(0);
  VNStageIntLLRInputS6xD(98)(5) <= CNStageIntLLROutputS6xD(356)(1);
  VNStageIntLLRInputS6xD(176)(6) <= CNStageIntLLROutputS6xD(356)(2);
  VNStageIntLLRInputS6xD(220)(6) <= CNStageIntLLROutputS6xD(356)(3);
  VNStageIntLLRInputS6xD(313)(3) <= CNStageIntLLROutputS6xD(356)(4);
  VNStageIntLLRInputS6xD(380)(5) <= CNStageIntLLROutputS6xD(356)(5);
  VNStageIntLLRInputS6xD(63)(3) <= CNStageIntLLROutputS6xD(357)(0);
  VNStageIntLLRInputS6xD(111)(6) <= CNStageIntLLROutputS6xD(357)(1);
  VNStageIntLLRInputS6xD(155)(6) <= CNStageIntLLROutputS6xD(357)(2);
  VNStageIntLLRInputS6xD(248)(6) <= CNStageIntLLROutputS6xD(357)(3);
  VNStageIntLLRInputS6xD(315)(5) <= CNStageIntLLROutputS6xD(357)(4);
  VNStageIntLLRInputS6xD(362)(6) <= CNStageIntLLROutputS6xD(357)(5);
  VNStageIntLLRInputS6xD(62)(5) <= CNStageIntLLROutputS6xD(358)(0);
  VNStageIntLLRInputS6xD(90)(6) <= CNStageIntLLROutputS6xD(358)(1);
  VNStageIntLLRInputS6xD(183)(4) <= CNStageIntLLROutputS6xD(358)(2);
  VNStageIntLLRInputS6xD(250)(4) <= CNStageIntLLROutputS6xD(358)(3);
  VNStageIntLLRInputS6xD(297)(6) <= CNStageIntLLROutputS6xD(358)(4);
  VNStageIntLLRInputS6xD(369)(4) <= CNStageIntLLROutputS6xD(358)(5);
  VNStageIntLLRInputS6xD(61)(5) <= CNStageIntLLROutputS6xD(359)(0);
  VNStageIntLLRInputS6xD(118)(5) <= CNStageIntLLROutputS6xD(359)(1);
  VNStageIntLLRInputS6xD(185)(3) <= CNStageIntLLROutputS6xD(359)(2);
  VNStageIntLLRInputS6xD(232)(5) <= CNStageIntLLROutputS6xD(359)(3);
  VNStageIntLLRInputS6xD(304)(6) <= CNStageIntLLROutputS6xD(359)(4);
  VNStageIntLLRInputS6xD(333)(5) <= CNStageIntLLROutputS6xD(359)(5);
  VNStageIntLLRInputS6xD(60)(5) <= CNStageIntLLROutputS6xD(360)(0);
  VNStageIntLLRInputS6xD(120)(3) <= CNStageIntLLROutputS6xD(360)(1);
  VNStageIntLLRInputS6xD(167)(6) <= CNStageIntLLROutputS6xD(360)(2);
  VNStageIntLLRInputS6xD(239)(6) <= CNStageIntLLROutputS6xD(360)(3);
  VNStageIntLLRInputS6xD(268)(6) <= CNStageIntLLROutputS6xD(360)(4);
  VNStageIntLLRInputS6xD(321)(6) <= CNStageIntLLROutputS6xD(360)(5);
  VNStageIntLLRInputS6xD(59)(4) <= CNStageIntLLROutputS6xD(361)(0);
  VNStageIntLLRInputS6xD(102)(5) <= CNStageIntLLROutputS6xD(361)(1);
  VNStageIntLLRInputS6xD(174)(4) <= CNStageIntLLROutputS6xD(361)(2);
  VNStageIntLLRInputS6xD(203)(6) <= CNStageIntLLROutputS6xD(361)(3);
  VNStageIntLLRInputS6xD(319)(6) <= CNStageIntLLROutputS6xD(361)(4);
  VNStageIntLLRInputS6xD(327)(6) <= CNStageIntLLROutputS6xD(361)(5);
  VNStageIntLLRInputS6xD(58)(4) <= CNStageIntLLROutputS6xD(362)(0);
  VNStageIntLLRInputS6xD(109)(5) <= CNStageIntLLROutputS6xD(362)(1);
  VNStageIntLLRInputS6xD(138)(6) <= CNStageIntLLROutputS6xD(362)(2);
  VNStageIntLLRInputS6xD(254)(4) <= CNStageIntLLROutputS6xD(362)(3);
  VNStageIntLLRInputS6xD(262)(5) <= CNStageIntLLROutputS6xD(362)(4);
  VNStageIntLLRInputS6xD(322)(5) <= CNStageIntLLROutputS6xD(362)(5);
  VNStageIntLLRInputS6xD(57)(5) <= CNStageIntLLROutputS6xD(363)(0);
  VNStageIntLLRInputS6xD(73)(5) <= CNStageIntLLROutputS6xD(363)(1);
  VNStageIntLLRInputS6xD(189)(5) <= CNStageIntLLROutputS6xD(363)(2);
  VNStageIntLLRInputS6xD(197)(6) <= CNStageIntLLROutputS6xD(363)(3);
  VNStageIntLLRInputS6xD(257)(6) <= CNStageIntLLROutputS6xD(363)(4);
  VNStageIntLLRInputS6xD(332)(5) <= CNStageIntLLROutputS6xD(363)(5);
  VNStageIntLLRInputS6xD(56)(6) <= CNStageIntLLROutputS6xD(364)(0);
  VNStageIntLLRInputS6xD(124)(4) <= CNStageIntLLROutputS6xD(364)(1);
  VNStageIntLLRInputS6xD(132)(5) <= CNStageIntLLROutputS6xD(364)(2);
  VNStageIntLLRInputS6xD(255)(6) <= CNStageIntLLROutputS6xD(364)(3);
  VNStageIntLLRInputS6xD(267)(6) <= CNStageIntLLROutputS6xD(364)(4);
  VNStageIntLLRInputS6xD(354)(5) <= CNStageIntLLROutputS6xD(364)(5);
  VNStageIntLLRInputS6xD(55)(6) <= CNStageIntLLROutputS6xD(365)(0);
  VNStageIntLLRInputS6xD(67)(3) <= CNStageIntLLROutputS6xD(365)(1);
  VNStageIntLLRInputS6xD(190)(4) <= CNStageIntLLROutputS6xD(365)(2);
  VNStageIntLLRInputS6xD(202)(5) <= CNStageIntLLROutputS6xD(365)(3);
  VNStageIntLLRInputS6xD(289)(6) <= CNStageIntLLROutputS6xD(365)(4);
  VNStageIntLLRInputS6xD(372)(5) <= CNStageIntLLROutputS6xD(365)(5);
  VNStageIntLLRInputS6xD(54)(5) <= CNStageIntLLROutputS6xD(366)(0);
  VNStageIntLLRInputS6xD(125)(3) <= CNStageIntLLROutputS6xD(366)(1);
  VNStageIntLLRInputS6xD(137)(6) <= CNStageIntLLROutputS6xD(366)(2);
  VNStageIntLLRInputS6xD(224)(6) <= CNStageIntLLROutputS6xD(366)(3);
  VNStageIntLLRInputS6xD(307)(6) <= CNStageIntLLROutputS6xD(366)(4);
  VNStageIntLLRInputS6xD(357)(6) <= CNStageIntLLROutputS6xD(366)(5);
  VNStageIntLLRInputS6xD(53)(5) <= CNStageIntLLROutputS6xD(367)(0);
  VNStageIntLLRInputS6xD(72)(5) <= CNStageIntLLROutputS6xD(367)(1);
  VNStageIntLLRInputS6xD(159)(4) <= CNStageIntLLROutputS6xD(367)(2);
  VNStageIntLLRInputS6xD(242)(6) <= CNStageIntLLROutputS6xD(367)(3);
  VNStageIntLLRInputS6xD(292)(6) <= CNStageIntLLROutputS6xD(367)(4);
  VNStageIntLLRInputS6xD(344)(6) <= CNStageIntLLROutputS6xD(367)(5);
  VNStageIntLLRInputS6xD(52)(4) <= CNStageIntLLROutputS6xD(368)(0);
  VNStageIntLLRInputS6xD(94)(4) <= CNStageIntLLROutputS6xD(368)(1);
  VNStageIntLLRInputS6xD(177)(6) <= CNStageIntLLROutputS6xD(368)(2);
  VNStageIntLLRInputS6xD(227)(6) <= CNStageIntLLROutputS6xD(368)(3);
  VNStageIntLLRInputS6xD(279)(5) <= CNStageIntLLROutputS6xD(368)(4);
  VNStageIntLLRInputS6xD(375)(5) <= CNStageIntLLROutputS6xD(368)(5);
  VNStageIntLLRInputS6xD(51)(5) <= CNStageIntLLROutputS6xD(369)(0);
  VNStageIntLLRInputS6xD(112)(6) <= CNStageIntLLROutputS6xD(369)(1);
  VNStageIntLLRInputS6xD(162)(6) <= CNStageIntLLROutputS6xD(369)(2);
  VNStageIntLLRInputS6xD(214)(6) <= CNStageIntLLROutputS6xD(369)(3);
  VNStageIntLLRInputS6xD(310)(5) <= CNStageIntLLROutputS6xD(369)(4);
  VNStageIntLLRInputS6xD(324)(6) <= CNStageIntLLROutputS6xD(369)(5);
  VNStageIntLLRInputS6xD(50)(6) <= CNStageIntLLROutputS6xD(370)(0);
  VNStageIntLLRInputS6xD(97)(6) <= CNStageIntLLROutputS6xD(370)(1);
  VNStageIntLLRInputS6xD(149)(6) <= CNStageIntLLROutputS6xD(370)(2);
  VNStageIntLLRInputS6xD(245)(6) <= CNStageIntLLROutputS6xD(370)(3);
  VNStageIntLLRInputS6xD(259)(4) <= CNStageIntLLROutputS6xD(370)(4);
  VNStageIntLLRInputS6xD(338)(4) <= CNStageIntLLROutputS6xD(370)(5);
  VNStageIntLLRInputS6xD(49)(6) <= CNStageIntLLROutputS6xD(371)(0);
  VNStageIntLLRInputS6xD(84)(5) <= CNStageIntLLROutputS6xD(371)(1);
  VNStageIntLLRInputS6xD(180)(4) <= CNStageIntLLROutputS6xD(371)(2);
  VNStageIntLLRInputS6xD(194)(6) <= CNStageIntLLROutputS6xD(371)(3);
  VNStageIntLLRInputS6xD(273)(5) <= CNStageIntLLROutputS6xD(371)(4);
  VNStageIntLLRInputS6xD(382)(5) <= CNStageIntLLROutputS6xD(371)(5);
  VNStageIntLLRInputS6xD(48)(3) <= CNStageIntLLROutputS6xD(372)(0);
  VNStageIntLLRInputS6xD(115)(6) <= CNStageIntLLROutputS6xD(372)(1);
  VNStageIntLLRInputS6xD(129)(6) <= CNStageIntLLROutputS6xD(372)(2);
  VNStageIntLLRInputS6xD(208)(5) <= CNStageIntLLROutputS6xD(372)(3);
  VNStageIntLLRInputS6xD(317)(3) <= CNStageIntLLROutputS6xD(372)(4);
  VNStageIntLLRInputS6xD(359)(6) <= CNStageIntLLROutputS6xD(372)(5);
  VNStageIntLLRInputS6xD(47)(3) <= CNStageIntLLROutputS6xD(373)(0);
  VNStageIntLLRInputS6xD(127)(6) <= CNStageIntLLROutputS6xD(373)(1);
  VNStageIntLLRInputS6xD(143)(6) <= CNStageIntLLROutputS6xD(373)(2);
  VNStageIntLLRInputS6xD(252)(5) <= CNStageIntLLROutputS6xD(373)(3);
  VNStageIntLLRInputS6xD(294)(6) <= CNStageIntLLROutputS6xD(373)(4);
  VNStageIntLLRInputS6xD(348)(6) <= CNStageIntLLROutputS6xD(373)(5);
  VNStageIntLLRInputS6xD(46)(6) <= CNStageIntLLROutputS6xD(374)(0);
  VNStageIntLLRInputS6xD(78)(6) <= CNStageIntLLROutputS6xD(374)(1);
  VNStageIntLLRInputS6xD(187)(5) <= CNStageIntLLROutputS6xD(374)(2);
  VNStageIntLLRInputS6xD(229)(4) <= CNStageIntLLROutputS6xD(374)(3);
  VNStageIntLLRInputS6xD(283)(6) <= CNStageIntLLROutputS6xD(374)(4);
  VNStageIntLLRInputS6xD(352)(6) <= CNStageIntLLROutputS6xD(374)(5);
  VNStageIntLLRInputS6xD(45)(6) <= CNStageIntLLROutputS6xD(375)(0);
  VNStageIntLLRInputS6xD(122)(5) <= CNStageIntLLROutputS6xD(375)(1);
  VNStageIntLLRInputS6xD(164)(5) <= CNStageIntLLROutputS6xD(375)(2);
  VNStageIntLLRInputS6xD(218)(6) <= CNStageIntLLROutputS6xD(375)(3);
  VNStageIntLLRInputS6xD(287)(6) <= CNStageIntLLROutputS6xD(375)(4);
  VNStageIntLLRInputS6xD(345)(5) <= CNStageIntLLROutputS6xD(375)(5);
  VNStageIntLLRInputS6xD(44)(6) <= CNStageIntLLROutputS6xD(376)(0);
  VNStageIntLLRInputS6xD(99)(6) <= CNStageIntLLROutputS6xD(376)(1);
  VNStageIntLLRInputS6xD(153)(6) <= CNStageIntLLROutputS6xD(376)(2);
  VNStageIntLLRInputS6xD(222)(3) <= CNStageIntLLROutputS6xD(376)(3);
  VNStageIntLLRInputS6xD(280)(6) <= CNStageIntLLROutputS6xD(376)(4);
  VNStageIntLLRInputS6xD(356)(5) <= CNStageIntLLROutputS6xD(376)(5);
  VNStageIntLLRInputS6xD(43)(5) <= CNStageIntLLROutputS6xD(377)(0);
  VNStageIntLLRInputS6xD(88)(6) <= CNStageIntLLROutputS6xD(377)(1);
  VNStageIntLLRInputS6xD(157)(5) <= CNStageIntLLROutputS6xD(377)(2);
  VNStageIntLLRInputS6xD(215)(6) <= CNStageIntLLROutputS6xD(377)(3);
  VNStageIntLLRInputS6xD(291)(5) <= CNStageIntLLROutputS6xD(377)(4);
  VNStageIntLLRInputS6xD(328)(4) <= CNStageIntLLROutputS6xD(377)(5);
  VNStageIntLLRInputS6xD(42)(6) <= CNStageIntLLROutputS6xD(378)(0);
  VNStageIntLLRInputS6xD(92)(6) <= CNStageIntLLROutputS6xD(378)(1);
  VNStageIntLLRInputS6xD(150)(5) <= CNStageIntLLROutputS6xD(378)(2);
  VNStageIntLLRInputS6xD(226)(2) <= CNStageIntLLROutputS6xD(378)(3);
  VNStageIntLLRInputS6xD(263)(6) <= CNStageIntLLROutputS6xD(378)(4);
  VNStageIntLLRInputS6xD(383)(6) <= CNStageIntLLROutputS6xD(378)(5);
  VNStageIntLLRInputS6xD(41)(6) <= CNStageIntLLROutputS6xD(379)(0);
  VNStageIntLLRInputS6xD(85)(5) <= CNStageIntLLROutputS6xD(379)(1);
  VNStageIntLLRInputS6xD(161)(6) <= CNStageIntLLROutputS6xD(379)(2);
  VNStageIntLLRInputS6xD(198)(6) <= CNStageIntLLROutputS6xD(379)(3);
  VNStageIntLLRInputS6xD(318)(3) <= CNStageIntLLROutputS6xD(379)(4);
  VNStageIntLLRInputS6xD(337)(6) <= CNStageIntLLROutputS6xD(379)(5);
  VNStageIntLLRInputS6xD(40)(4) <= CNStageIntLLROutputS6xD(380)(0);
  VNStageIntLLRInputS6xD(96)(5) <= CNStageIntLLROutputS6xD(380)(1);
  VNStageIntLLRInputS6xD(133)(4) <= CNStageIntLLROutputS6xD(380)(2);
  VNStageIntLLRInputS6xD(253)(5) <= CNStageIntLLROutputS6xD(380)(3);
  VNStageIntLLRInputS6xD(272)(6) <= CNStageIntLLROutputS6xD(380)(4);
  VNStageIntLLRInputS6xD(334)(4) <= CNStageIntLLROutputS6xD(380)(5);
  VNStageIntLLRInputS6xD(39)(6) <= CNStageIntLLROutputS6xD(381)(0);
  VNStageIntLLRInputS6xD(68)(5) <= CNStageIntLLROutputS6xD(381)(1);
  VNStageIntLLRInputS6xD(188)(4) <= CNStageIntLLROutputS6xD(381)(2);
  VNStageIntLLRInputS6xD(207)(5) <= CNStageIntLLROutputS6xD(381)(3);
  VNStageIntLLRInputS6xD(269)(5) <= CNStageIntLLROutputS6xD(381)(4);
  VNStageIntLLRInputS6xD(368)(2) <= CNStageIntLLROutputS6xD(381)(5);
  VNStageIntLLRInputS6xD(38)(6) <= CNStageIntLLROutputS6xD(382)(0);
  VNStageIntLLRInputS6xD(123)(4) <= CNStageIntLLROutputS6xD(382)(1);
  VNStageIntLLRInputS6xD(142)(4) <= CNStageIntLLROutputS6xD(382)(2);
  VNStageIntLLRInputS6xD(204)(6) <= CNStageIntLLROutputS6xD(382)(3);
  VNStageIntLLRInputS6xD(303)(6) <= CNStageIntLLROutputS6xD(382)(4);
  VNStageIntLLRInputS6xD(325)(6) <= CNStageIntLLROutputS6xD(382)(5);
  VNStageIntLLRInputS6xD(37)(6) <= CNStageIntLLROutputS6xD(383)(0);
  VNStageIntLLRInputS6xD(77)(4) <= CNStageIntLLROutputS6xD(383)(1);
  VNStageIntLLRInputS6xD(139)(6) <= CNStageIntLLROutputS6xD(383)(2);
  VNStageIntLLRInputS6xD(238)(6) <= CNStageIntLLROutputS6xD(383)(3);
  VNStageIntLLRInputS6xD(260)(5) <= CNStageIntLLROutputS6xD(383)(4);
  VNStageIntLLRInputS6xD(374)(6) <= CNStageIntLLROutputS6xD(383)(5);

  -- Check Nodes (Iteration 7)
  CNStageIntLLRInputS7xD(53)(0) <= VNStageIntLLROutputS6xD(0)(0);
  CNStageIntLLRInputS7xD(110)(0) <= VNStageIntLLROutputS6xD(0)(1);
  CNStageIntLLRInputS7xD(170)(0) <= VNStageIntLLROutputS6xD(0)(2);
  CNStageIntLLRInputS7xD(224)(0) <= VNStageIntLLROutputS6xD(0)(3);
  CNStageIntLLRInputS7xD(279)(0) <= VNStageIntLLROutputS6xD(0)(4);
  CNStageIntLLRInputS7xD(332)(0) <= VNStageIntLLROutputS6xD(0)(5);
  CNStageIntLLRInputS7xD(51)(0) <= VNStageIntLLROutputS6xD(1)(0);
  CNStageIntLLRInputS7xD(139)(0) <= VNStageIntLLROutputS6xD(1)(1);
  CNStageIntLLRInputS7xD(223)(0) <= VNStageIntLLROutputS6xD(1)(2);
  CNStageIntLLRInputS7xD(241)(0) <= VNStageIntLLROutputS6xD(1)(3);
  CNStageIntLLRInputS7xD(307)(0) <= VNStageIntLLROutputS6xD(1)(4);
  CNStageIntLLRInputS7xD(356)(0) <= VNStageIntLLROutputS6xD(1)(5);
  CNStageIntLLRInputS7xD(50)(0) <= VNStageIntLLROutputS6xD(2)(0);
  CNStageIntLLRInputS7xD(92)(0) <= VNStageIntLLROutputS6xD(2)(1);
  CNStageIntLLRInputS7xD(138)(0) <= VNStageIntLLROutputS6xD(2)(2);
  CNStageIntLLRInputS7xD(222)(0) <= VNStageIntLLROutputS6xD(2)(3);
  CNStageIntLLRInputS7xD(240)(0) <= VNStageIntLLROutputS6xD(2)(4);
  CNStageIntLLRInputS7xD(306)(0) <= VNStageIntLLROutputS6xD(2)(5);
  CNStageIntLLRInputS7xD(355)(0) <= VNStageIntLLROutputS6xD(2)(6);
  CNStageIntLLRInputS7xD(91)(0) <= VNStageIntLLROutputS6xD(3)(0);
  CNStageIntLLRInputS7xD(137)(0) <= VNStageIntLLROutputS6xD(3)(1);
  CNStageIntLLRInputS7xD(221)(0) <= VNStageIntLLROutputS6xD(3)(2);
  CNStageIntLLRInputS7xD(239)(0) <= VNStageIntLLROutputS6xD(3)(3);
  CNStageIntLLRInputS7xD(305)(0) <= VNStageIntLLROutputS6xD(3)(4);
  CNStageIntLLRInputS7xD(49)(0) <= VNStageIntLLROutputS6xD(4)(0);
  CNStageIntLLRInputS7xD(90)(0) <= VNStageIntLLROutputS6xD(4)(1);
  CNStageIntLLRInputS7xD(220)(0) <= VNStageIntLLROutputS6xD(4)(2);
  CNStageIntLLRInputS7xD(238)(0) <= VNStageIntLLROutputS6xD(4)(3);
  CNStageIntLLRInputS7xD(304)(0) <= VNStageIntLLROutputS6xD(4)(4);
  CNStageIntLLRInputS7xD(354)(0) <= VNStageIntLLROutputS6xD(4)(5);
  CNStageIntLLRInputS7xD(48)(0) <= VNStageIntLLROutputS6xD(5)(0);
  CNStageIntLLRInputS7xD(89)(0) <= VNStageIntLLROutputS6xD(5)(1);
  CNStageIntLLRInputS7xD(136)(0) <= VNStageIntLLROutputS6xD(5)(2);
  CNStageIntLLRInputS7xD(219)(0) <= VNStageIntLLROutputS6xD(5)(3);
  CNStageIntLLRInputS7xD(237)(0) <= VNStageIntLLROutputS6xD(5)(4);
  CNStageIntLLRInputS7xD(303)(0) <= VNStageIntLLROutputS6xD(5)(5);
  CNStageIntLLRInputS7xD(353)(0) <= VNStageIntLLROutputS6xD(5)(6);
  CNStageIntLLRInputS7xD(47)(0) <= VNStageIntLLROutputS6xD(6)(0);
  CNStageIntLLRInputS7xD(88)(0) <= VNStageIntLLROutputS6xD(6)(1);
  CNStageIntLLRInputS7xD(135)(0) <= VNStageIntLLROutputS6xD(6)(2);
  CNStageIntLLRInputS7xD(218)(0) <= VNStageIntLLROutputS6xD(6)(3);
  CNStageIntLLRInputS7xD(236)(0) <= VNStageIntLLROutputS6xD(6)(4);
  CNStageIntLLRInputS7xD(302)(0) <= VNStageIntLLROutputS6xD(6)(5);
  CNStageIntLLRInputS7xD(352)(0) <= VNStageIntLLROutputS6xD(6)(6);
  CNStageIntLLRInputS7xD(46)(0) <= VNStageIntLLROutputS6xD(7)(0);
  CNStageIntLLRInputS7xD(87)(0) <= VNStageIntLLROutputS6xD(7)(1);
  CNStageIntLLRInputS7xD(134)(0) <= VNStageIntLLROutputS6xD(7)(2);
  CNStageIntLLRInputS7xD(217)(0) <= VNStageIntLLROutputS6xD(7)(3);
  CNStageIntLLRInputS7xD(235)(0) <= VNStageIntLLROutputS6xD(7)(4);
  CNStageIntLLRInputS7xD(301)(0) <= VNStageIntLLROutputS6xD(7)(5);
  CNStageIntLLRInputS7xD(351)(0) <= VNStageIntLLROutputS6xD(7)(6);
  CNStageIntLLRInputS7xD(45)(0) <= VNStageIntLLROutputS6xD(8)(0);
  CNStageIntLLRInputS7xD(133)(0) <= VNStageIntLLROutputS6xD(8)(1);
  CNStageIntLLRInputS7xD(216)(0) <= VNStageIntLLROutputS6xD(8)(2);
  CNStageIntLLRInputS7xD(44)(0) <= VNStageIntLLROutputS6xD(9)(0);
  CNStageIntLLRInputS7xD(86)(0) <= VNStageIntLLROutputS6xD(9)(1);
  CNStageIntLLRInputS7xD(132)(0) <= VNStageIntLLROutputS6xD(9)(2);
  CNStageIntLLRInputS7xD(215)(0) <= VNStageIntLLROutputS6xD(9)(3);
  CNStageIntLLRInputS7xD(234)(0) <= VNStageIntLLROutputS6xD(9)(4);
  CNStageIntLLRInputS7xD(300)(0) <= VNStageIntLLROutputS6xD(9)(5);
  CNStageIntLLRInputS7xD(350)(0) <= VNStageIntLLROutputS6xD(9)(6);
  CNStageIntLLRInputS7xD(43)(0) <= VNStageIntLLROutputS6xD(10)(0);
  CNStageIntLLRInputS7xD(85)(0) <= VNStageIntLLROutputS6xD(10)(1);
  CNStageIntLLRInputS7xD(131)(0) <= VNStageIntLLROutputS6xD(10)(2);
  CNStageIntLLRInputS7xD(233)(0) <= VNStageIntLLROutputS6xD(10)(3);
  CNStageIntLLRInputS7xD(349)(0) <= VNStageIntLLROutputS6xD(10)(4);
  CNStageIntLLRInputS7xD(42)(0) <= VNStageIntLLROutputS6xD(11)(0);
  CNStageIntLLRInputS7xD(84)(0) <= VNStageIntLLROutputS6xD(11)(1);
  CNStageIntLLRInputS7xD(130)(0) <= VNStageIntLLROutputS6xD(11)(2);
  CNStageIntLLRInputS7xD(214)(0) <= VNStageIntLLROutputS6xD(11)(3);
  CNStageIntLLRInputS7xD(232)(0) <= VNStageIntLLROutputS6xD(11)(4);
  CNStageIntLLRInputS7xD(348)(0) <= VNStageIntLLROutputS6xD(11)(5);
  CNStageIntLLRInputS7xD(41)(0) <= VNStageIntLLROutputS6xD(12)(0);
  CNStageIntLLRInputS7xD(83)(0) <= VNStageIntLLROutputS6xD(12)(1);
  CNStageIntLLRInputS7xD(129)(0) <= VNStageIntLLROutputS6xD(12)(2);
  CNStageIntLLRInputS7xD(213)(0) <= VNStageIntLLROutputS6xD(12)(3);
  CNStageIntLLRInputS7xD(231)(0) <= VNStageIntLLROutputS6xD(12)(4);
  CNStageIntLLRInputS7xD(299)(0) <= VNStageIntLLROutputS6xD(12)(5);
  CNStageIntLLRInputS7xD(347)(0) <= VNStageIntLLROutputS6xD(12)(6);
  CNStageIntLLRInputS7xD(82)(0) <= VNStageIntLLROutputS6xD(13)(0);
  CNStageIntLLRInputS7xD(128)(0) <= VNStageIntLLROutputS6xD(13)(1);
  CNStageIntLLRInputS7xD(212)(0) <= VNStageIntLLROutputS6xD(13)(2);
  CNStageIntLLRInputS7xD(230)(0) <= VNStageIntLLROutputS6xD(13)(3);
  CNStageIntLLRInputS7xD(298)(0) <= VNStageIntLLROutputS6xD(13)(4);
  CNStageIntLLRInputS7xD(346)(0) <= VNStageIntLLROutputS6xD(13)(5);
  CNStageIntLLRInputS7xD(40)(0) <= VNStageIntLLROutputS6xD(14)(0);
  CNStageIntLLRInputS7xD(81)(0) <= VNStageIntLLROutputS6xD(14)(1);
  CNStageIntLLRInputS7xD(127)(0) <= VNStageIntLLROutputS6xD(14)(2);
  CNStageIntLLRInputS7xD(211)(0) <= VNStageIntLLROutputS6xD(14)(3);
  CNStageIntLLRInputS7xD(229)(0) <= VNStageIntLLROutputS6xD(14)(4);
  CNStageIntLLRInputS7xD(297)(0) <= VNStageIntLLROutputS6xD(14)(5);
  CNStageIntLLRInputS7xD(345)(0) <= VNStageIntLLROutputS6xD(14)(6);
  CNStageIntLLRInputS7xD(39)(0) <= VNStageIntLLROutputS6xD(15)(0);
  CNStageIntLLRInputS7xD(80)(0) <= VNStageIntLLROutputS6xD(15)(1);
  CNStageIntLLRInputS7xD(126)(0) <= VNStageIntLLROutputS6xD(15)(2);
  CNStageIntLLRInputS7xD(210)(0) <= VNStageIntLLROutputS6xD(15)(3);
  CNStageIntLLRInputS7xD(228)(0) <= VNStageIntLLROutputS6xD(15)(4);
  CNStageIntLLRInputS7xD(296)(0) <= VNStageIntLLROutputS6xD(15)(5);
  CNStageIntLLRInputS7xD(344)(0) <= VNStageIntLLROutputS6xD(15)(6);
  CNStageIntLLRInputS7xD(38)(0) <= VNStageIntLLROutputS6xD(16)(0);
  CNStageIntLLRInputS7xD(125)(0) <= VNStageIntLLROutputS6xD(16)(1);
  CNStageIntLLRInputS7xD(209)(0) <= VNStageIntLLROutputS6xD(16)(2);
  CNStageIntLLRInputS7xD(227)(0) <= VNStageIntLLROutputS6xD(16)(3);
  CNStageIntLLRInputS7xD(295)(0) <= VNStageIntLLROutputS6xD(16)(4);
  CNStageIntLLRInputS7xD(343)(0) <= VNStageIntLLROutputS6xD(16)(5);
  CNStageIntLLRInputS7xD(37)(0) <= VNStageIntLLROutputS6xD(17)(0);
  CNStageIntLLRInputS7xD(79)(0) <= VNStageIntLLROutputS6xD(17)(1);
  CNStageIntLLRInputS7xD(124)(0) <= VNStageIntLLROutputS6xD(17)(2);
  CNStageIntLLRInputS7xD(208)(0) <= VNStageIntLLROutputS6xD(17)(3);
  CNStageIntLLRInputS7xD(226)(0) <= VNStageIntLLROutputS6xD(17)(4);
  CNStageIntLLRInputS7xD(294)(0) <= VNStageIntLLROutputS6xD(17)(5);
  CNStageIntLLRInputS7xD(342)(0) <= VNStageIntLLROutputS6xD(17)(6);
  CNStageIntLLRInputS7xD(36)(0) <= VNStageIntLLROutputS6xD(18)(0);
  CNStageIntLLRInputS7xD(78)(0) <= VNStageIntLLROutputS6xD(18)(1);
  CNStageIntLLRInputS7xD(123)(0) <= VNStageIntLLROutputS6xD(18)(2);
  CNStageIntLLRInputS7xD(207)(0) <= VNStageIntLLROutputS6xD(18)(3);
  CNStageIntLLRInputS7xD(225)(0) <= VNStageIntLLROutputS6xD(18)(4);
  CNStageIntLLRInputS7xD(293)(0) <= VNStageIntLLROutputS6xD(18)(5);
  CNStageIntLLRInputS7xD(341)(0) <= VNStageIntLLROutputS6xD(18)(6);
  CNStageIntLLRInputS7xD(35)(0) <= VNStageIntLLROutputS6xD(19)(0);
  CNStageIntLLRInputS7xD(77)(0) <= VNStageIntLLROutputS6xD(19)(1);
  CNStageIntLLRInputS7xD(122)(0) <= VNStageIntLLROutputS6xD(19)(2);
  CNStageIntLLRInputS7xD(278)(0) <= VNStageIntLLROutputS6xD(19)(3);
  CNStageIntLLRInputS7xD(340)(0) <= VNStageIntLLROutputS6xD(19)(4);
  CNStageIntLLRInputS7xD(34)(0) <= VNStageIntLLROutputS6xD(20)(0);
  CNStageIntLLRInputS7xD(76)(0) <= VNStageIntLLROutputS6xD(20)(1);
  CNStageIntLLRInputS7xD(277)(0) <= VNStageIntLLROutputS6xD(20)(2);
  CNStageIntLLRInputS7xD(292)(0) <= VNStageIntLLROutputS6xD(20)(3);
  CNStageIntLLRInputS7xD(339)(0) <= VNStageIntLLROutputS6xD(20)(4);
  CNStageIntLLRInputS7xD(33)(0) <= VNStageIntLLROutputS6xD(21)(0);
  CNStageIntLLRInputS7xD(75)(0) <= VNStageIntLLROutputS6xD(21)(1);
  CNStageIntLLRInputS7xD(121)(0) <= VNStageIntLLROutputS6xD(21)(2);
  CNStageIntLLRInputS7xD(206)(0) <= VNStageIntLLROutputS6xD(21)(3);
  CNStageIntLLRInputS7xD(276)(0) <= VNStageIntLLROutputS6xD(21)(4);
  CNStageIntLLRInputS7xD(291)(0) <= VNStageIntLLROutputS6xD(21)(5);
  CNStageIntLLRInputS7xD(338)(0) <= VNStageIntLLROutputS6xD(21)(6);
  CNStageIntLLRInputS7xD(32)(0) <= VNStageIntLLROutputS6xD(22)(0);
  CNStageIntLLRInputS7xD(74)(0) <= VNStageIntLLROutputS6xD(22)(1);
  CNStageIntLLRInputS7xD(120)(0) <= VNStageIntLLROutputS6xD(22)(2);
  CNStageIntLLRInputS7xD(205)(0) <= VNStageIntLLROutputS6xD(22)(3);
  CNStageIntLLRInputS7xD(275)(0) <= VNStageIntLLROutputS6xD(22)(4);
  CNStageIntLLRInputS7xD(290)(0) <= VNStageIntLLROutputS6xD(22)(5);
  CNStageIntLLRInputS7xD(337)(0) <= VNStageIntLLROutputS6xD(22)(6);
  CNStageIntLLRInputS7xD(31)(0) <= VNStageIntLLROutputS6xD(23)(0);
  CNStageIntLLRInputS7xD(73)(0) <= VNStageIntLLROutputS6xD(23)(1);
  CNStageIntLLRInputS7xD(119)(0) <= VNStageIntLLROutputS6xD(23)(2);
  CNStageIntLLRInputS7xD(204)(0) <= VNStageIntLLROutputS6xD(23)(3);
  CNStageIntLLRInputS7xD(274)(0) <= VNStageIntLLROutputS6xD(23)(4);
  CNStageIntLLRInputS7xD(289)(0) <= VNStageIntLLROutputS6xD(23)(5);
  CNStageIntLLRInputS7xD(336)(0) <= VNStageIntLLROutputS6xD(23)(6);
  CNStageIntLLRInputS7xD(30)(0) <= VNStageIntLLROutputS6xD(24)(0);
  CNStageIntLLRInputS7xD(72)(0) <= VNStageIntLLROutputS6xD(24)(1);
  CNStageIntLLRInputS7xD(118)(0) <= VNStageIntLLROutputS6xD(24)(2);
  CNStageIntLLRInputS7xD(203)(0) <= VNStageIntLLROutputS6xD(24)(3);
  CNStageIntLLRInputS7xD(273)(0) <= VNStageIntLLROutputS6xD(24)(4);
  CNStageIntLLRInputS7xD(288)(0) <= VNStageIntLLROutputS6xD(24)(5);
  CNStageIntLLRInputS7xD(335)(0) <= VNStageIntLLROutputS6xD(24)(6);
  CNStageIntLLRInputS7xD(29)(0) <= VNStageIntLLROutputS6xD(25)(0);
  CNStageIntLLRInputS7xD(71)(0) <= VNStageIntLLROutputS6xD(25)(1);
  CNStageIntLLRInputS7xD(117)(0) <= VNStageIntLLROutputS6xD(25)(2);
  CNStageIntLLRInputS7xD(202)(0) <= VNStageIntLLROutputS6xD(25)(3);
  CNStageIntLLRInputS7xD(287)(0) <= VNStageIntLLROutputS6xD(25)(4);
  CNStageIntLLRInputS7xD(28)(0) <= VNStageIntLLROutputS6xD(26)(0);
  CNStageIntLLRInputS7xD(70)(0) <= VNStageIntLLROutputS6xD(26)(1);
  CNStageIntLLRInputS7xD(116)(0) <= VNStageIntLLROutputS6xD(26)(2);
  CNStageIntLLRInputS7xD(201)(0) <= VNStageIntLLROutputS6xD(26)(3);
  CNStageIntLLRInputS7xD(272)(0) <= VNStageIntLLROutputS6xD(26)(4);
  CNStageIntLLRInputS7xD(286)(0) <= VNStageIntLLROutputS6xD(26)(5);
  CNStageIntLLRInputS7xD(334)(0) <= VNStageIntLLROutputS6xD(26)(6);
  CNStageIntLLRInputS7xD(27)(0) <= VNStageIntLLROutputS6xD(27)(0);
  CNStageIntLLRInputS7xD(69)(0) <= VNStageIntLLROutputS6xD(27)(1);
  CNStageIntLLRInputS7xD(115)(0) <= VNStageIntLLROutputS6xD(27)(2);
  CNStageIntLLRInputS7xD(200)(0) <= VNStageIntLLROutputS6xD(27)(3);
  CNStageIntLLRInputS7xD(285)(0) <= VNStageIntLLROutputS6xD(27)(4);
  CNStageIntLLRInputS7xD(26)(0) <= VNStageIntLLROutputS6xD(28)(0);
  CNStageIntLLRInputS7xD(68)(0) <= VNStageIntLLROutputS6xD(28)(1);
  CNStageIntLLRInputS7xD(114)(0) <= VNStageIntLLROutputS6xD(28)(2);
  CNStageIntLLRInputS7xD(199)(0) <= VNStageIntLLROutputS6xD(28)(3);
  CNStageIntLLRInputS7xD(271)(0) <= VNStageIntLLROutputS6xD(28)(4);
  CNStageIntLLRInputS7xD(333)(0) <= VNStageIntLLROutputS6xD(28)(5);
  CNStageIntLLRInputS7xD(25)(0) <= VNStageIntLLROutputS6xD(29)(0);
  CNStageIntLLRInputS7xD(67)(0) <= VNStageIntLLROutputS6xD(29)(1);
  CNStageIntLLRInputS7xD(113)(0) <= VNStageIntLLROutputS6xD(29)(2);
  CNStageIntLLRInputS7xD(270)(0) <= VNStageIntLLROutputS6xD(29)(3);
  CNStageIntLLRInputS7xD(24)(0) <= VNStageIntLLROutputS6xD(30)(0);
  CNStageIntLLRInputS7xD(66)(0) <= VNStageIntLLROutputS6xD(30)(1);
  CNStageIntLLRInputS7xD(112)(0) <= VNStageIntLLROutputS6xD(30)(2);
  CNStageIntLLRInputS7xD(198)(0) <= VNStageIntLLROutputS6xD(30)(3);
  CNStageIntLLRInputS7xD(269)(0) <= VNStageIntLLROutputS6xD(30)(4);
  CNStageIntLLRInputS7xD(284)(0) <= VNStageIntLLROutputS6xD(30)(5);
  CNStageIntLLRInputS7xD(23)(0) <= VNStageIntLLROutputS6xD(31)(0);
  CNStageIntLLRInputS7xD(65)(0) <= VNStageIntLLROutputS6xD(31)(1);
  CNStageIntLLRInputS7xD(197)(0) <= VNStageIntLLROutputS6xD(31)(2);
  CNStageIntLLRInputS7xD(283)(0) <= VNStageIntLLROutputS6xD(31)(3);
  CNStageIntLLRInputS7xD(22)(0) <= VNStageIntLLROutputS6xD(32)(0);
  CNStageIntLLRInputS7xD(64)(0) <= VNStageIntLLROutputS6xD(32)(1);
  CNStageIntLLRInputS7xD(111)(0) <= VNStageIntLLROutputS6xD(32)(2);
  CNStageIntLLRInputS7xD(268)(0) <= VNStageIntLLROutputS6xD(32)(3);
  CNStageIntLLRInputS7xD(21)(0) <= VNStageIntLLROutputS6xD(33)(0);
  CNStageIntLLRInputS7xD(63)(0) <= VNStageIntLLROutputS6xD(33)(1);
  CNStageIntLLRInputS7xD(169)(0) <= VNStageIntLLROutputS6xD(33)(2);
  CNStageIntLLRInputS7xD(196)(0) <= VNStageIntLLROutputS6xD(33)(3);
  CNStageIntLLRInputS7xD(267)(0) <= VNStageIntLLROutputS6xD(33)(4);
  CNStageIntLLRInputS7xD(282)(0) <= VNStageIntLLROutputS6xD(33)(5);
  CNStageIntLLRInputS7xD(20)(0) <= VNStageIntLLROutputS6xD(34)(0);
  CNStageIntLLRInputS7xD(62)(0) <= VNStageIntLLROutputS6xD(34)(1);
  CNStageIntLLRInputS7xD(168)(0) <= VNStageIntLLROutputS6xD(34)(2);
  CNStageIntLLRInputS7xD(195)(0) <= VNStageIntLLROutputS6xD(34)(3);
  CNStageIntLLRInputS7xD(266)(0) <= VNStageIntLLROutputS6xD(34)(4);
  CNStageIntLLRInputS7xD(281)(0) <= VNStageIntLLROutputS6xD(34)(5);
  CNStageIntLLRInputS7xD(19)(0) <= VNStageIntLLROutputS6xD(35)(0);
  CNStageIntLLRInputS7xD(61)(0) <= VNStageIntLLROutputS6xD(35)(1);
  CNStageIntLLRInputS7xD(167)(0) <= VNStageIntLLROutputS6xD(35)(2);
  CNStageIntLLRInputS7xD(194)(0) <= VNStageIntLLROutputS6xD(35)(3);
  CNStageIntLLRInputS7xD(265)(0) <= VNStageIntLLROutputS6xD(35)(4);
  CNStageIntLLRInputS7xD(280)(0) <= VNStageIntLLROutputS6xD(35)(5);
  CNStageIntLLRInputS7xD(18)(0) <= VNStageIntLLROutputS6xD(36)(0);
  CNStageIntLLRInputS7xD(60)(0) <= VNStageIntLLROutputS6xD(36)(1);
  CNStageIntLLRInputS7xD(166)(0) <= VNStageIntLLROutputS6xD(36)(2);
  CNStageIntLLRInputS7xD(264)(0) <= VNStageIntLLROutputS6xD(36)(3);
  CNStageIntLLRInputS7xD(17)(0) <= VNStageIntLLROutputS6xD(37)(0);
  CNStageIntLLRInputS7xD(59)(0) <= VNStageIntLLROutputS6xD(37)(1);
  CNStageIntLLRInputS7xD(165)(0) <= VNStageIntLLROutputS6xD(37)(2);
  CNStageIntLLRInputS7xD(193)(0) <= VNStageIntLLROutputS6xD(37)(3);
  CNStageIntLLRInputS7xD(263)(0) <= VNStageIntLLROutputS6xD(37)(4);
  CNStageIntLLRInputS7xD(331)(0) <= VNStageIntLLROutputS6xD(37)(5);
  CNStageIntLLRInputS7xD(383)(0) <= VNStageIntLLROutputS6xD(37)(6);
  CNStageIntLLRInputS7xD(16)(0) <= VNStageIntLLROutputS6xD(38)(0);
  CNStageIntLLRInputS7xD(58)(0) <= VNStageIntLLROutputS6xD(38)(1);
  CNStageIntLLRInputS7xD(164)(0) <= VNStageIntLLROutputS6xD(38)(2);
  CNStageIntLLRInputS7xD(192)(0) <= VNStageIntLLROutputS6xD(38)(3);
  CNStageIntLLRInputS7xD(262)(0) <= VNStageIntLLROutputS6xD(38)(4);
  CNStageIntLLRInputS7xD(330)(0) <= VNStageIntLLROutputS6xD(38)(5);
  CNStageIntLLRInputS7xD(382)(0) <= VNStageIntLLROutputS6xD(38)(6);
  CNStageIntLLRInputS7xD(15)(0) <= VNStageIntLLROutputS6xD(39)(0);
  CNStageIntLLRInputS7xD(57)(0) <= VNStageIntLLROutputS6xD(39)(1);
  CNStageIntLLRInputS7xD(163)(0) <= VNStageIntLLROutputS6xD(39)(2);
  CNStageIntLLRInputS7xD(191)(0) <= VNStageIntLLROutputS6xD(39)(3);
  CNStageIntLLRInputS7xD(261)(0) <= VNStageIntLLROutputS6xD(39)(4);
  CNStageIntLLRInputS7xD(329)(0) <= VNStageIntLLROutputS6xD(39)(5);
  CNStageIntLLRInputS7xD(381)(0) <= VNStageIntLLROutputS6xD(39)(6);
  CNStageIntLLRInputS7xD(14)(0) <= VNStageIntLLROutputS6xD(40)(0);
  CNStageIntLLRInputS7xD(56)(0) <= VNStageIntLLROutputS6xD(40)(1);
  CNStageIntLLRInputS7xD(162)(0) <= VNStageIntLLROutputS6xD(40)(2);
  CNStageIntLLRInputS7xD(260)(0) <= VNStageIntLLROutputS6xD(40)(3);
  CNStageIntLLRInputS7xD(380)(0) <= VNStageIntLLROutputS6xD(40)(4);
  CNStageIntLLRInputS7xD(13)(0) <= VNStageIntLLROutputS6xD(41)(0);
  CNStageIntLLRInputS7xD(55)(0) <= VNStageIntLLROutputS6xD(41)(1);
  CNStageIntLLRInputS7xD(161)(0) <= VNStageIntLLROutputS6xD(41)(2);
  CNStageIntLLRInputS7xD(190)(0) <= VNStageIntLLROutputS6xD(41)(3);
  CNStageIntLLRInputS7xD(259)(0) <= VNStageIntLLROutputS6xD(41)(4);
  CNStageIntLLRInputS7xD(328)(0) <= VNStageIntLLROutputS6xD(41)(5);
  CNStageIntLLRInputS7xD(379)(0) <= VNStageIntLLROutputS6xD(41)(6);
  CNStageIntLLRInputS7xD(12)(0) <= VNStageIntLLROutputS6xD(42)(0);
  CNStageIntLLRInputS7xD(54)(0) <= VNStageIntLLROutputS6xD(42)(1);
  CNStageIntLLRInputS7xD(160)(0) <= VNStageIntLLROutputS6xD(42)(2);
  CNStageIntLLRInputS7xD(189)(0) <= VNStageIntLLROutputS6xD(42)(3);
  CNStageIntLLRInputS7xD(258)(0) <= VNStageIntLLROutputS6xD(42)(4);
  CNStageIntLLRInputS7xD(327)(0) <= VNStageIntLLROutputS6xD(42)(5);
  CNStageIntLLRInputS7xD(378)(0) <= VNStageIntLLROutputS6xD(42)(6);
  CNStageIntLLRInputS7xD(109)(0) <= VNStageIntLLROutputS6xD(43)(0);
  CNStageIntLLRInputS7xD(159)(0) <= VNStageIntLLROutputS6xD(43)(1);
  CNStageIntLLRInputS7xD(188)(0) <= VNStageIntLLROutputS6xD(43)(2);
  CNStageIntLLRInputS7xD(257)(0) <= VNStageIntLLROutputS6xD(43)(3);
  CNStageIntLLRInputS7xD(326)(0) <= VNStageIntLLROutputS6xD(43)(4);
  CNStageIntLLRInputS7xD(377)(0) <= VNStageIntLLROutputS6xD(43)(5);
  CNStageIntLLRInputS7xD(11)(0) <= VNStageIntLLROutputS6xD(44)(0);
  CNStageIntLLRInputS7xD(108)(0) <= VNStageIntLLROutputS6xD(44)(1);
  CNStageIntLLRInputS7xD(158)(0) <= VNStageIntLLROutputS6xD(44)(2);
  CNStageIntLLRInputS7xD(187)(0) <= VNStageIntLLROutputS6xD(44)(3);
  CNStageIntLLRInputS7xD(256)(0) <= VNStageIntLLROutputS6xD(44)(4);
  CNStageIntLLRInputS7xD(325)(0) <= VNStageIntLLROutputS6xD(44)(5);
  CNStageIntLLRInputS7xD(376)(0) <= VNStageIntLLROutputS6xD(44)(6);
  CNStageIntLLRInputS7xD(10)(0) <= VNStageIntLLROutputS6xD(45)(0);
  CNStageIntLLRInputS7xD(107)(0) <= VNStageIntLLROutputS6xD(45)(1);
  CNStageIntLLRInputS7xD(157)(0) <= VNStageIntLLROutputS6xD(45)(2);
  CNStageIntLLRInputS7xD(186)(0) <= VNStageIntLLROutputS6xD(45)(3);
  CNStageIntLLRInputS7xD(255)(0) <= VNStageIntLLROutputS6xD(45)(4);
  CNStageIntLLRInputS7xD(324)(0) <= VNStageIntLLROutputS6xD(45)(5);
  CNStageIntLLRInputS7xD(375)(0) <= VNStageIntLLROutputS6xD(45)(6);
  CNStageIntLLRInputS7xD(9)(0) <= VNStageIntLLROutputS6xD(46)(0);
  CNStageIntLLRInputS7xD(106)(0) <= VNStageIntLLROutputS6xD(46)(1);
  CNStageIntLLRInputS7xD(156)(0) <= VNStageIntLLROutputS6xD(46)(2);
  CNStageIntLLRInputS7xD(185)(0) <= VNStageIntLLROutputS6xD(46)(3);
  CNStageIntLLRInputS7xD(254)(0) <= VNStageIntLLROutputS6xD(46)(4);
  CNStageIntLLRInputS7xD(323)(0) <= VNStageIntLLROutputS6xD(46)(5);
  CNStageIntLLRInputS7xD(374)(0) <= VNStageIntLLROutputS6xD(46)(6);
  CNStageIntLLRInputS7xD(8)(0) <= VNStageIntLLROutputS6xD(47)(0);
  CNStageIntLLRInputS7xD(155)(0) <= VNStageIntLLROutputS6xD(47)(1);
  CNStageIntLLRInputS7xD(253)(0) <= VNStageIntLLROutputS6xD(47)(2);
  CNStageIntLLRInputS7xD(373)(0) <= VNStageIntLLROutputS6xD(47)(3);
  CNStageIntLLRInputS7xD(7)(0) <= VNStageIntLLROutputS6xD(48)(0);
  CNStageIntLLRInputS7xD(154)(0) <= VNStageIntLLROutputS6xD(48)(1);
  CNStageIntLLRInputS7xD(322)(0) <= VNStageIntLLROutputS6xD(48)(2);
  CNStageIntLLRInputS7xD(372)(0) <= VNStageIntLLROutputS6xD(48)(3);
  CNStageIntLLRInputS7xD(6)(0) <= VNStageIntLLROutputS6xD(49)(0);
  CNStageIntLLRInputS7xD(105)(0) <= VNStageIntLLROutputS6xD(49)(1);
  CNStageIntLLRInputS7xD(153)(0) <= VNStageIntLLROutputS6xD(49)(2);
  CNStageIntLLRInputS7xD(184)(0) <= VNStageIntLLROutputS6xD(49)(3);
  CNStageIntLLRInputS7xD(252)(0) <= VNStageIntLLROutputS6xD(49)(4);
  CNStageIntLLRInputS7xD(321)(0) <= VNStageIntLLROutputS6xD(49)(5);
  CNStageIntLLRInputS7xD(371)(0) <= VNStageIntLLROutputS6xD(49)(6);
  CNStageIntLLRInputS7xD(5)(0) <= VNStageIntLLROutputS6xD(50)(0);
  CNStageIntLLRInputS7xD(104)(0) <= VNStageIntLLROutputS6xD(50)(1);
  CNStageIntLLRInputS7xD(152)(0) <= VNStageIntLLROutputS6xD(50)(2);
  CNStageIntLLRInputS7xD(183)(0) <= VNStageIntLLROutputS6xD(50)(3);
  CNStageIntLLRInputS7xD(251)(0) <= VNStageIntLLROutputS6xD(50)(4);
  CNStageIntLLRInputS7xD(320)(0) <= VNStageIntLLROutputS6xD(50)(5);
  CNStageIntLLRInputS7xD(370)(0) <= VNStageIntLLROutputS6xD(50)(6);
  CNStageIntLLRInputS7xD(4)(0) <= VNStageIntLLROutputS6xD(51)(0);
  CNStageIntLLRInputS7xD(103)(0) <= VNStageIntLLROutputS6xD(51)(1);
  CNStageIntLLRInputS7xD(182)(0) <= VNStageIntLLROutputS6xD(51)(2);
  CNStageIntLLRInputS7xD(250)(0) <= VNStageIntLLROutputS6xD(51)(3);
  CNStageIntLLRInputS7xD(319)(0) <= VNStageIntLLROutputS6xD(51)(4);
  CNStageIntLLRInputS7xD(369)(0) <= VNStageIntLLROutputS6xD(51)(5);
  CNStageIntLLRInputS7xD(102)(0) <= VNStageIntLLROutputS6xD(52)(0);
  CNStageIntLLRInputS7xD(151)(0) <= VNStageIntLLROutputS6xD(52)(1);
  CNStageIntLLRInputS7xD(181)(0) <= VNStageIntLLROutputS6xD(52)(2);
  CNStageIntLLRInputS7xD(318)(0) <= VNStageIntLLROutputS6xD(52)(3);
  CNStageIntLLRInputS7xD(368)(0) <= VNStageIntLLROutputS6xD(52)(4);
  CNStageIntLLRInputS7xD(3)(0) <= VNStageIntLLROutputS6xD(53)(0);
  CNStageIntLLRInputS7xD(150)(0) <= VNStageIntLLROutputS6xD(53)(1);
  CNStageIntLLRInputS7xD(180)(0) <= VNStageIntLLROutputS6xD(53)(2);
  CNStageIntLLRInputS7xD(249)(0) <= VNStageIntLLROutputS6xD(53)(3);
  CNStageIntLLRInputS7xD(317)(0) <= VNStageIntLLROutputS6xD(53)(4);
  CNStageIntLLRInputS7xD(367)(0) <= VNStageIntLLROutputS6xD(53)(5);
  CNStageIntLLRInputS7xD(2)(0) <= VNStageIntLLROutputS6xD(54)(0);
  CNStageIntLLRInputS7xD(101)(0) <= VNStageIntLLROutputS6xD(54)(1);
  CNStageIntLLRInputS7xD(149)(0) <= VNStageIntLLROutputS6xD(54)(2);
  CNStageIntLLRInputS7xD(179)(0) <= VNStageIntLLROutputS6xD(54)(3);
  CNStageIntLLRInputS7xD(316)(0) <= VNStageIntLLROutputS6xD(54)(4);
  CNStageIntLLRInputS7xD(366)(0) <= VNStageIntLLROutputS6xD(54)(5);
  CNStageIntLLRInputS7xD(1)(0) <= VNStageIntLLROutputS6xD(55)(0);
  CNStageIntLLRInputS7xD(100)(0) <= VNStageIntLLROutputS6xD(55)(1);
  CNStageIntLLRInputS7xD(148)(0) <= VNStageIntLLROutputS6xD(55)(2);
  CNStageIntLLRInputS7xD(178)(0) <= VNStageIntLLROutputS6xD(55)(3);
  CNStageIntLLRInputS7xD(248)(0) <= VNStageIntLLROutputS6xD(55)(4);
  CNStageIntLLRInputS7xD(315)(0) <= VNStageIntLLROutputS6xD(55)(5);
  CNStageIntLLRInputS7xD(365)(0) <= VNStageIntLLROutputS6xD(55)(6);
  CNStageIntLLRInputS7xD(0)(0) <= VNStageIntLLROutputS6xD(56)(0);
  CNStageIntLLRInputS7xD(99)(0) <= VNStageIntLLROutputS6xD(56)(1);
  CNStageIntLLRInputS7xD(147)(0) <= VNStageIntLLROutputS6xD(56)(2);
  CNStageIntLLRInputS7xD(177)(0) <= VNStageIntLLROutputS6xD(56)(3);
  CNStageIntLLRInputS7xD(247)(0) <= VNStageIntLLROutputS6xD(56)(4);
  CNStageIntLLRInputS7xD(314)(0) <= VNStageIntLLROutputS6xD(56)(5);
  CNStageIntLLRInputS7xD(364)(0) <= VNStageIntLLROutputS6xD(56)(6);
  CNStageIntLLRInputS7xD(98)(0) <= VNStageIntLLROutputS6xD(57)(0);
  CNStageIntLLRInputS7xD(146)(0) <= VNStageIntLLROutputS6xD(57)(1);
  CNStageIntLLRInputS7xD(176)(0) <= VNStageIntLLROutputS6xD(57)(2);
  CNStageIntLLRInputS7xD(246)(0) <= VNStageIntLLROutputS6xD(57)(3);
  CNStageIntLLRInputS7xD(313)(0) <= VNStageIntLLROutputS6xD(57)(4);
  CNStageIntLLRInputS7xD(363)(0) <= VNStageIntLLROutputS6xD(57)(5);
  CNStageIntLLRInputS7xD(97)(0) <= VNStageIntLLROutputS6xD(58)(0);
  CNStageIntLLRInputS7xD(145)(0) <= VNStageIntLLROutputS6xD(58)(1);
  CNStageIntLLRInputS7xD(175)(0) <= VNStageIntLLROutputS6xD(58)(2);
  CNStageIntLLRInputS7xD(312)(0) <= VNStageIntLLROutputS6xD(58)(3);
  CNStageIntLLRInputS7xD(362)(0) <= VNStageIntLLROutputS6xD(58)(4);
  CNStageIntLLRInputS7xD(144)(0) <= VNStageIntLLROutputS6xD(59)(0);
  CNStageIntLLRInputS7xD(174)(0) <= VNStageIntLLROutputS6xD(59)(1);
  CNStageIntLLRInputS7xD(245)(0) <= VNStageIntLLROutputS6xD(59)(2);
  CNStageIntLLRInputS7xD(311)(0) <= VNStageIntLLROutputS6xD(59)(3);
  CNStageIntLLRInputS7xD(361)(0) <= VNStageIntLLROutputS6xD(59)(4);
  CNStageIntLLRInputS7xD(96)(0) <= VNStageIntLLROutputS6xD(60)(0);
  CNStageIntLLRInputS7xD(143)(0) <= VNStageIntLLROutputS6xD(60)(1);
  CNStageIntLLRInputS7xD(173)(0) <= VNStageIntLLROutputS6xD(60)(2);
  CNStageIntLLRInputS7xD(244)(0) <= VNStageIntLLROutputS6xD(60)(3);
  CNStageIntLLRInputS7xD(310)(0) <= VNStageIntLLROutputS6xD(60)(4);
  CNStageIntLLRInputS7xD(360)(0) <= VNStageIntLLROutputS6xD(60)(5);
  CNStageIntLLRInputS7xD(95)(0) <= VNStageIntLLROutputS6xD(61)(0);
  CNStageIntLLRInputS7xD(142)(0) <= VNStageIntLLROutputS6xD(61)(1);
  CNStageIntLLRInputS7xD(172)(0) <= VNStageIntLLROutputS6xD(61)(2);
  CNStageIntLLRInputS7xD(243)(0) <= VNStageIntLLROutputS6xD(61)(3);
  CNStageIntLLRInputS7xD(309)(0) <= VNStageIntLLROutputS6xD(61)(4);
  CNStageIntLLRInputS7xD(359)(0) <= VNStageIntLLROutputS6xD(61)(5);
  CNStageIntLLRInputS7xD(94)(0) <= VNStageIntLLROutputS6xD(62)(0);
  CNStageIntLLRInputS7xD(141)(0) <= VNStageIntLLROutputS6xD(62)(1);
  CNStageIntLLRInputS7xD(171)(0) <= VNStageIntLLROutputS6xD(62)(2);
  CNStageIntLLRInputS7xD(242)(0) <= VNStageIntLLROutputS6xD(62)(3);
  CNStageIntLLRInputS7xD(308)(0) <= VNStageIntLLROutputS6xD(62)(4);
  CNStageIntLLRInputS7xD(358)(0) <= VNStageIntLLROutputS6xD(62)(5);
  CNStageIntLLRInputS7xD(52)(0) <= VNStageIntLLROutputS6xD(63)(0);
  CNStageIntLLRInputS7xD(93)(0) <= VNStageIntLLROutputS6xD(63)(1);
  CNStageIntLLRInputS7xD(140)(0) <= VNStageIntLLROutputS6xD(63)(2);
  CNStageIntLLRInputS7xD(357)(0) <= VNStageIntLLROutputS6xD(63)(3);
  CNStageIntLLRInputS7xD(53)(1) <= VNStageIntLLROutputS6xD(64)(0);
  CNStageIntLLRInputS7xD(109)(1) <= VNStageIntLLROutputS6xD(64)(1);
  CNStageIntLLRInputS7xD(130)(1) <= VNStageIntLLROutputS6xD(64)(2);
  CNStageIntLLRInputS7xD(245)(1) <= VNStageIntLLROutputS6xD(64)(3);
  CNStageIntLLRInputS7xD(299)(1) <= VNStageIntLLROutputS6xD(64)(4);
  CNStageIntLLRInputS7xD(342)(1) <= VNStageIntLLROutputS6xD(64)(5);
  CNStageIntLLRInputS7xD(51)(1) <= VNStageIntLLROutputS6xD(65)(0);
  CNStageIntLLRInputS7xD(74)(1) <= VNStageIntLLROutputS6xD(65)(1);
  CNStageIntLLRInputS7xD(141)(1) <= VNStageIntLLROutputS6xD(65)(2);
  CNStageIntLLRInputS7xD(189)(1) <= VNStageIntLLROutputS6xD(65)(3);
  CNStageIntLLRInputS7xD(286)(1) <= VNStageIntLLROutputS6xD(65)(4);
  CNStageIntLLRInputS7xD(50)(1) <= VNStageIntLLROutputS6xD(66)(0);
  CNStageIntLLRInputS7xD(66)(1) <= VNStageIntLLROutputS6xD(66)(1);
  CNStageIntLLRInputS7xD(155)(1) <= VNStageIntLLROutputS6xD(66)(2);
  CNStageIntLLRInputS7xD(244)(1) <= VNStageIntLLROutputS6xD(66)(3);
  CNStageIntLLRInputS7xD(97)(1) <= VNStageIntLLROutputS6xD(67)(0);
  CNStageIntLLRInputS7xD(275)(1) <= VNStageIntLLROutputS6xD(67)(1);
  CNStageIntLLRInputS7xD(322)(1) <= VNStageIntLLROutputS6xD(67)(2);
  CNStageIntLLRInputS7xD(365)(1) <= VNStageIntLLROutputS6xD(67)(3);
  CNStageIntLLRInputS7xD(49)(1) <= VNStageIntLLROutputS6xD(68)(0);
  CNStageIntLLRInputS7xD(112)(1) <= VNStageIntLLROutputS6xD(68)(1);
  CNStageIntLLRInputS7xD(210)(1) <= VNStageIntLLROutputS6xD(68)(2);
  CNStageIntLLRInputS7xD(256)(1) <= VNStageIntLLROutputS6xD(68)(3);
  CNStageIntLLRInputS7xD(318)(1) <= VNStageIntLLROutputS6xD(68)(4);
  CNStageIntLLRInputS7xD(381)(1) <= VNStageIntLLROutputS6xD(68)(5);
  CNStageIntLLRInputS7xD(48)(1) <= VNStageIntLLROutputS6xD(69)(0);
  CNStageIntLLRInputS7xD(101)(1) <= VNStageIntLLROutputS6xD(69)(1);
  CNStageIntLLRInputS7xD(135)(1) <= VNStageIntLLROutputS6xD(69)(2);
  CNStageIntLLRInputS7xD(215)(1) <= VNStageIntLLROutputS6xD(69)(3);
  CNStageIntLLRInputS7xD(259)(1) <= VNStageIntLLROutputS6xD(69)(4);
  CNStageIntLLRInputS7xD(283)(1) <= VNStageIntLLROutputS6xD(69)(5);
  CNStageIntLLRInputS7xD(351)(1) <= VNStageIntLLROutputS6xD(69)(6);
  CNStageIntLLRInputS7xD(47)(1) <= VNStageIntLLROutputS6xD(70)(0);
  CNStageIntLLRInputS7xD(104)(1) <= VNStageIntLLROutputS6xD(70)(1);
  CNStageIntLLRInputS7xD(136)(1) <= VNStageIntLLROutputS6xD(70)(2);
  CNStageIntLLRInputS7xD(206)(1) <= VNStageIntLLROutputS6xD(70)(3);
  CNStageIntLLRInputS7xD(246)(1) <= VNStageIntLLROutputS6xD(70)(4);
  CNStageIntLLRInputS7xD(301)(1) <= VNStageIntLLROutputS6xD(70)(5);
  CNStageIntLLRInputS7xD(46)(1) <= VNStageIntLLROutputS6xD(71)(0);
  CNStageIntLLRInputS7xD(95)(1) <= VNStageIntLLROutputS6xD(71)(1);
  CNStageIntLLRInputS7xD(176)(1) <= VNStageIntLLROutputS6xD(71)(2);
  CNStageIntLLRInputS7xD(276)(1) <= VNStageIntLLROutputS6xD(71)(3);
  CNStageIntLLRInputS7xD(302)(1) <= VNStageIntLLROutputS6xD(71)(4);
  CNStageIntLLRInputS7xD(353)(1) <= VNStageIntLLROutputS6xD(71)(5);
  CNStageIntLLRInputS7xD(45)(1) <= VNStageIntLLROutputS6xD(72)(0);
  CNStageIntLLRInputS7xD(75)(1) <= VNStageIntLLROutputS6xD(72)(1);
  CNStageIntLLRInputS7xD(162)(1) <= VNStageIntLLROutputS6xD(72)(2);
  CNStageIntLLRInputS7xD(183)(1) <= VNStageIntLLROutputS6xD(72)(3);
  CNStageIntLLRInputS7xD(243)(1) <= VNStageIntLLROutputS6xD(72)(4);
  CNStageIntLLRInputS7xD(367)(1) <= VNStageIntLLROutputS6xD(72)(5);
  CNStageIntLLRInputS7xD(44)(1) <= VNStageIntLLROutputS6xD(73)(0);
  CNStageIntLLRInputS7xD(56)(1) <= VNStageIntLLROutputS6xD(73)(1);
  CNStageIntLLRInputS7xD(121)(1) <= VNStageIntLLROutputS6xD(73)(2);
  CNStageIntLLRInputS7xD(219)(1) <= VNStageIntLLROutputS6xD(73)(3);
  CNStageIntLLRInputS7xD(328)(1) <= VNStageIntLLROutputS6xD(73)(4);
  CNStageIntLLRInputS7xD(363)(1) <= VNStageIntLLROutputS6xD(73)(5);
  CNStageIntLLRInputS7xD(43)(1) <= VNStageIntLLROutputS6xD(74)(0);
  CNStageIntLLRInputS7xD(70)(1) <= VNStageIntLLROutputS6xD(74)(1);
  CNStageIntLLRInputS7xD(125)(1) <= VNStageIntLLROutputS6xD(74)(2);
  CNStageIntLLRInputS7xD(221)(1) <= VNStageIntLLROutputS6xD(74)(3);
  CNStageIntLLRInputS7xD(290)(1) <= VNStageIntLLROutputS6xD(74)(4);
  CNStageIntLLRInputS7xD(42)(1) <= VNStageIntLLROutputS6xD(75)(0);
  CNStageIntLLRInputS7xD(81)(1) <= VNStageIntLLROutputS6xD(75)(1);
  CNStageIntLLRInputS7xD(170)(1) <= VNStageIntLLROutputS6xD(75)(2);
  CNStageIntLLRInputS7xD(192)(1) <= VNStageIntLLROutputS6xD(75)(3);
  CNStageIntLLRInputS7xD(278)(1) <= VNStageIntLLROutputS6xD(75)(4);
  CNStageIntLLRInputS7xD(294)(1) <= VNStageIntLLROutputS6xD(75)(5);
  CNStageIntLLRInputS7xD(347)(1) <= VNStageIntLLROutputS6xD(75)(6);
  CNStageIntLLRInputS7xD(41)(1) <= VNStageIntLLROutputS6xD(76)(0);
  CNStageIntLLRInputS7xD(106)(1) <= VNStageIntLLROutputS6xD(76)(1);
  CNStageIntLLRInputS7xD(124)(1) <= VNStageIntLLROutputS6xD(76)(2);
  CNStageIntLLRInputS7xD(174)(1) <= VNStageIntLLROutputS6xD(76)(3);
  CNStageIntLLRInputS7xD(270)(1) <= VNStageIntLLROutputS6xD(76)(4);
  CNStageIntLLRInputS7xD(332)(1) <= VNStageIntLLROutputS6xD(76)(5);
  CNStageIntLLRInputS7xD(348)(1) <= VNStageIntLLROutputS6xD(76)(6);
  CNStageIntLLRInputS7xD(119)(1) <= VNStageIntLLROutputS6xD(77)(0);
  CNStageIntLLRInputS7xD(185)(1) <= VNStageIntLLROutputS6xD(77)(1);
  CNStageIntLLRInputS7xD(257)(1) <= VNStageIntLLROutputS6xD(77)(2);
  CNStageIntLLRInputS7xD(293)(1) <= VNStageIntLLROutputS6xD(77)(3);
  CNStageIntLLRInputS7xD(383)(1) <= VNStageIntLLROutputS6xD(77)(4);
  CNStageIntLLRInputS7xD(40)(1) <= VNStageIntLLROutputS6xD(78)(0);
  CNStageIntLLRInputS7xD(84)(1) <= VNStageIntLLROutputS6xD(78)(1);
  CNStageIntLLRInputS7xD(159)(1) <= VNStageIntLLROutputS6xD(78)(2);
  CNStageIntLLRInputS7xD(193)(1) <= VNStageIntLLROutputS6xD(78)(3);
  CNStageIntLLRInputS7xD(274)(1) <= VNStageIntLLROutputS6xD(78)(4);
  CNStageIntLLRInputS7xD(288)(1) <= VNStageIntLLROutputS6xD(78)(5);
  CNStageIntLLRInputS7xD(374)(1) <= VNStageIntLLROutputS6xD(78)(6);
  CNStageIntLLRInputS7xD(39)(1) <= VNStageIntLLROutputS6xD(79)(0);
  CNStageIntLLRInputS7xD(99)(1) <= VNStageIntLLROutputS6xD(79)(1);
  CNStageIntLLRInputS7xD(167)(1) <= VNStageIntLLROutputS6xD(79)(2);
  CNStageIntLLRInputS7xD(220)(1) <= VNStageIntLLROutputS6xD(79)(3);
  CNStageIntLLRInputS7xD(325)(1) <= VNStageIntLLROutputS6xD(79)(4);
  CNStageIntLLRInputS7xD(38)(1) <= VNStageIntLLROutputS6xD(80)(0);
  CNStageIntLLRInputS7xD(62)(1) <= VNStageIntLLROutputS6xD(80)(1);
  CNStageIntLLRInputS7xD(131)(1) <= VNStageIntLLROutputS6xD(80)(2);
  CNStageIntLLRInputS7xD(182)(1) <= VNStageIntLLROutputS6xD(80)(3);
  CNStageIntLLRInputS7xD(248)(1) <= VNStageIntLLROutputS6xD(80)(4);
  CNStageIntLLRInputS7xD(337)(1) <= VNStageIntLLROutputS6xD(80)(5);
  CNStageIntLLRInputS7xD(37)(1) <= VNStageIntLLROutputS6xD(81)(0);
  CNStageIntLLRInputS7xD(72)(1) <= VNStageIntLLROutputS6xD(81)(1);
  CNStageIntLLRInputS7xD(129)(1) <= VNStageIntLLROutputS6xD(81)(2);
  CNStageIntLLRInputS7xD(262)(1) <= VNStageIntLLROutputS6xD(81)(3);
  CNStageIntLLRInputS7xD(36)(1) <= VNStageIntLLROutputS6xD(82)(0);
  CNStageIntLLRInputS7xD(67)(1) <= VNStageIntLLROutputS6xD(82)(1);
  CNStageIntLLRInputS7xD(165)(1) <= VNStageIntLLROutputS6xD(82)(2);
  CNStageIntLLRInputS7xD(188)(1) <= VNStageIntLLROutputS6xD(82)(3);
  CNStageIntLLRInputS7xD(254)(1) <= VNStageIntLLROutputS6xD(82)(4);
  CNStageIntLLRInputS7xD(298)(1) <= VNStageIntLLROutputS6xD(82)(5);
  CNStageIntLLRInputS7xD(336)(1) <= VNStageIntLLROutputS6xD(82)(6);
  CNStageIntLLRInputS7xD(35)(1) <= VNStageIntLLROutputS6xD(83)(0);
  CNStageIntLLRInputS7xD(73)(1) <= VNStageIntLLROutputS6xD(83)(1);
  CNStageIntLLRInputS7xD(144)(1) <= VNStageIntLLROutputS6xD(83)(2);
  CNStageIntLLRInputS7xD(208)(1) <= VNStageIntLLROutputS6xD(83)(3);
  CNStageIntLLRInputS7xD(232)(1) <= VNStageIntLLROutputS6xD(83)(4);
  CNStageIntLLRInputS7xD(330)(1) <= VNStageIntLLROutputS6xD(83)(5);
  CNStageIntLLRInputS7xD(34)(1) <= VNStageIntLLROutputS6xD(84)(0);
  CNStageIntLLRInputS7xD(61)(1) <= VNStageIntLLROutputS6xD(84)(1);
  CNStageIntLLRInputS7xD(147)(1) <= VNStageIntLLROutputS6xD(84)(2);
  CNStageIntLLRInputS7xD(222)(1) <= VNStageIntLLROutputS6xD(84)(3);
  CNStageIntLLRInputS7xD(310)(1) <= VNStageIntLLROutputS6xD(84)(4);
  CNStageIntLLRInputS7xD(371)(1) <= VNStageIntLLROutputS6xD(84)(5);
  CNStageIntLLRInputS7xD(33)(1) <= VNStageIntLLROutputS6xD(85)(0);
  CNStageIntLLRInputS7xD(132)(1) <= VNStageIntLLROutputS6xD(85)(1);
  CNStageIntLLRInputS7xD(218)(1) <= VNStageIntLLROutputS6xD(85)(2);
  CNStageIntLLRInputS7xD(235)(1) <= VNStageIntLLROutputS6xD(85)(3);
  CNStageIntLLRInputS7xD(313)(1) <= VNStageIntLLROutputS6xD(85)(4);
  CNStageIntLLRInputS7xD(379)(1) <= VNStageIntLLROutputS6xD(85)(5);
  CNStageIntLLRInputS7xD(32)(1) <= VNStageIntLLROutputS6xD(86)(0);
  CNStageIntLLRInputS7xD(166)(1) <= VNStageIntLLROutputS6xD(86)(1);
  CNStageIntLLRInputS7xD(239)(1) <= VNStageIntLLROutputS6xD(86)(2);
  CNStageIntLLRInputS7xD(343)(1) <= VNStageIntLLROutputS6xD(86)(3);
  CNStageIntLLRInputS7xD(31)(1) <= VNStageIntLLROutputS6xD(87)(0);
  CNStageIntLLRInputS7xD(77)(1) <= VNStageIntLLROutputS6xD(87)(1);
  CNStageIntLLRInputS7xD(128)(1) <= VNStageIntLLROutputS6xD(87)(2);
  CNStageIntLLRInputS7xD(203)(1) <= VNStageIntLLROutputS6xD(87)(3);
  CNStageIntLLRInputS7xD(229)(1) <= VNStageIntLLROutputS6xD(87)(4);
  CNStageIntLLRInputS7xD(331)(1) <= VNStageIntLLROutputS6xD(87)(5);
  CNStageIntLLRInputS7xD(341)(1) <= VNStageIntLLROutputS6xD(87)(6);
  CNStageIntLLRInputS7xD(30)(1) <= VNStageIntLLROutputS6xD(88)(0);
  CNStageIntLLRInputS7xD(79)(1) <= VNStageIntLLROutputS6xD(88)(1);
  CNStageIntLLRInputS7xD(156)(1) <= VNStageIntLLROutputS6xD(88)(2);
  CNStageIntLLRInputS7xD(204)(1) <= VNStageIntLLROutputS6xD(88)(3);
  CNStageIntLLRInputS7xD(263)(1) <= VNStageIntLLROutputS6xD(88)(4);
  CNStageIntLLRInputS7xD(297)(1) <= VNStageIntLLROutputS6xD(88)(5);
  CNStageIntLLRInputS7xD(377)(1) <= VNStageIntLLROutputS6xD(88)(6);
  CNStageIntLLRInputS7xD(29)(1) <= VNStageIntLLROutputS6xD(89)(0);
  CNStageIntLLRInputS7xD(102)(1) <= VNStageIntLLROutputS6xD(89)(1);
  CNStageIntLLRInputS7xD(140)(1) <= VNStageIntLLROutputS6xD(89)(2);
  CNStageIntLLRInputS7xD(184)(1) <= VNStageIntLLROutputS6xD(89)(3);
  CNStageIntLLRInputS7xD(247)(1) <= VNStageIntLLROutputS6xD(89)(4);
  CNStageIntLLRInputS7xD(355)(1) <= VNStageIntLLROutputS6xD(89)(5);
  CNStageIntLLRInputS7xD(28)(1) <= VNStageIntLLROutputS6xD(90)(0);
  CNStageIntLLRInputS7xD(85)(1) <= VNStageIntLLROutputS6xD(90)(1);
  CNStageIntLLRInputS7xD(168)(1) <= VNStageIntLLROutputS6xD(90)(2);
  CNStageIntLLRInputS7xD(175)(1) <= VNStageIntLLROutputS6xD(90)(3);
  CNStageIntLLRInputS7xD(258)(1) <= VNStageIntLLROutputS6xD(90)(4);
  CNStageIntLLRInputS7xD(307)(1) <= VNStageIntLLROutputS6xD(90)(5);
  CNStageIntLLRInputS7xD(358)(1) <= VNStageIntLLROutputS6xD(90)(6);
  CNStageIntLLRInputS7xD(27)(1) <= VNStageIntLLROutputS6xD(91)(0);
  CNStageIntLLRInputS7xD(96)(1) <= VNStageIntLLROutputS6xD(91)(1);
  CNStageIntLLRInputS7xD(158)(1) <= VNStageIntLLROutputS6xD(91)(2);
  CNStageIntLLRInputS7xD(191)(1) <= VNStageIntLLROutputS6xD(91)(3);
  CNStageIntLLRInputS7xD(269)(1) <= VNStageIntLLROutputS6xD(91)(4);
  CNStageIntLLRInputS7xD(280)(1) <= VNStageIntLLROutputS6xD(91)(5);
  CNStageIntLLRInputS7xD(344)(1) <= VNStageIntLLROutputS6xD(91)(6);
  CNStageIntLLRInputS7xD(26)(1) <= VNStageIntLLROutputS6xD(92)(0);
  CNStageIntLLRInputS7xD(103)(1) <= VNStageIntLLROutputS6xD(92)(1);
  CNStageIntLLRInputS7xD(145)(1) <= VNStageIntLLROutputS6xD(92)(2);
  CNStageIntLLRInputS7xD(195)(1) <= VNStageIntLLROutputS6xD(92)(3);
  CNStageIntLLRInputS7xD(242)(1) <= VNStageIntLLROutputS6xD(92)(4);
  CNStageIntLLRInputS7xD(324)(1) <= VNStageIntLLROutputS6xD(92)(5);
  CNStageIntLLRInputS7xD(378)(1) <= VNStageIntLLROutputS6xD(92)(6);
  CNStageIntLLRInputS7xD(25)(1) <= VNStageIntLLROutputS6xD(93)(0);
  CNStageIntLLRInputS7xD(78)(1) <= VNStageIntLLROutputS6xD(93)(1);
  CNStageIntLLRInputS7xD(164)(1) <= VNStageIntLLROutputS6xD(93)(2);
  CNStageIntLLRInputS7xD(224)(1) <= VNStageIntLLROutputS6xD(93)(3);
  CNStageIntLLRInputS7xD(231)(1) <= VNStageIntLLROutputS6xD(93)(4);
  CNStageIntLLRInputS7xD(311)(1) <= VNStageIntLLROutputS6xD(93)(5);
  CNStageIntLLRInputS7xD(340)(1) <= VNStageIntLLROutputS6xD(93)(6);
  CNStageIntLLRInputS7xD(24)(1) <= VNStageIntLLROutputS6xD(94)(0);
  CNStageIntLLRInputS7xD(92)(1) <= VNStageIntLLROutputS6xD(94)(1);
  CNStageIntLLRInputS7xD(194)(1) <= VNStageIntLLROutputS6xD(94)(2);
  CNStageIntLLRInputS7xD(329)(1) <= VNStageIntLLROutputS6xD(94)(3);
  CNStageIntLLRInputS7xD(368)(1) <= VNStageIntLLROutputS6xD(94)(4);
  CNStageIntLLRInputS7xD(23)(1) <= VNStageIntLLROutputS6xD(95)(0);
  CNStageIntLLRInputS7xD(63)(1) <= VNStageIntLLROutputS6xD(95)(1);
  CNStageIntLLRInputS7xD(134)(1) <= VNStageIntLLROutputS6xD(95)(2);
  CNStageIntLLRInputS7xD(190)(1) <= VNStageIntLLROutputS6xD(95)(3);
  CNStageIntLLRInputS7xD(234)(1) <= VNStageIntLLROutputS6xD(95)(4);
  CNStageIntLLRInputS7xD(303)(1) <= VNStageIntLLROutputS6xD(95)(5);
  CNStageIntLLRInputS7xD(352)(1) <= VNStageIntLLROutputS6xD(95)(6);
  CNStageIntLLRInputS7xD(22)(1) <= VNStageIntLLROutputS6xD(96)(0);
  CNStageIntLLRInputS7xD(98)(1) <= VNStageIntLLROutputS6xD(96)(1);
  CNStageIntLLRInputS7xD(150)(1) <= VNStageIntLLROutputS6xD(96)(2);
  CNStageIntLLRInputS7xD(172)(1) <= VNStageIntLLROutputS6xD(96)(3);
  CNStageIntLLRInputS7xD(251)(1) <= VNStageIntLLROutputS6xD(96)(4);
  CNStageIntLLRInputS7xD(380)(1) <= VNStageIntLLROutputS6xD(96)(5);
  CNStageIntLLRInputS7xD(21)(1) <= VNStageIntLLROutputS6xD(97)(0);
  CNStageIntLLRInputS7xD(65)(1) <= VNStageIntLLROutputS6xD(97)(1);
  CNStageIntLLRInputS7xD(142)(1) <= VNStageIntLLROutputS6xD(97)(2);
  CNStageIntLLRInputS7xD(180)(1) <= VNStageIntLLROutputS6xD(97)(3);
  CNStageIntLLRInputS7xD(260)(1) <= VNStageIntLLROutputS6xD(97)(4);
  CNStageIntLLRInputS7xD(316)(1) <= VNStageIntLLROutputS6xD(97)(5);
  CNStageIntLLRInputS7xD(370)(1) <= VNStageIntLLROutputS6xD(97)(6);
  CNStageIntLLRInputS7xD(20)(1) <= VNStageIntLLROutputS6xD(98)(0);
  CNStageIntLLRInputS7xD(116)(1) <= VNStageIntLLROutputS6xD(98)(1);
  CNStageIntLLRInputS7xD(199)(1) <= VNStageIntLLROutputS6xD(98)(2);
  CNStageIntLLRInputS7xD(255)(1) <= VNStageIntLLROutputS6xD(98)(3);
  CNStageIntLLRInputS7xD(308)(1) <= VNStageIntLLROutputS6xD(98)(4);
  CNStageIntLLRInputS7xD(356)(1) <= VNStageIntLLROutputS6xD(98)(5);
  CNStageIntLLRInputS7xD(19)(1) <= VNStageIntLLROutputS6xD(99)(0);
  CNStageIntLLRInputS7xD(76)(1) <= VNStageIntLLROutputS6xD(99)(1);
  CNStageIntLLRInputS7xD(126)(1) <= VNStageIntLLROutputS6xD(99)(2);
  CNStageIntLLRInputS7xD(198)(1) <= VNStageIntLLROutputS6xD(99)(3);
  CNStageIntLLRInputS7xD(261)(1) <= VNStageIntLLROutputS6xD(99)(4);
  CNStageIntLLRInputS7xD(285)(1) <= VNStageIntLLROutputS6xD(99)(5);
  CNStageIntLLRInputS7xD(376)(1) <= VNStageIntLLROutputS6xD(99)(6);
  CNStageIntLLRInputS7xD(18)(1) <= VNStageIntLLROutputS6xD(100)(0);
  CNStageIntLLRInputS7xD(94)(1) <= VNStageIntLLROutputS6xD(100)(1);
  CNStageIntLLRInputS7xD(120)(1) <= VNStageIntLLROutputS6xD(100)(2);
  CNStageIntLLRInputS7xD(178)(1) <= VNStageIntLLROutputS6xD(100)(3);
  CNStageIntLLRInputS7xD(250)(1) <= VNStageIntLLROutputS6xD(100)(4);
  CNStageIntLLRInputS7xD(295)(1) <= VNStageIntLLROutputS6xD(100)(5);
  CNStageIntLLRInputS7xD(349)(1) <= VNStageIntLLROutputS6xD(100)(6);
  CNStageIntLLRInputS7xD(17)(1) <= VNStageIntLLROutputS6xD(101)(0);
  CNStageIntLLRInputS7xD(58)(1) <= VNStageIntLLROutputS6xD(101)(1);
  CNStageIntLLRInputS7xD(123)(1) <= VNStageIntLLROutputS6xD(101)(2);
  CNStageIntLLRInputS7xD(211)(1) <= VNStageIntLLROutputS6xD(101)(3);
  CNStageIntLLRInputS7xD(273)(1) <= VNStageIntLLROutputS6xD(101)(4);
  CNStageIntLLRInputS7xD(289)(1) <= VNStageIntLLROutputS6xD(101)(5);
  CNStageIntLLRInputS7xD(346)(1) <= VNStageIntLLROutputS6xD(101)(6);
  CNStageIntLLRInputS7xD(16)(1) <= VNStageIntLLROutputS6xD(102)(0);
  CNStageIntLLRInputS7xD(59)(1) <= VNStageIntLLROutputS6xD(102)(1);
  CNStageIntLLRInputS7xD(113)(1) <= VNStageIntLLROutputS6xD(102)(2);
  CNStageIntLLRInputS7xD(214)(1) <= VNStageIntLLROutputS6xD(102)(3);
  CNStageIntLLRInputS7xD(226)(1) <= VNStageIntLLROutputS6xD(102)(4);
  CNStageIntLLRInputS7xD(361)(1) <= VNStageIntLLROutputS6xD(102)(5);
  CNStageIntLLRInputS7xD(15)(1) <= VNStageIntLLROutputS6xD(103)(0);
  CNStageIntLLRInputS7xD(93)(1) <= VNStageIntLLROutputS6xD(103)(1);
  CNStageIntLLRInputS7xD(151)(1) <= VNStageIntLLROutputS6xD(103)(2);
  CNStageIntLLRInputS7xD(200)(1) <= VNStageIntLLROutputS6xD(103)(3);
  CNStageIntLLRInputS7xD(265)(1) <= VNStageIntLLROutputS6xD(103)(4);
  CNStageIntLLRInputS7xD(284)(1) <= VNStageIntLLROutputS6xD(103)(5);
  CNStageIntLLRInputS7xD(354)(1) <= VNStageIntLLROutputS6xD(103)(6);
  CNStageIntLLRInputS7xD(14)(1) <= VNStageIntLLROutputS6xD(104)(0);
  CNStageIntLLRInputS7xD(86)(1) <= VNStageIntLLROutputS6xD(104)(1);
  CNStageIntLLRInputS7xD(133)(1) <= VNStageIntLLROutputS6xD(104)(2);
  CNStageIntLLRInputS7xD(179)(1) <= VNStageIntLLROutputS6xD(104)(3);
  CNStageIntLLRInputS7xD(267)(1) <= VNStageIntLLROutputS6xD(104)(4);
  CNStageIntLLRInputS7xD(317)(1) <= VNStageIntLLROutputS6xD(104)(5);
  CNStageIntLLRInputS7xD(13)(1) <= VNStageIntLLROutputS6xD(105)(0);
  CNStageIntLLRInputS7xD(146)(1) <= VNStageIntLLROutputS6xD(105)(1);
  CNStageIntLLRInputS7xD(197)(1) <= VNStageIntLLROutputS6xD(105)(2);
  CNStageIntLLRInputS7xD(237)(1) <= VNStageIntLLROutputS6xD(105)(3);
  CNStageIntLLRInputS7xD(300)(1) <= VNStageIntLLROutputS6xD(105)(4);
  CNStageIntLLRInputS7xD(338)(1) <= VNStageIntLLROutputS6xD(105)(5);
  CNStageIntLLRInputS7xD(12)(1) <= VNStageIntLLROutputS6xD(106)(0);
  CNStageIntLLRInputS7xD(157)(1) <= VNStageIntLLROutputS6xD(106)(1);
  CNStageIntLLRInputS7xD(223)(1) <= VNStageIntLLROutputS6xD(106)(2);
  CNStageIntLLRInputS7xD(272)(1) <= VNStageIntLLROutputS6xD(106)(3);
  CNStageIntLLRInputS7xD(312)(1) <= VNStageIntLLROutputS6xD(106)(4);
  CNStageIntLLRInputS7xD(333)(1) <= VNStageIntLLROutputS6xD(106)(5);
  CNStageIntLLRInputS7xD(110)(1) <= VNStageIntLLROutputS6xD(107)(0);
  CNStageIntLLRInputS7xD(127)(1) <= VNStageIntLLROutputS6xD(107)(1);
  CNStageIntLLRInputS7xD(207)(1) <= VNStageIntLLROutputS6xD(107)(2);
  CNStageIntLLRInputS7xD(230)(1) <= VNStageIntLLROutputS6xD(107)(3);
  CNStageIntLLRInputS7xD(323)(1) <= VNStageIntLLROutputS6xD(107)(4);
  CNStageIntLLRInputS7xD(335)(1) <= VNStageIntLLROutputS6xD(107)(5);
  CNStageIntLLRInputS7xD(11)(1) <= VNStageIntLLROutputS6xD(108)(0);
  CNStageIntLLRInputS7xD(105)(1) <= VNStageIntLLROutputS6xD(108)(1);
  CNStageIntLLRInputS7xD(115)(1) <= VNStageIntLLROutputS6xD(108)(2);
  CNStageIntLLRInputS7xD(181)(1) <= VNStageIntLLROutputS6xD(108)(3);
  CNStageIntLLRInputS7xD(238)(1) <= VNStageIntLLROutputS6xD(108)(4);
  CNStageIntLLRInputS7xD(296)(1) <= VNStageIntLLROutputS6xD(108)(5);
  CNStageIntLLRInputS7xD(10)(1) <= VNStageIntLLROutputS6xD(109)(0);
  CNStageIntLLRInputS7xD(100)(1) <= VNStageIntLLROutputS6xD(109)(1);
  CNStageIntLLRInputS7xD(160)(1) <= VNStageIntLLROutputS6xD(109)(2);
  CNStageIntLLRInputS7xD(171)(1) <= VNStageIntLLROutputS6xD(109)(3);
  CNStageIntLLRInputS7xD(266)(1) <= VNStageIntLLROutputS6xD(109)(4);
  CNStageIntLLRInputS7xD(362)(1) <= VNStageIntLLROutputS6xD(109)(5);
  CNStageIntLLRInputS7xD(9)(1) <= VNStageIntLLROutputS6xD(110)(0);
  CNStageIntLLRInputS7xD(83)(1) <= VNStageIntLLROutputS6xD(110)(1);
  CNStageIntLLRInputS7xD(118)(1) <= VNStageIntLLROutputS6xD(110)(2);
  CNStageIntLLRInputS7xD(212)(1) <= VNStageIntLLROutputS6xD(110)(3);
  CNStageIntLLRInputS7xD(225)(1) <= VNStageIntLLROutputS6xD(110)(4);
  CNStageIntLLRInputS7xD(326)(1) <= VNStageIntLLROutputS6xD(110)(5);
  CNStageIntLLRInputS7xD(345)(1) <= VNStageIntLLROutputS6xD(110)(6);
  CNStageIntLLRInputS7xD(8)(1) <= VNStageIntLLROutputS6xD(111)(0);
  CNStageIntLLRInputS7xD(90)(1) <= VNStageIntLLROutputS6xD(111)(1);
  CNStageIntLLRInputS7xD(138)(1) <= VNStageIntLLROutputS6xD(111)(2);
  CNStageIntLLRInputS7xD(177)(1) <= VNStageIntLLROutputS6xD(111)(3);
  CNStageIntLLRInputS7xD(252)(1) <= VNStageIntLLROutputS6xD(111)(4);
  CNStageIntLLRInputS7xD(287)(1) <= VNStageIntLLROutputS6xD(111)(5);
  CNStageIntLLRInputS7xD(357)(1) <= VNStageIntLLROutputS6xD(111)(6);
  CNStageIntLLRInputS7xD(7)(1) <= VNStageIntLLROutputS6xD(112)(0);
  CNStageIntLLRInputS7xD(54)(1) <= VNStageIntLLROutputS6xD(112)(1);
  CNStageIntLLRInputS7xD(148)(1) <= VNStageIntLLROutputS6xD(112)(2);
  CNStageIntLLRInputS7xD(205)(1) <= VNStageIntLLROutputS6xD(112)(3);
  CNStageIntLLRInputS7xD(233)(1) <= VNStageIntLLROutputS6xD(112)(4);
  CNStageIntLLRInputS7xD(305)(1) <= VNStageIntLLROutputS6xD(112)(5);
  CNStageIntLLRInputS7xD(369)(1) <= VNStageIntLLROutputS6xD(112)(6);
  CNStageIntLLRInputS7xD(6)(1) <= VNStageIntLLROutputS6xD(113)(0);
  CNStageIntLLRInputS7xD(108)(1) <= VNStageIntLLROutputS6xD(113)(1);
  CNStageIntLLRInputS7xD(143)(1) <= VNStageIntLLROutputS6xD(113)(2);
  CNStageIntLLRInputS7xD(202)(1) <= VNStageIntLLROutputS6xD(113)(3);
  CNStageIntLLRInputS7xD(253)(1) <= VNStageIntLLROutputS6xD(113)(4);
  CNStageIntLLRInputS7xD(314)(1) <= VNStageIntLLROutputS6xD(113)(5);
  CNStageIntLLRInputS7xD(339)(1) <= VNStageIntLLROutputS6xD(113)(6);
  CNStageIntLLRInputS7xD(5)(1) <= VNStageIntLLROutputS6xD(114)(0);
  CNStageIntLLRInputS7xD(88)(1) <= VNStageIntLLROutputS6xD(114)(1);
  CNStageIntLLRInputS7xD(149)(1) <= VNStageIntLLROutputS6xD(114)(2);
  CNStageIntLLRInputS7xD(216)(1) <= VNStageIntLLROutputS6xD(114)(3);
  CNStageIntLLRInputS7xD(268)(1) <= VNStageIntLLROutputS6xD(114)(4);
  CNStageIntLLRInputS7xD(309)(1) <= VNStageIntLLROutputS6xD(114)(5);
  CNStageIntLLRInputS7xD(4)(1) <= VNStageIntLLROutputS6xD(115)(0);
  CNStageIntLLRInputS7xD(68)(1) <= VNStageIntLLROutputS6xD(115)(1);
  CNStageIntLLRInputS7xD(137)(1) <= VNStageIntLLROutputS6xD(115)(2);
  CNStageIntLLRInputS7xD(209)(1) <= VNStageIntLLROutputS6xD(115)(3);
  CNStageIntLLRInputS7xD(264)(1) <= VNStageIntLLROutputS6xD(115)(4);
  CNStageIntLLRInputS7xD(315)(1) <= VNStageIntLLROutputS6xD(115)(5);
  CNStageIntLLRInputS7xD(372)(1) <= VNStageIntLLROutputS6xD(115)(6);
  CNStageIntLLRInputS7xD(71)(1) <= VNStageIntLLROutputS6xD(116)(0);
  CNStageIntLLRInputS7xD(163)(1) <= VNStageIntLLROutputS6xD(116)(1);
  CNStageIntLLRInputS7xD(187)(1) <= VNStageIntLLROutputS6xD(116)(2);
  CNStageIntLLRInputS7xD(228)(1) <= VNStageIntLLROutputS6xD(116)(3);
  CNStageIntLLRInputS7xD(304)(1) <= VNStageIntLLROutputS6xD(116)(4);
  CNStageIntLLRInputS7xD(3)(1) <= VNStageIntLLROutputS6xD(117)(0);
  CNStageIntLLRInputS7xD(55)(1) <= VNStageIntLLROutputS6xD(117)(1);
  CNStageIntLLRInputS7xD(111)(1) <= VNStageIntLLROutputS6xD(117)(2);
  CNStageIntLLRInputS7xD(196)(1) <= VNStageIntLLROutputS6xD(117)(3);
  CNStageIntLLRInputS7xD(2)(1) <= VNStageIntLLROutputS6xD(118)(0);
  CNStageIntLLRInputS7xD(89)(1) <= VNStageIntLLROutputS6xD(118)(1);
  CNStageIntLLRInputS7xD(152)(1) <= VNStageIntLLROutputS6xD(118)(2);
  CNStageIntLLRInputS7xD(249)(1) <= VNStageIntLLROutputS6xD(118)(3);
  CNStageIntLLRInputS7xD(282)(1) <= VNStageIntLLROutputS6xD(118)(4);
  CNStageIntLLRInputS7xD(359)(1) <= VNStageIntLLROutputS6xD(118)(5);
  CNStageIntLLRInputS7xD(1)(1) <= VNStageIntLLROutputS6xD(119)(0);
  CNStageIntLLRInputS7xD(107)(1) <= VNStageIntLLROutputS6xD(119)(1);
  CNStageIntLLRInputS7xD(154)(1) <= VNStageIntLLROutputS6xD(119)(2);
  CNStageIntLLRInputS7xD(227)(1) <= VNStageIntLLROutputS6xD(119)(3);
  CNStageIntLLRInputS7xD(319)(1) <= VNStageIntLLROutputS6xD(119)(4);
  CNStageIntLLRInputS7xD(0)(1) <= VNStageIntLLROutputS6xD(120)(0);
  CNStageIntLLRInputS7xD(80)(1) <= VNStageIntLLROutputS6xD(120)(1);
  CNStageIntLLRInputS7xD(321)(1) <= VNStageIntLLROutputS6xD(120)(2);
  CNStageIntLLRInputS7xD(360)(1) <= VNStageIntLLROutputS6xD(120)(3);
  CNStageIntLLRInputS7xD(64)(1) <= VNStageIntLLROutputS6xD(121)(0);
  CNStageIntLLRInputS7xD(161)(1) <= VNStageIntLLROutputS6xD(121)(1);
  CNStageIntLLRInputS7xD(217)(1) <= VNStageIntLLROutputS6xD(121)(2);
  CNStageIntLLRInputS7xD(236)(1) <= VNStageIntLLROutputS6xD(121)(3);
  CNStageIntLLRInputS7xD(291)(1) <= VNStageIntLLROutputS6xD(121)(4);
  CNStageIntLLRInputS7xD(350)(1) <= VNStageIntLLROutputS6xD(121)(5);
  CNStageIntLLRInputS7xD(91)(1) <= VNStageIntLLROutputS6xD(122)(0);
  CNStageIntLLRInputS7xD(114)(1) <= VNStageIntLLROutputS6xD(122)(1);
  CNStageIntLLRInputS7xD(201)(1) <= VNStageIntLLROutputS6xD(122)(2);
  CNStageIntLLRInputS7xD(241)(1) <= VNStageIntLLROutputS6xD(122)(3);
  CNStageIntLLRInputS7xD(327)(1) <= VNStageIntLLROutputS6xD(122)(4);
  CNStageIntLLRInputS7xD(375)(1) <= VNStageIntLLROutputS6xD(122)(5);
  CNStageIntLLRInputS7xD(82)(1) <= VNStageIntLLROutputS6xD(123)(0);
  CNStageIntLLRInputS7xD(122)(1) <= VNStageIntLLROutputS6xD(123)(1);
  CNStageIntLLRInputS7xD(213)(1) <= VNStageIntLLROutputS6xD(123)(2);
  CNStageIntLLRInputS7xD(279)(1) <= VNStageIntLLROutputS6xD(123)(3);
  CNStageIntLLRInputS7xD(382)(1) <= VNStageIntLLROutputS6xD(123)(4);
  CNStageIntLLRInputS7xD(69)(1) <= VNStageIntLLROutputS6xD(124)(0);
  CNStageIntLLRInputS7xD(153)(1) <= VNStageIntLLROutputS6xD(124)(1);
  CNStageIntLLRInputS7xD(240)(1) <= VNStageIntLLROutputS6xD(124)(2);
  CNStageIntLLRInputS7xD(292)(1) <= VNStageIntLLROutputS6xD(124)(3);
  CNStageIntLLRInputS7xD(364)(1) <= VNStageIntLLROutputS6xD(124)(4);
  CNStageIntLLRInputS7xD(87)(1) <= VNStageIntLLROutputS6xD(125)(0);
  CNStageIntLLRInputS7xD(169)(1) <= VNStageIntLLROutputS6xD(125)(1);
  CNStageIntLLRInputS7xD(320)(1) <= VNStageIntLLROutputS6xD(125)(2);
  CNStageIntLLRInputS7xD(366)(1) <= VNStageIntLLROutputS6xD(125)(3);
  CNStageIntLLRInputS7xD(60)(1) <= VNStageIntLLROutputS6xD(126)(0);
  CNStageIntLLRInputS7xD(139)(1) <= VNStageIntLLROutputS6xD(126)(1);
  CNStageIntLLRInputS7xD(186)(1) <= VNStageIntLLROutputS6xD(126)(2);
  CNStageIntLLRInputS7xD(271)(1) <= VNStageIntLLROutputS6xD(126)(3);
  CNStageIntLLRInputS7xD(281)(1) <= VNStageIntLLROutputS6xD(126)(4);
  CNStageIntLLRInputS7xD(334)(1) <= VNStageIntLLROutputS6xD(126)(5);
  CNStageIntLLRInputS7xD(52)(1) <= VNStageIntLLROutputS6xD(127)(0);
  CNStageIntLLRInputS7xD(57)(1) <= VNStageIntLLROutputS6xD(127)(1);
  CNStageIntLLRInputS7xD(117)(1) <= VNStageIntLLROutputS6xD(127)(2);
  CNStageIntLLRInputS7xD(173)(1) <= VNStageIntLLROutputS6xD(127)(3);
  CNStageIntLLRInputS7xD(277)(1) <= VNStageIntLLROutputS6xD(127)(4);
  CNStageIntLLRInputS7xD(306)(1) <= VNStageIntLLROutputS6xD(127)(5);
  CNStageIntLLRInputS7xD(373)(1) <= VNStageIntLLROutputS6xD(127)(6);
  CNStageIntLLRInputS7xD(53)(2) <= VNStageIntLLROutputS6xD(128)(0);
  CNStageIntLLRInputS7xD(108)(2) <= VNStageIntLLROutputS6xD(128)(1);
  CNStageIntLLRInputS7xD(129)(2) <= VNStageIntLLROutputS6xD(128)(2);
  CNStageIntLLRInputS7xD(198)(2) <= VNStageIntLLROutputS6xD(128)(3);
  CNStageIntLLRInputS7xD(244)(2) <= VNStageIntLLROutputS6xD(128)(4);
  CNStageIntLLRInputS7xD(298)(2) <= VNStageIntLLROutputS6xD(128)(5);
  CNStageIntLLRInputS7xD(341)(2) <= VNStageIntLLROutputS6xD(128)(6);
  CNStageIntLLRInputS7xD(51)(2) <= VNStageIntLLROutputS6xD(129)(0);
  CNStageIntLLRInputS7xD(56)(2) <= VNStageIntLLROutputS6xD(129)(1);
  CNStageIntLLRInputS7xD(116)(2) <= VNStageIntLLROutputS6xD(129)(2);
  CNStageIntLLRInputS7xD(172)(2) <= VNStageIntLLROutputS6xD(129)(3);
  CNStageIntLLRInputS7xD(276)(2) <= VNStageIntLLROutputS6xD(129)(4);
  CNStageIntLLRInputS7xD(305)(2) <= VNStageIntLLROutputS6xD(129)(5);
  CNStageIntLLRInputS7xD(372)(2) <= VNStageIntLLROutputS6xD(129)(6);
  CNStageIntLLRInputS7xD(50)(2) <= VNStageIntLLROutputS6xD(130)(0);
  CNStageIntLLRInputS7xD(73)(2) <= VNStageIntLLROutputS6xD(130)(1);
  CNStageIntLLRInputS7xD(140)(2) <= VNStageIntLLROutputS6xD(130)(2);
  CNStageIntLLRInputS7xD(188)(2) <= VNStageIntLLROutputS6xD(130)(3);
  CNStageIntLLRInputS7xD(245)(2) <= VNStageIntLLROutputS6xD(130)(4);
  CNStageIntLLRInputS7xD(285)(2) <= VNStageIntLLROutputS6xD(130)(5);
  CNStageIntLLRInputS7xD(65)(2) <= VNStageIntLLROutputS6xD(131)(0);
  CNStageIntLLRInputS7xD(154)(2) <= VNStageIntLLROutputS6xD(131)(1);
  CNStageIntLLRInputS7xD(206)(2) <= VNStageIntLLROutputS6xD(131)(2);
  CNStageIntLLRInputS7xD(243)(2) <= VNStageIntLLROutputS6xD(131)(3);
  CNStageIntLLRInputS7xD(307)(2) <= VNStageIntLLROutputS6xD(131)(4);
  CNStageIntLLRInputS7xD(334)(2) <= VNStageIntLLROutputS6xD(131)(5);
  CNStageIntLLRInputS7xD(49)(2) <= VNStageIntLLROutputS6xD(132)(0);
  CNStageIntLLRInputS7xD(151)(2) <= VNStageIntLLROutputS6xD(132)(1);
  CNStageIntLLRInputS7xD(214)(2) <= VNStageIntLLROutputS6xD(132)(2);
  CNStageIntLLRInputS7xD(274)(2) <= VNStageIntLLROutputS6xD(132)(3);
  CNStageIntLLRInputS7xD(321)(2) <= VNStageIntLLROutputS6xD(132)(4);
  CNStageIntLLRInputS7xD(364)(2) <= VNStageIntLLROutputS6xD(132)(5);
  CNStageIntLLRInputS7xD(48)(2) <= VNStageIntLLROutputS6xD(133)(0);
  CNStageIntLLRInputS7xD(209)(2) <= VNStageIntLLROutputS6xD(133)(1);
  CNStageIntLLRInputS7xD(255)(2) <= VNStageIntLLROutputS6xD(133)(2);
  CNStageIntLLRInputS7xD(317)(2) <= VNStageIntLLROutputS6xD(133)(3);
  CNStageIntLLRInputS7xD(380)(2) <= VNStageIntLLROutputS6xD(133)(4);
  CNStageIntLLRInputS7xD(47)(2) <= VNStageIntLLROutputS6xD(134)(0);
  CNStageIntLLRInputS7xD(100)(2) <= VNStageIntLLROutputS6xD(134)(1);
  CNStageIntLLRInputS7xD(134)(2) <= VNStageIntLLROutputS6xD(134)(2);
  CNStageIntLLRInputS7xD(258)(2) <= VNStageIntLLROutputS6xD(134)(3);
  CNStageIntLLRInputS7xD(46)(2) <= VNStageIntLLROutputS6xD(135)(0);
  CNStageIntLLRInputS7xD(103)(2) <= VNStageIntLLROutputS6xD(135)(1);
  CNStageIntLLRInputS7xD(135)(2) <= VNStageIntLLROutputS6xD(135)(2);
  CNStageIntLLRInputS7xD(205)(2) <= VNStageIntLLROutputS6xD(135)(3);
  CNStageIntLLRInputS7xD(45)(2) <= VNStageIntLLROutputS6xD(136)(0);
  CNStageIntLLRInputS7xD(94)(2) <= VNStageIntLLROutputS6xD(136)(1);
  CNStageIntLLRInputS7xD(111)(2) <= VNStageIntLLROutputS6xD(136)(2);
  CNStageIntLLRInputS7xD(175)(2) <= VNStageIntLLROutputS6xD(136)(3);
  CNStageIntLLRInputS7xD(275)(2) <= VNStageIntLLROutputS6xD(136)(4);
  CNStageIntLLRInputS7xD(301)(2) <= VNStageIntLLROutputS6xD(136)(5);
  CNStageIntLLRInputS7xD(352)(2) <= VNStageIntLLROutputS6xD(136)(6);
  CNStageIntLLRInputS7xD(44)(2) <= VNStageIntLLROutputS6xD(137)(0);
  CNStageIntLLRInputS7xD(74)(2) <= VNStageIntLLROutputS6xD(137)(1);
  CNStageIntLLRInputS7xD(161)(2) <= VNStageIntLLROutputS6xD(137)(2);
  CNStageIntLLRInputS7xD(182)(2) <= VNStageIntLLROutputS6xD(137)(3);
  CNStageIntLLRInputS7xD(242)(2) <= VNStageIntLLROutputS6xD(137)(4);
  CNStageIntLLRInputS7xD(282)(2) <= VNStageIntLLROutputS6xD(137)(5);
  CNStageIntLLRInputS7xD(366)(2) <= VNStageIntLLROutputS6xD(137)(6);
  CNStageIntLLRInputS7xD(43)(2) <= VNStageIntLLROutputS6xD(138)(0);
  CNStageIntLLRInputS7xD(55)(2) <= VNStageIntLLROutputS6xD(138)(1);
  CNStageIntLLRInputS7xD(120)(2) <= VNStageIntLLROutputS6xD(138)(2);
  CNStageIntLLRInputS7xD(218)(2) <= VNStageIntLLROutputS6xD(138)(3);
  CNStageIntLLRInputS7xD(268)(2) <= VNStageIntLLROutputS6xD(138)(4);
  CNStageIntLLRInputS7xD(327)(2) <= VNStageIntLLROutputS6xD(138)(5);
  CNStageIntLLRInputS7xD(362)(2) <= VNStageIntLLROutputS6xD(138)(6);
  CNStageIntLLRInputS7xD(42)(2) <= VNStageIntLLROutputS6xD(139)(0);
  CNStageIntLLRInputS7xD(69)(2) <= VNStageIntLLROutputS6xD(139)(1);
  CNStageIntLLRInputS7xD(124)(2) <= VNStageIntLLROutputS6xD(139)(2);
  CNStageIntLLRInputS7xD(220)(2) <= VNStageIntLLROutputS6xD(139)(3);
  CNStageIntLLRInputS7xD(252)(2) <= VNStageIntLLROutputS6xD(139)(4);
  CNStageIntLLRInputS7xD(289)(2) <= VNStageIntLLROutputS6xD(139)(5);
  CNStageIntLLRInputS7xD(383)(2) <= VNStageIntLLROutputS6xD(139)(6);
  CNStageIntLLRInputS7xD(41)(2) <= VNStageIntLLROutputS6xD(140)(0);
  CNStageIntLLRInputS7xD(80)(2) <= VNStageIntLLROutputS6xD(140)(1);
  CNStageIntLLRInputS7xD(170)(2) <= VNStageIntLLROutputS6xD(140)(2);
  CNStageIntLLRInputS7xD(191)(2) <= VNStageIntLLROutputS6xD(140)(3);
  CNStageIntLLRInputS7xD(277)(2) <= VNStageIntLLROutputS6xD(140)(4);
  CNStageIntLLRInputS7xD(293)(2) <= VNStageIntLLROutputS6xD(140)(5);
  CNStageIntLLRInputS7xD(346)(2) <= VNStageIntLLROutputS6xD(140)(6);
  CNStageIntLLRInputS7xD(123)(2) <= VNStageIntLLROutputS6xD(141)(0);
  CNStageIntLLRInputS7xD(173)(2) <= VNStageIntLLROutputS6xD(141)(1);
  CNStageIntLLRInputS7xD(269)(2) <= VNStageIntLLROutputS6xD(141)(2);
  CNStageIntLLRInputS7xD(332)(2) <= VNStageIntLLROutputS6xD(141)(3);
  CNStageIntLLRInputS7xD(347)(2) <= VNStageIntLLROutputS6xD(141)(4);
  CNStageIntLLRInputS7xD(40)(2) <= VNStageIntLLROutputS6xD(142)(0);
  CNStageIntLLRInputS7xD(96)(2) <= VNStageIntLLROutputS6xD(142)(1);
  CNStageIntLLRInputS7xD(118)(2) <= VNStageIntLLROutputS6xD(142)(2);
  CNStageIntLLRInputS7xD(256)(2) <= VNStageIntLLROutputS6xD(142)(3);
  CNStageIntLLRInputS7xD(382)(2) <= VNStageIntLLROutputS6xD(142)(4);
  CNStageIntLLRInputS7xD(39)(2) <= VNStageIntLLROutputS6xD(143)(0);
  CNStageIntLLRInputS7xD(83)(2) <= VNStageIntLLROutputS6xD(143)(1);
  CNStageIntLLRInputS7xD(158)(2) <= VNStageIntLLROutputS6xD(143)(2);
  CNStageIntLLRInputS7xD(192)(2) <= VNStageIntLLROutputS6xD(143)(3);
  CNStageIntLLRInputS7xD(273)(2) <= VNStageIntLLROutputS6xD(143)(4);
  CNStageIntLLRInputS7xD(287)(2) <= VNStageIntLLROutputS6xD(143)(5);
  CNStageIntLLRInputS7xD(373)(2) <= VNStageIntLLROutputS6xD(143)(6);
  CNStageIntLLRInputS7xD(38)(2) <= VNStageIntLLROutputS6xD(144)(0);
  CNStageIntLLRInputS7xD(98)(2) <= VNStageIntLLROutputS6xD(144)(1);
  CNStageIntLLRInputS7xD(166)(2) <= VNStageIntLLROutputS6xD(144)(2);
  CNStageIntLLRInputS7xD(219)(2) <= VNStageIntLLROutputS6xD(144)(3);
  CNStageIntLLRInputS7xD(249)(2) <= VNStageIntLLROutputS6xD(144)(4);
  CNStageIntLLRInputS7xD(324)(2) <= VNStageIntLLROutputS6xD(144)(5);
  CNStageIntLLRInputS7xD(333)(2) <= VNStageIntLLROutputS6xD(144)(6);
  CNStageIntLLRInputS7xD(37)(2) <= VNStageIntLLROutputS6xD(145)(0);
  CNStageIntLLRInputS7xD(61)(2) <= VNStageIntLLROutputS6xD(145)(1);
  CNStageIntLLRInputS7xD(130)(2) <= VNStageIntLLROutputS6xD(145)(2);
  CNStageIntLLRInputS7xD(181)(2) <= VNStageIntLLROutputS6xD(145)(3);
  CNStageIntLLRInputS7xD(247)(2) <= VNStageIntLLROutputS6xD(145)(4);
  CNStageIntLLRInputS7xD(331)(2) <= VNStageIntLLROutputS6xD(145)(5);
  CNStageIntLLRInputS7xD(336)(2) <= VNStageIntLLROutputS6xD(145)(6);
  CNStageIntLLRInputS7xD(36)(2) <= VNStageIntLLROutputS6xD(146)(0);
  CNStageIntLLRInputS7xD(71)(2) <= VNStageIntLLROutputS6xD(146)(1);
  CNStageIntLLRInputS7xD(128)(2) <= VNStageIntLLROutputS6xD(146)(2);
  CNStageIntLLRInputS7xD(261)(2) <= VNStageIntLLROutputS6xD(146)(3);
  CNStageIntLLRInputS7xD(299)(2) <= VNStageIntLLROutputS6xD(146)(4);
  CNStageIntLLRInputS7xD(35)(2) <= VNStageIntLLROutputS6xD(147)(0);
  CNStageIntLLRInputS7xD(66)(2) <= VNStageIntLLROutputS6xD(147)(1);
  CNStageIntLLRInputS7xD(164)(2) <= VNStageIntLLROutputS6xD(147)(2);
  CNStageIntLLRInputS7xD(187)(2) <= VNStageIntLLROutputS6xD(147)(3);
  CNStageIntLLRInputS7xD(253)(2) <= VNStageIntLLROutputS6xD(147)(4);
  CNStageIntLLRInputS7xD(297)(2) <= VNStageIntLLROutputS6xD(147)(5);
  CNStageIntLLRInputS7xD(335)(2) <= VNStageIntLLROutputS6xD(147)(6);
  CNStageIntLLRInputS7xD(34)(2) <= VNStageIntLLROutputS6xD(148)(0);
  CNStageIntLLRInputS7xD(72)(2) <= VNStageIntLLROutputS6xD(148)(1);
  CNStageIntLLRInputS7xD(143)(2) <= VNStageIntLLROutputS6xD(148)(2);
  CNStageIntLLRInputS7xD(207)(2) <= VNStageIntLLROutputS6xD(148)(3);
  CNStageIntLLRInputS7xD(231)(2) <= VNStageIntLLROutputS6xD(148)(4);
  CNStageIntLLRInputS7xD(329)(2) <= VNStageIntLLROutputS6xD(148)(5);
  CNStageIntLLRInputS7xD(33)(2) <= VNStageIntLLROutputS6xD(149)(0);
  CNStageIntLLRInputS7xD(60)(2) <= VNStageIntLLROutputS6xD(149)(1);
  CNStageIntLLRInputS7xD(146)(2) <= VNStageIntLLROutputS6xD(149)(2);
  CNStageIntLLRInputS7xD(221)(2) <= VNStageIntLLROutputS6xD(149)(3);
  CNStageIntLLRInputS7xD(241)(2) <= VNStageIntLLROutputS6xD(149)(4);
  CNStageIntLLRInputS7xD(309)(2) <= VNStageIntLLROutputS6xD(149)(5);
  CNStageIntLLRInputS7xD(370)(2) <= VNStageIntLLROutputS6xD(149)(6);
  CNStageIntLLRInputS7xD(32)(2) <= VNStageIntLLROutputS6xD(150)(0);
  CNStageIntLLRInputS7xD(86)(2) <= VNStageIntLLROutputS6xD(150)(1);
  CNStageIntLLRInputS7xD(131)(2) <= VNStageIntLLROutputS6xD(150)(2);
  CNStageIntLLRInputS7xD(217)(2) <= VNStageIntLLROutputS6xD(150)(3);
  CNStageIntLLRInputS7xD(312)(2) <= VNStageIntLLROutputS6xD(150)(4);
  CNStageIntLLRInputS7xD(378)(2) <= VNStageIntLLROutputS6xD(150)(5);
  CNStageIntLLRInputS7xD(31)(2) <= VNStageIntLLROutputS6xD(151)(0);
  CNStageIntLLRInputS7xD(92)(2) <= VNStageIntLLROutputS6xD(151)(1);
  CNStageIntLLRInputS7xD(165)(2) <= VNStageIntLLROutputS6xD(151)(2);
  CNStageIntLLRInputS7xD(184)(2) <= VNStageIntLLROutputS6xD(151)(3);
  CNStageIntLLRInputS7xD(238)(2) <= VNStageIntLLROutputS6xD(151)(4);
  CNStageIntLLRInputS7xD(342)(2) <= VNStageIntLLROutputS6xD(151)(5);
  CNStageIntLLRInputS7xD(30)(2) <= VNStageIntLLROutputS6xD(152)(0);
  CNStageIntLLRInputS7xD(76)(2) <= VNStageIntLLROutputS6xD(152)(1);
  CNStageIntLLRInputS7xD(127)(2) <= VNStageIntLLROutputS6xD(152)(2);
  CNStageIntLLRInputS7xD(202)(2) <= VNStageIntLLROutputS6xD(152)(3);
  CNStageIntLLRInputS7xD(228)(2) <= VNStageIntLLROutputS6xD(152)(4);
  CNStageIntLLRInputS7xD(330)(2) <= VNStageIntLLROutputS6xD(152)(5);
  CNStageIntLLRInputS7xD(340)(2) <= VNStageIntLLROutputS6xD(152)(6);
  CNStageIntLLRInputS7xD(29)(2) <= VNStageIntLLROutputS6xD(153)(0);
  CNStageIntLLRInputS7xD(78)(2) <= VNStageIntLLROutputS6xD(153)(1);
  CNStageIntLLRInputS7xD(155)(2) <= VNStageIntLLROutputS6xD(153)(2);
  CNStageIntLLRInputS7xD(203)(2) <= VNStageIntLLROutputS6xD(153)(3);
  CNStageIntLLRInputS7xD(262)(2) <= VNStageIntLLROutputS6xD(153)(4);
  CNStageIntLLRInputS7xD(296)(2) <= VNStageIntLLROutputS6xD(153)(5);
  CNStageIntLLRInputS7xD(376)(2) <= VNStageIntLLROutputS6xD(153)(6);
  CNStageIntLLRInputS7xD(28)(2) <= VNStageIntLLROutputS6xD(154)(0);
  CNStageIntLLRInputS7xD(139)(2) <= VNStageIntLLROutputS6xD(154)(1);
  CNStageIntLLRInputS7xD(183)(2) <= VNStageIntLLROutputS6xD(154)(2);
  CNStageIntLLRInputS7xD(246)(2) <= VNStageIntLLROutputS6xD(154)(3);
  CNStageIntLLRInputS7xD(322)(2) <= VNStageIntLLROutputS6xD(154)(4);
  CNStageIntLLRInputS7xD(27)(2) <= VNStageIntLLROutputS6xD(155)(0);
  CNStageIntLLRInputS7xD(84)(2) <= VNStageIntLLROutputS6xD(155)(1);
  CNStageIntLLRInputS7xD(167)(2) <= VNStageIntLLROutputS6xD(155)(2);
  CNStageIntLLRInputS7xD(174)(2) <= VNStageIntLLROutputS6xD(155)(3);
  CNStageIntLLRInputS7xD(257)(2) <= VNStageIntLLROutputS6xD(155)(4);
  CNStageIntLLRInputS7xD(306)(2) <= VNStageIntLLROutputS6xD(155)(5);
  CNStageIntLLRInputS7xD(357)(2) <= VNStageIntLLROutputS6xD(155)(6);
  CNStageIntLLRInputS7xD(26)(2) <= VNStageIntLLROutputS6xD(156)(0);
  CNStageIntLLRInputS7xD(95)(2) <= VNStageIntLLROutputS6xD(156)(1);
  CNStageIntLLRInputS7xD(157)(2) <= VNStageIntLLROutputS6xD(156)(2);
  CNStageIntLLRInputS7xD(343)(2) <= VNStageIntLLROutputS6xD(156)(3);
  CNStageIntLLRInputS7xD(25)(2) <= VNStageIntLLROutputS6xD(157)(0);
  CNStageIntLLRInputS7xD(102)(2) <= VNStageIntLLROutputS6xD(157)(1);
  CNStageIntLLRInputS7xD(144)(2) <= VNStageIntLLROutputS6xD(157)(2);
  CNStageIntLLRInputS7xD(194)(2) <= VNStageIntLLROutputS6xD(157)(3);
  CNStageIntLLRInputS7xD(323)(2) <= VNStageIntLLROutputS6xD(157)(4);
  CNStageIntLLRInputS7xD(377)(2) <= VNStageIntLLROutputS6xD(157)(5);
  CNStageIntLLRInputS7xD(24)(2) <= VNStageIntLLROutputS6xD(158)(0);
  CNStageIntLLRInputS7xD(77)(2) <= VNStageIntLLROutputS6xD(158)(1);
  CNStageIntLLRInputS7xD(163)(2) <= VNStageIntLLROutputS6xD(158)(2);
  CNStageIntLLRInputS7xD(224)(2) <= VNStageIntLLROutputS6xD(158)(3);
  CNStageIntLLRInputS7xD(230)(2) <= VNStageIntLLROutputS6xD(158)(4);
  CNStageIntLLRInputS7xD(310)(2) <= VNStageIntLLROutputS6xD(158)(5);
  CNStageIntLLRInputS7xD(339)(2) <= VNStageIntLLROutputS6xD(158)(6);
  CNStageIntLLRInputS7xD(23)(2) <= VNStageIntLLROutputS6xD(159)(0);
  CNStageIntLLRInputS7xD(91)(2) <= VNStageIntLLROutputS6xD(159)(1);
  CNStageIntLLRInputS7xD(136)(2) <= VNStageIntLLROutputS6xD(159)(2);
  CNStageIntLLRInputS7xD(271)(2) <= VNStageIntLLROutputS6xD(159)(3);
  CNStageIntLLRInputS7xD(367)(2) <= VNStageIntLLROutputS6xD(159)(4);
  CNStageIntLLRInputS7xD(22)(2) <= VNStageIntLLROutputS6xD(160)(0);
  CNStageIntLLRInputS7xD(62)(2) <= VNStageIntLLROutputS6xD(160)(1);
  CNStageIntLLRInputS7xD(133)(2) <= VNStageIntLLROutputS6xD(160)(2);
  CNStageIntLLRInputS7xD(189)(2) <= VNStageIntLLROutputS6xD(160)(3);
  CNStageIntLLRInputS7xD(233)(2) <= VNStageIntLLROutputS6xD(160)(4);
  CNStageIntLLRInputS7xD(302)(2) <= VNStageIntLLROutputS6xD(160)(5);
  CNStageIntLLRInputS7xD(351)(2) <= VNStageIntLLROutputS6xD(160)(6);
  CNStageIntLLRInputS7xD(21)(2) <= VNStageIntLLROutputS6xD(161)(0);
  CNStageIntLLRInputS7xD(97)(2) <= VNStageIntLLROutputS6xD(161)(1);
  CNStageIntLLRInputS7xD(149)(2) <= VNStageIntLLROutputS6xD(161)(2);
  CNStageIntLLRInputS7xD(171)(2) <= VNStageIntLLROutputS6xD(161)(3);
  CNStageIntLLRInputS7xD(250)(2) <= VNStageIntLLROutputS6xD(161)(4);
  CNStageIntLLRInputS7xD(300)(2) <= VNStageIntLLROutputS6xD(161)(5);
  CNStageIntLLRInputS7xD(379)(2) <= VNStageIntLLROutputS6xD(161)(6);
  CNStageIntLLRInputS7xD(20)(2) <= VNStageIntLLROutputS6xD(162)(0);
  CNStageIntLLRInputS7xD(64)(2) <= VNStageIntLLROutputS6xD(162)(1);
  CNStageIntLLRInputS7xD(141)(2) <= VNStageIntLLROutputS6xD(162)(2);
  CNStageIntLLRInputS7xD(179)(2) <= VNStageIntLLROutputS6xD(162)(3);
  CNStageIntLLRInputS7xD(259)(2) <= VNStageIntLLROutputS6xD(162)(4);
  CNStageIntLLRInputS7xD(315)(2) <= VNStageIntLLROutputS6xD(162)(5);
  CNStageIntLLRInputS7xD(369)(2) <= VNStageIntLLROutputS6xD(162)(6);
  CNStageIntLLRInputS7xD(19)(2) <= VNStageIntLLROutputS6xD(163)(0);
  CNStageIntLLRInputS7xD(79)(2) <= VNStageIntLLROutputS6xD(163)(1);
  CNStageIntLLRInputS7xD(115)(2) <= VNStageIntLLROutputS6xD(163)(2);
  CNStageIntLLRInputS7xD(254)(2) <= VNStageIntLLROutputS6xD(163)(3);
  CNStageIntLLRInputS7xD(355)(2) <= VNStageIntLLROutputS6xD(163)(4);
  CNStageIntLLRInputS7xD(18)(2) <= VNStageIntLLROutputS6xD(164)(0);
  CNStageIntLLRInputS7xD(75)(2) <= VNStageIntLLROutputS6xD(164)(1);
  CNStageIntLLRInputS7xD(125)(2) <= VNStageIntLLROutputS6xD(164)(2);
  CNStageIntLLRInputS7xD(197)(2) <= VNStageIntLLROutputS6xD(164)(3);
  CNStageIntLLRInputS7xD(260)(2) <= VNStageIntLLROutputS6xD(164)(4);
  CNStageIntLLRInputS7xD(375)(2) <= VNStageIntLLROutputS6xD(164)(5);
  CNStageIntLLRInputS7xD(17)(2) <= VNStageIntLLROutputS6xD(165)(0);
  CNStageIntLLRInputS7xD(93)(2) <= VNStageIntLLROutputS6xD(165)(1);
  CNStageIntLLRInputS7xD(119)(2) <= VNStageIntLLROutputS6xD(165)(2);
  CNStageIntLLRInputS7xD(177)(2) <= VNStageIntLLROutputS6xD(165)(3);
  CNStageIntLLRInputS7xD(294)(2) <= VNStageIntLLROutputS6xD(165)(4);
  CNStageIntLLRInputS7xD(348)(2) <= VNStageIntLLROutputS6xD(165)(5);
  CNStageIntLLRInputS7xD(16)(2) <= VNStageIntLLROutputS6xD(166)(0);
  CNStageIntLLRInputS7xD(57)(2) <= VNStageIntLLROutputS6xD(166)(1);
  CNStageIntLLRInputS7xD(122)(2) <= VNStageIntLLROutputS6xD(166)(2);
  CNStageIntLLRInputS7xD(210)(2) <= VNStageIntLLROutputS6xD(166)(3);
  CNStageIntLLRInputS7xD(288)(2) <= VNStageIntLLROutputS6xD(166)(4);
  CNStageIntLLRInputS7xD(345)(2) <= VNStageIntLLROutputS6xD(166)(5);
  CNStageIntLLRInputS7xD(15)(2) <= VNStageIntLLROutputS6xD(167)(0);
  CNStageIntLLRInputS7xD(58)(2) <= VNStageIntLLROutputS6xD(167)(1);
  CNStageIntLLRInputS7xD(112)(2) <= VNStageIntLLROutputS6xD(167)(2);
  CNStageIntLLRInputS7xD(213)(2) <= VNStageIntLLROutputS6xD(167)(3);
  CNStageIntLLRInputS7xD(225)(2) <= VNStageIntLLROutputS6xD(167)(4);
  CNStageIntLLRInputS7xD(292)(2) <= VNStageIntLLROutputS6xD(167)(5);
  CNStageIntLLRInputS7xD(360)(2) <= VNStageIntLLROutputS6xD(167)(6);
  CNStageIntLLRInputS7xD(14)(2) <= VNStageIntLLROutputS6xD(168)(0);
  CNStageIntLLRInputS7xD(150)(2) <= VNStageIntLLROutputS6xD(168)(1);
  CNStageIntLLRInputS7xD(199)(2) <= VNStageIntLLROutputS6xD(168)(2);
  CNStageIntLLRInputS7xD(264)(2) <= VNStageIntLLROutputS6xD(168)(3);
  CNStageIntLLRInputS7xD(283)(2) <= VNStageIntLLROutputS6xD(168)(4);
  CNStageIntLLRInputS7xD(353)(2) <= VNStageIntLLROutputS6xD(168)(5);
  CNStageIntLLRInputS7xD(13)(2) <= VNStageIntLLROutputS6xD(169)(0);
  CNStageIntLLRInputS7xD(85)(2) <= VNStageIntLLROutputS6xD(169)(1);
  CNStageIntLLRInputS7xD(132)(2) <= VNStageIntLLROutputS6xD(169)(2);
  CNStageIntLLRInputS7xD(178)(2) <= VNStageIntLLROutputS6xD(169)(3);
  CNStageIntLLRInputS7xD(266)(2) <= VNStageIntLLROutputS6xD(169)(4);
  CNStageIntLLRInputS7xD(316)(2) <= VNStageIntLLROutputS6xD(169)(5);
  CNStageIntLLRInputS7xD(12)(2) <= VNStageIntLLROutputS6xD(170)(0);
  CNStageIntLLRInputS7xD(101)(2) <= VNStageIntLLROutputS6xD(170)(1);
  CNStageIntLLRInputS7xD(145)(2) <= VNStageIntLLROutputS6xD(170)(2);
  CNStageIntLLRInputS7xD(236)(2) <= VNStageIntLLROutputS6xD(170)(3);
  CNStageIntLLRInputS7xD(337)(2) <= VNStageIntLLROutputS6xD(170)(4);
  CNStageIntLLRInputS7xD(105)(2) <= VNStageIntLLROutputS6xD(171)(0);
  CNStageIntLLRInputS7xD(156)(2) <= VNStageIntLLROutputS6xD(171)(1);
  CNStageIntLLRInputS7xD(222)(2) <= VNStageIntLLROutputS6xD(171)(2);
  CNStageIntLLRInputS7xD(311)(2) <= VNStageIntLLROutputS6xD(171)(3);
  CNStageIntLLRInputS7xD(11)(2) <= VNStageIntLLROutputS6xD(172)(0);
  CNStageIntLLRInputS7xD(110)(2) <= VNStageIntLLROutputS6xD(172)(1);
  CNStageIntLLRInputS7xD(126)(2) <= VNStageIntLLROutputS6xD(172)(2);
  CNStageIntLLRInputS7xD(229)(2) <= VNStageIntLLROutputS6xD(172)(3);
  CNStageIntLLRInputS7xD(10)(2) <= VNStageIntLLROutputS6xD(173)(0);
  CNStageIntLLRInputS7xD(104)(2) <= VNStageIntLLROutputS6xD(173)(1);
  CNStageIntLLRInputS7xD(114)(2) <= VNStageIntLLROutputS6xD(173)(2);
  CNStageIntLLRInputS7xD(180)(2) <= VNStageIntLLROutputS6xD(173)(3);
  CNStageIntLLRInputS7xD(237)(2) <= VNStageIntLLROutputS6xD(173)(4);
  CNStageIntLLRInputS7xD(295)(2) <= VNStageIntLLROutputS6xD(173)(5);
  CNStageIntLLRInputS7xD(9)(2) <= VNStageIntLLROutputS6xD(174)(0);
  CNStageIntLLRInputS7xD(99)(2) <= VNStageIntLLROutputS6xD(174)(1);
  CNStageIntLLRInputS7xD(159)(2) <= VNStageIntLLROutputS6xD(174)(2);
  CNStageIntLLRInputS7xD(265)(2) <= VNStageIntLLROutputS6xD(174)(3);
  CNStageIntLLRInputS7xD(361)(2) <= VNStageIntLLROutputS6xD(174)(4);
  CNStageIntLLRInputS7xD(8)(2) <= VNStageIntLLROutputS6xD(175)(0);
  CNStageIntLLRInputS7xD(82)(2) <= VNStageIntLLROutputS6xD(175)(1);
  CNStageIntLLRInputS7xD(117)(2) <= VNStageIntLLROutputS6xD(175)(2);
  CNStageIntLLRInputS7xD(211)(2) <= VNStageIntLLROutputS6xD(175)(3);
  CNStageIntLLRInputS7xD(278)(2) <= VNStageIntLLROutputS6xD(175)(4);
  CNStageIntLLRInputS7xD(325)(2) <= VNStageIntLLROutputS6xD(175)(5);
  CNStageIntLLRInputS7xD(344)(2) <= VNStageIntLLROutputS6xD(175)(6);
  CNStageIntLLRInputS7xD(7)(2) <= VNStageIntLLROutputS6xD(176)(0);
  CNStageIntLLRInputS7xD(89)(2) <= VNStageIntLLROutputS6xD(176)(1);
  CNStageIntLLRInputS7xD(137)(2) <= VNStageIntLLROutputS6xD(176)(2);
  CNStageIntLLRInputS7xD(176)(2) <= VNStageIntLLROutputS6xD(176)(3);
  CNStageIntLLRInputS7xD(251)(2) <= VNStageIntLLROutputS6xD(176)(4);
  CNStageIntLLRInputS7xD(286)(2) <= VNStageIntLLROutputS6xD(176)(5);
  CNStageIntLLRInputS7xD(356)(2) <= VNStageIntLLROutputS6xD(176)(6);
  CNStageIntLLRInputS7xD(6)(2) <= VNStageIntLLROutputS6xD(177)(0);
  CNStageIntLLRInputS7xD(109)(2) <= VNStageIntLLROutputS6xD(177)(1);
  CNStageIntLLRInputS7xD(147)(2) <= VNStageIntLLROutputS6xD(177)(2);
  CNStageIntLLRInputS7xD(204)(2) <= VNStageIntLLROutputS6xD(177)(3);
  CNStageIntLLRInputS7xD(232)(2) <= VNStageIntLLROutputS6xD(177)(4);
  CNStageIntLLRInputS7xD(304)(2) <= VNStageIntLLROutputS6xD(177)(5);
  CNStageIntLLRInputS7xD(368)(2) <= VNStageIntLLROutputS6xD(177)(6);
  CNStageIntLLRInputS7xD(5)(2) <= VNStageIntLLROutputS6xD(178)(0);
  CNStageIntLLRInputS7xD(107)(2) <= VNStageIntLLROutputS6xD(178)(1);
  CNStageIntLLRInputS7xD(142)(2) <= VNStageIntLLROutputS6xD(178)(2);
  CNStageIntLLRInputS7xD(201)(2) <= VNStageIntLLROutputS6xD(178)(3);
  CNStageIntLLRInputS7xD(313)(2) <= VNStageIntLLROutputS6xD(178)(4);
  CNStageIntLLRInputS7xD(338)(2) <= VNStageIntLLROutputS6xD(178)(5);
  CNStageIntLLRInputS7xD(4)(2) <= VNStageIntLLROutputS6xD(179)(0);
  CNStageIntLLRInputS7xD(87)(2) <= VNStageIntLLROutputS6xD(179)(1);
  CNStageIntLLRInputS7xD(148)(2) <= VNStageIntLLROutputS6xD(179)(2);
  CNStageIntLLRInputS7xD(215)(2) <= VNStageIntLLROutputS6xD(179)(3);
  CNStageIntLLRInputS7xD(267)(2) <= VNStageIntLLROutputS6xD(179)(4);
  CNStageIntLLRInputS7xD(308)(2) <= VNStageIntLLROutputS6xD(179)(5);
  CNStageIntLLRInputS7xD(67)(2) <= VNStageIntLLROutputS6xD(180)(0);
  CNStageIntLLRInputS7xD(208)(2) <= VNStageIntLLROutputS6xD(180)(1);
  CNStageIntLLRInputS7xD(263)(2) <= VNStageIntLLROutputS6xD(180)(2);
  CNStageIntLLRInputS7xD(314)(2) <= VNStageIntLLROutputS6xD(180)(3);
  CNStageIntLLRInputS7xD(371)(2) <= VNStageIntLLROutputS6xD(180)(4);
  CNStageIntLLRInputS7xD(3)(2) <= VNStageIntLLROutputS6xD(181)(0);
  CNStageIntLLRInputS7xD(70)(2) <= VNStageIntLLROutputS6xD(181)(1);
  CNStageIntLLRInputS7xD(162)(2) <= VNStageIntLLROutputS6xD(181)(2);
  CNStageIntLLRInputS7xD(186)(2) <= VNStageIntLLROutputS6xD(181)(3);
  CNStageIntLLRInputS7xD(227)(2) <= VNStageIntLLROutputS6xD(181)(4);
  CNStageIntLLRInputS7xD(303)(2) <= VNStageIntLLROutputS6xD(181)(5);
  CNStageIntLLRInputS7xD(2)(2) <= VNStageIntLLROutputS6xD(182)(0);
  CNStageIntLLRInputS7xD(54)(2) <= VNStageIntLLROutputS6xD(182)(1);
  CNStageIntLLRInputS7xD(169)(2) <= VNStageIntLLROutputS6xD(182)(2);
  CNStageIntLLRInputS7xD(195)(2) <= VNStageIntLLROutputS6xD(182)(3);
  CNStageIntLLRInputS7xD(248)(2) <= VNStageIntLLROutputS6xD(182)(4);
  CNStageIntLLRInputS7xD(328)(2) <= VNStageIntLLROutputS6xD(182)(5);
  CNStageIntLLRInputS7xD(350)(2) <= VNStageIntLLROutputS6xD(182)(6);
  CNStageIntLLRInputS7xD(1)(2) <= VNStageIntLLROutputS6xD(183)(0);
  CNStageIntLLRInputS7xD(88)(2) <= VNStageIntLLROutputS6xD(183)(1);
  CNStageIntLLRInputS7xD(190)(2) <= VNStageIntLLROutputS6xD(183)(2);
  CNStageIntLLRInputS7xD(281)(2) <= VNStageIntLLROutputS6xD(183)(3);
  CNStageIntLLRInputS7xD(358)(2) <= VNStageIntLLROutputS6xD(183)(4);
  CNStageIntLLRInputS7xD(0)(2) <= VNStageIntLLROutputS6xD(184)(0);
  CNStageIntLLRInputS7xD(106)(2) <= VNStageIntLLROutputS6xD(184)(1);
  CNStageIntLLRInputS7xD(153)(2) <= VNStageIntLLROutputS6xD(184)(2);
  CNStageIntLLRInputS7xD(193)(2) <= VNStageIntLLROutputS6xD(184)(3);
  CNStageIntLLRInputS7xD(226)(2) <= VNStageIntLLROutputS6xD(184)(4);
  CNStageIntLLRInputS7xD(318)(2) <= VNStageIntLLROutputS6xD(184)(5);
  CNStageIntLLRInputS7xD(354)(2) <= VNStageIntLLROutputS6xD(184)(6);
  CNStageIntLLRInputS7xD(121)(2) <= VNStageIntLLROutputS6xD(185)(0);
  CNStageIntLLRInputS7xD(272)(2) <= VNStageIntLLROutputS6xD(185)(1);
  CNStageIntLLRInputS7xD(320)(2) <= VNStageIntLLROutputS6xD(185)(2);
  CNStageIntLLRInputS7xD(359)(2) <= VNStageIntLLROutputS6xD(185)(3);
  CNStageIntLLRInputS7xD(63)(2) <= VNStageIntLLROutputS6xD(186)(0);
  CNStageIntLLRInputS7xD(160)(2) <= VNStageIntLLROutputS6xD(186)(1);
  CNStageIntLLRInputS7xD(216)(2) <= VNStageIntLLROutputS6xD(186)(2);
  CNStageIntLLRInputS7xD(235)(2) <= VNStageIntLLROutputS6xD(186)(3);
  CNStageIntLLRInputS7xD(290)(2) <= VNStageIntLLROutputS6xD(186)(4);
  CNStageIntLLRInputS7xD(349)(2) <= VNStageIntLLROutputS6xD(186)(5);
  CNStageIntLLRInputS7xD(90)(2) <= VNStageIntLLROutputS6xD(187)(0);
  CNStageIntLLRInputS7xD(113)(2) <= VNStageIntLLROutputS6xD(187)(1);
  CNStageIntLLRInputS7xD(200)(2) <= VNStageIntLLROutputS6xD(187)(2);
  CNStageIntLLRInputS7xD(240)(2) <= VNStageIntLLROutputS6xD(187)(3);
  CNStageIntLLRInputS7xD(326)(2) <= VNStageIntLLROutputS6xD(187)(4);
  CNStageIntLLRInputS7xD(374)(2) <= VNStageIntLLROutputS6xD(187)(5);
  CNStageIntLLRInputS7xD(81)(2) <= VNStageIntLLROutputS6xD(188)(0);
  CNStageIntLLRInputS7xD(212)(2) <= VNStageIntLLROutputS6xD(188)(1);
  CNStageIntLLRInputS7xD(279)(2) <= VNStageIntLLROutputS6xD(188)(2);
  CNStageIntLLRInputS7xD(284)(2) <= VNStageIntLLROutputS6xD(188)(3);
  CNStageIntLLRInputS7xD(381)(2) <= VNStageIntLLROutputS6xD(188)(4);
  CNStageIntLLRInputS7xD(68)(2) <= VNStageIntLLROutputS6xD(189)(0);
  CNStageIntLLRInputS7xD(152)(2) <= VNStageIntLLROutputS6xD(189)(1);
  CNStageIntLLRInputS7xD(223)(2) <= VNStageIntLLROutputS6xD(189)(2);
  CNStageIntLLRInputS7xD(239)(2) <= VNStageIntLLROutputS6xD(189)(3);
  CNStageIntLLRInputS7xD(291)(2) <= VNStageIntLLROutputS6xD(189)(4);
  CNStageIntLLRInputS7xD(363)(2) <= VNStageIntLLROutputS6xD(189)(5);
  CNStageIntLLRInputS7xD(168)(2) <= VNStageIntLLROutputS6xD(190)(0);
  CNStageIntLLRInputS7xD(196)(2) <= VNStageIntLLROutputS6xD(190)(1);
  CNStageIntLLRInputS7xD(234)(2) <= VNStageIntLLROutputS6xD(190)(2);
  CNStageIntLLRInputS7xD(319)(2) <= VNStageIntLLROutputS6xD(190)(3);
  CNStageIntLLRInputS7xD(365)(2) <= VNStageIntLLROutputS6xD(190)(4);
  CNStageIntLLRInputS7xD(52)(2) <= VNStageIntLLROutputS6xD(191)(0);
  CNStageIntLLRInputS7xD(59)(2) <= VNStageIntLLROutputS6xD(191)(1);
  CNStageIntLLRInputS7xD(138)(2) <= VNStageIntLLROutputS6xD(191)(2);
  CNStageIntLLRInputS7xD(185)(2) <= VNStageIntLLROutputS6xD(191)(3);
  CNStageIntLLRInputS7xD(270)(2) <= VNStageIntLLROutputS6xD(191)(4);
  CNStageIntLLRInputS7xD(280)(2) <= VNStageIntLLROutputS6xD(191)(5);
  CNStageIntLLRInputS7xD(53)(3) <= VNStageIntLLROutputS6xD(192)(0);
  CNStageIntLLRInputS7xD(107)(3) <= VNStageIntLLROutputS6xD(192)(1);
  CNStageIntLLRInputS7xD(128)(3) <= VNStageIntLLROutputS6xD(192)(2);
  CNStageIntLLRInputS7xD(197)(3) <= VNStageIntLLROutputS6xD(192)(3);
  CNStageIntLLRInputS7xD(243)(3) <= VNStageIntLLROutputS6xD(192)(4);
  CNStageIntLLRInputS7xD(297)(3) <= VNStageIntLLROutputS6xD(192)(5);
  CNStageIntLLRInputS7xD(340)(3) <= VNStageIntLLROutputS6xD(192)(6);
  CNStageIntLLRInputS7xD(51)(3) <= VNStageIntLLROutputS6xD(193)(0);
  CNStageIntLLRInputS7xD(58)(3) <= VNStageIntLLROutputS6xD(193)(1);
  CNStageIntLLRInputS7xD(137)(3) <= VNStageIntLLROutputS6xD(193)(2);
  CNStageIntLLRInputS7xD(269)(3) <= VNStageIntLLROutputS6xD(193)(3);
  CNStageIntLLRInputS7xD(333)(3) <= VNStageIntLLROutputS6xD(193)(4);
  CNStageIntLLRInputS7xD(50)(3) <= VNStageIntLLROutputS6xD(194)(0);
  CNStageIntLLRInputS7xD(55)(3) <= VNStageIntLLROutputS6xD(194)(1);
  CNStageIntLLRInputS7xD(115)(3) <= VNStageIntLLROutputS6xD(194)(2);
  CNStageIntLLRInputS7xD(171)(3) <= VNStageIntLLROutputS6xD(194)(3);
  CNStageIntLLRInputS7xD(275)(3) <= VNStageIntLLROutputS6xD(194)(4);
  CNStageIntLLRInputS7xD(304)(3) <= VNStageIntLLROutputS6xD(194)(5);
  CNStageIntLLRInputS7xD(371)(3) <= VNStageIntLLROutputS6xD(194)(6);
  CNStageIntLLRInputS7xD(72)(3) <= VNStageIntLLROutputS6xD(195)(0);
  CNStageIntLLRInputS7xD(139)(3) <= VNStageIntLLROutputS6xD(195)(1);
  CNStageIntLLRInputS7xD(187)(3) <= VNStageIntLLROutputS6xD(195)(2);
  CNStageIntLLRInputS7xD(244)(3) <= VNStageIntLLROutputS6xD(195)(3);
  CNStageIntLLRInputS7xD(49)(3) <= VNStageIntLLROutputS6xD(196)(0);
  CNStageIntLLRInputS7xD(64)(3) <= VNStageIntLLROutputS6xD(196)(1);
  CNStageIntLLRInputS7xD(153)(3) <= VNStageIntLLROutputS6xD(196)(2);
  CNStageIntLLRInputS7xD(205)(3) <= VNStageIntLLROutputS6xD(196)(3);
  CNStageIntLLRInputS7xD(242)(3) <= VNStageIntLLROutputS6xD(196)(4);
  CNStageIntLLRInputS7xD(306)(3) <= VNStageIntLLROutputS6xD(196)(5);
  CNStageIntLLRInputS7xD(48)(3) <= VNStageIntLLROutputS6xD(197)(0);
  CNStageIntLLRInputS7xD(96)(3) <= VNStageIntLLROutputS6xD(197)(1);
  CNStageIntLLRInputS7xD(150)(3) <= VNStageIntLLROutputS6xD(197)(2);
  CNStageIntLLRInputS7xD(213)(3) <= VNStageIntLLROutputS6xD(197)(3);
  CNStageIntLLRInputS7xD(273)(3) <= VNStageIntLLROutputS6xD(197)(4);
  CNStageIntLLRInputS7xD(320)(3) <= VNStageIntLLROutputS6xD(197)(5);
  CNStageIntLLRInputS7xD(363)(3) <= VNStageIntLLROutputS6xD(197)(6);
  CNStageIntLLRInputS7xD(47)(3) <= VNStageIntLLROutputS6xD(198)(0);
  CNStageIntLLRInputS7xD(105)(3) <= VNStageIntLLROutputS6xD(198)(1);
  CNStageIntLLRInputS7xD(111)(3) <= VNStageIntLLROutputS6xD(198)(2);
  CNStageIntLLRInputS7xD(208)(3) <= VNStageIntLLROutputS6xD(198)(3);
  CNStageIntLLRInputS7xD(254)(3) <= VNStageIntLLROutputS6xD(198)(4);
  CNStageIntLLRInputS7xD(316)(3) <= VNStageIntLLROutputS6xD(198)(5);
  CNStageIntLLRInputS7xD(379)(3) <= VNStageIntLLROutputS6xD(198)(6);
  CNStageIntLLRInputS7xD(46)(3) <= VNStageIntLLROutputS6xD(199)(0);
  CNStageIntLLRInputS7xD(99)(3) <= VNStageIntLLROutputS6xD(199)(1);
  CNStageIntLLRInputS7xD(133)(3) <= VNStageIntLLROutputS6xD(199)(2);
  CNStageIntLLRInputS7xD(214)(3) <= VNStageIntLLROutputS6xD(199)(3);
  CNStageIntLLRInputS7xD(257)(3) <= VNStageIntLLROutputS6xD(199)(4);
  CNStageIntLLRInputS7xD(282)(3) <= VNStageIntLLROutputS6xD(199)(5);
  CNStageIntLLRInputS7xD(350)(3) <= VNStageIntLLROutputS6xD(199)(6);
  CNStageIntLLRInputS7xD(45)(3) <= VNStageIntLLROutputS6xD(200)(0);
  CNStageIntLLRInputS7xD(102)(3) <= VNStageIntLLROutputS6xD(200)(1);
  CNStageIntLLRInputS7xD(134)(3) <= VNStageIntLLROutputS6xD(200)(2);
  CNStageIntLLRInputS7xD(204)(3) <= VNStageIntLLROutputS6xD(200)(3);
  CNStageIntLLRInputS7xD(245)(3) <= VNStageIntLLROutputS6xD(200)(4);
  CNStageIntLLRInputS7xD(300)(3) <= VNStageIntLLROutputS6xD(200)(5);
  CNStageIntLLRInputS7xD(44)(3) <= VNStageIntLLROutputS6xD(201)(0);
  CNStageIntLLRInputS7xD(93)(3) <= VNStageIntLLROutputS6xD(201)(1);
  CNStageIntLLRInputS7xD(169)(3) <= VNStageIntLLROutputS6xD(201)(2);
  CNStageIntLLRInputS7xD(174)(3) <= VNStageIntLLROutputS6xD(201)(3);
  CNStageIntLLRInputS7xD(274)(3) <= VNStageIntLLROutputS6xD(201)(4);
  CNStageIntLLRInputS7xD(351)(3) <= VNStageIntLLROutputS6xD(201)(5);
  CNStageIntLLRInputS7xD(43)(3) <= VNStageIntLLROutputS6xD(202)(0);
  CNStageIntLLRInputS7xD(73)(3) <= VNStageIntLLROutputS6xD(202)(1);
  CNStageIntLLRInputS7xD(160)(3) <= VNStageIntLLROutputS6xD(202)(2);
  CNStageIntLLRInputS7xD(181)(3) <= VNStageIntLLROutputS6xD(202)(3);
  CNStageIntLLRInputS7xD(281)(3) <= VNStageIntLLROutputS6xD(202)(4);
  CNStageIntLLRInputS7xD(365)(3) <= VNStageIntLLROutputS6xD(202)(5);
  CNStageIntLLRInputS7xD(42)(3) <= VNStageIntLLROutputS6xD(203)(0);
  CNStageIntLLRInputS7xD(54)(3) <= VNStageIntLLROutputS6xD(203)(1);
  CNStageIntLLRInputS7xD(119)(3) <= VNStageIntLLROutputS6xD(203)(2);
  CNStageIntLLRInputS7xD(217)(3) <= VNStageIntLLROutputS6xD(203)(3);
  CNStageIntLLRInputS7xD(267)(3) <= VNStageIntLLROutputS6xD(203)(4);
  CNStageIntLLRInputS7xD(326)(3) <= VNStageIntLLROutputS6xD(203)(5);
  CNStageIntLLRInputS7xD(361)(3) <= VNStageIntLLROutputS6xD(203)(6);
  CNStageIntLLRInputS7xD(41)(3) <= VNStageIntLLROutputS6xD(204)(0);
  CNStageIntLLRInputS7xD(68)(3) <= VNStageIntLLROutputS6xD(204)(1);
  CNStageIntLLRInputS7xD(123)(3) <= VNStageIntLLROutputS6xD(204)(2);
  CNStageIntLLRInputS7xD(219)(3) <= VNStageIntLLROutputS6xD(204)(3);
  CNStageIntLLRInputS7xD(251)(3) <= VNStageIntLLROutputS6xD(204)(4);
  CNStageIntLLRInputS7xD(288)(3) <= VNStageIntLLROutputS6xD(204)(5);
  CNStageIntLLRInputS7xD(382)(3) <= VNStageIntLLROutputS6xD(204)(6);
  CNStageIntLLRInputS7xD(170)(3) <= VNStageIntLLROutputS6xD(205)(0);
  CNStageIntLLRInputS7xD(276)(3) <= VNStageIntLLROutputS6xD(205)(1);
  CNStageIntLLRInputS7xD(345)(3) <= VNStageIntLLROutputS6xD(205)(2);
  CNStageIntLLRInputS7xD(40)(3) <= VNStageIntLLROutputS6xD(206)(0);
  CNStageIntLLRInputS7xD(122)(3) <= VNStageIntLLROutputS6xD(206)(1);
  CNStageIntLLRInputS7xD(172)(3) <= VNStageIntLLROutputS6xD(206)(2);
  CNStageIntLLRInputS7xD(332)(3) <= VNStageIntLLROutputS6xD(206)(3);
  CNStageIntLLRInputS7xD(346)(3) <= VNStageIntLLROutputS6xD(206)(4);
  CNStageIntLLRInputS7xD(39)(3) <= VNStageIntLLROutputS6xD(207)(0);
  CNStageIntLLRInputS7xD(95)(3) <= VNStageIntLLROutputS6xD(207)(1);
  CNStageIntLLRInputS7xD(117)(3) <= VNStageIntLLROutputS6xD(207)(2);
  CNStageIntLLRInputS7xD(255)(3) <= VNStageIntLLROutputS6xD(207)(3);
  CNStageIntLLRInputS7xD(292)(3) <= VNStageIntLLROutputS6xD(207)(4);
  CNStageIntLLRInputS7xD(381)(3) <= VNStageIntLLROutputS6xD(207)(5);
  CNStageIntLLRInputS7xD(38)(3) <= VNStageIntLLROutputS6xD(208)(0);
  CNStageIntLLRInputS7xD(82)(3) <= VNStageIntLLROutputS6xD(208)(1);
  CNStageIntLLRInputS7xD(157)(3) <= VNStageIntLLROutputS6xD(208)(2);
  CNStageIntLLRInputS7xD(191)(3) <= VNStageIntLLROutputS6xD(208)(3);
  CNStageIntLLRInputS7xD(286)(3) <= VNStageIntLLROutputS6xD(208)(4);
  CNStageIntLLRInputS7xD(372)(3) <= VNStageIntLLROutputS6xD(208)(5);
  CNStageIntLLRInputS7xD(37)(3) <= VNStageIntLLROutputS6xD(209)(0);
  CNStageIntLLRInputS7xD(97)(3) <= VNStageIntLLROutputS6xD(209)(1);
  CNStageIntLLRInputS7xD(165)(3) <= VNStageIntLLROutputS6xD(209)(2);
  CNStageIntLLRInputS7xD(218)(3) <= VNStageIntLLROutputS6xD(209)(3);
  CNStageIntLLRInputS7xD(323)(3) <= VNStageIntLLROutputS6xD(209)(4);
  CNStageIntLLRInputS7xD(36)(3) <= VNStageIntLLROutputS6xD(210)(0);
  CNStageIntLLRInputS7xD(60)(3) <= VNStageIntLLROutputS6xD(210)(1);
  CNStageIntLLRInputS7xD(129)(3) <= VNStageIntLLROutputS6xD(210)(2);
  CNStageIntLLRInputS7xD(180)(3) <= VNStageIntLLROutputS6xD(210)(3);
  CNStageIntLLRInputS7xD(246)(3) <= VNStageIntLLROutputS6xD(210)(4);
  CNStageIntLLRInputS7xD(330)(3) <= VNStageIntLLROutputS6xD(210)(5);
  CNStageIntLLRInputS7xD(335)(3) <= VNStageIntLLROutputS6xD(210)(6);
  CNStageIntLLRInputS7xD(35)(3) <= VNStageIntLLROutputS6xD(211)(0);
  CNStageIntLLRInputS7xD(70)(3) <= VNStageIntLLROutputS6xD(211)(1);
  CNStageIntLLRInputS7xD(127)(3) <= VNStageIntLLROutputS6xD(211)(2);
  CNStageIntLLRInputS7xD(206)(3) <= VNStageIntLLROutputS6xD(211)(3);
  CNStageIntLLRInputS7xD(260)(3) <= VNStageIntLLROutputS6xD(211)(4);
  CNStageIntLLRInputS7xD(298)(3) <= VNStageIntLLROutputS6xD(211)(5);
  CNStageIntLLRInputS7xD(34)(3) <= VNStageIntLLROutputS6xD(212)(0);
  CNStageIntLLRInputS7xD(65)(3) <= VNStageIntLLROutputS6xD(212)(1);
  CNStageIntLLRInputS7xD(163)(3) <= VNStageIntLLROutputS6xD(212)(2);
  CNStageIntLLRInputS7xD(186)(3) <= VNStageIntLLROutputS6xD(212)(3);
  CNStageIntLLRInputS7xD(296)(3) <= VNStageIntLLROutputS6xD(212)(4);
  CNStageIntLLRInputS7xD(33)(3) <= VNStageIntLLROutputS6xD(213)(0);
  CNStageIntLLRInputS7xD(71)(3) <= VNStageIntLLROutputS6xD(213)(1);
  CNStageIntLLRInputS7xD(142)(3) <= VNStageIntLLROutputS6xD(213)(2);
  CNStageIntLLRInputS7xD(230)(3) <= VNStageIntLLROutputS6xD(213)(3);
  CNStageIntLLRInputS7xD(32)(3) <= VNStageIntLLROutputS6xD(214)(0);
  CNStageIntLLRInputS7xD(59)(3) <= VNStageIntLLROutputS6xD(214)(1);
  CNStageIntLLRInputS7xD(145)(3) <= VNStageIntLLROutputS6xD(214)(2);
  CNStageIntLLRInputS7xD(220)(3) <= VNStageIntLLROutputS6xD(214)(3);
  CNStageIntLLRInputS7xD(240)(3) <= VNStageIntLLROutputS6xD(214)(4);
  CNStageIntLLRInputS7xD(308)(3) <= VNStageIntLLROutputS6xD(214)(5);
  CNStageIntLLRInputS7xD(369)(3) <= VNStageIntLLROutputS6xD(214)(6);
  CNStageIntLLRInputS7xD(31)(3) <= VNStageIntLLROutputS6xD(215)(0);
  CNStageIntLLRInputS7xD(85)(3) <= VNStageIntLLROutputS6xD(215)(1);
  CNStageIntLLRInputS7xD(130)(3) <= VNStageIntLLROutputS6xD(215)(2);
  CNStageIntLLRInputS7xD(216)(3) <= VNStageIntLLROutputS6xD(215)(3);
  CNStageIntLLRInputS7xD(234)(3) <= VNStageIntLLROutputS6xD(215)(4);
  CNStageIntLLRInputS7xD(311)(3) <= VNStageIntLLROutputS6xD(215)(5);
  CNStageIntLLRInputS7xD(377)(3) <= VNStageIntLLROutputS6xD(215)(6);
  CNStageIntLLRInputS7xD(30)(3) <= VNStageIntLLROutputS6xD(216)(0);
  CNStageIntLLRInputS7xD(91)(3) <= VNStageIntLLROutputS6xD(216)(1);
  CNStageIntLLRInputS7xD(164)(3) <= VNStageIntLLROutputS6xD(216)(2);
  CNStageIntLLRInputS7xD(183)(3) <= VNStageIntLLROutputS6xD(216)(3);
  CNStageIntLLRInputS7xD(237)(3) <= VNStageIntLLROutputS6xD(216)(4);
  CNStageIntLLRInputS7xD(299)(3) <= VNStageIntLLROutputS6xD(216)(5);
  CNStageIntLLRInputS7xD(341)(3) <= VNStageIntLLROutputS6xD(216)(6);
  CNStageIntLLRInputS7xD(29)(3) <= VNStageIntLLROutputS6xD(217)(0);
  CNStageIntLLRInputS7xD(75)(3) <= VNStageIntLLROutputS6xD(217)(1);
  CNStageIntLLRInputS7xD(126)(3) <= VNStageIntLLROutputS6xD(217)(2);
  CNStageIntLLRInputS7xD(201)(3) <= VNStageIntLLROutputS6xD(217)(3);
  CNStageIntLLRInputS7xD(227)(3) <= VNStageIntLLROutputS6xD(217)(4);
  CNStageIntLLRInputS7xD(329)(3) <= VNStageIntLLROutputS6xD(217)(5);
  CNStageIntLLRInputS7xD(339)(3) <= VNStageIntLLROutputS6xD(217)(6);
  CNStageIntLLRInputS7xD(28)(3) <= VNStageIntLLROutputS6xD(218)(0);
  CNStageIntLLRInputS7xD(77)(3) <= VNStageIntLLROutputS6xD(218)(1);
  CNStageIntLLRInputS7xD(154)(3) <= VNStageIntLLROutputS6xD(218)(2);
  CNStageIntLLRInputS7xD(202)(3) <= VNStageIntLLROutputS6xD(218)(3);
  CNStageIntLLRInputS7xD(261)(3) <= VNStageIntLLROutputS6xD(218)(4);
  CNStageIntLLRInputS7xD(295)(3) <= VNStageIntLLROutputS6xD(218)(5);
  CNStageIntLLRInputS7xD(375)(3) <= VNStageIntLLROutputS6xD(218)(6);
  CNStageIntLLRInputS7xD(27)(3) <= VNStageIntLLROutputS6xD(219)(0);
  CNStageIntLLRInputS7xD(101)(3) <= VNStageIntLLROutputS6xD(219)(1);
  CNStageIntLLRInputS7xD(138)(3) <= VNStageIntLLROutputS6xD(219)(2);
  CNStageIntLLRInputS7xD(182)(3) <= VNStageIntLLROutputS6xD(219)(3);
  CNStageIntLLRInputS7xD(321)(3) <= VNStageIntLLROutputS6xD(219)(4);
  CNStageIntLLRInputS7xD(354)(3) <= VNStageIntLLROutputS6xD(219)(5);
  CNStageIntLLRInputS7xD(26)(3) <= VNStageIntLLROutputS6xD(220)(0);
  CNStageIntLLRInputS7xD(83)(3) <= VNStageIntLLROutputS6xD(220)(1);
  CNStageIntLLRInputS7xD(166)(3) <= VNStageIntLLROutputS6xD(220)(2);
  CNStageIntLLRInputS7xD(173)(3) <= VNStageIntLLROutputS6xD(220)(3);
  CNStageIntLLRInputS7xD(256)(3) <= VNStageIntLLROutputS6xD(220)(4);
  CNStageIntLLRInputS7xD(305)(3) <= VNStageIntLLROutputS6xD(220)(5);
  CNStageIntLLRInputS7xD(356)(3) <= VNStageIntLLROutputS6xD(220)(6);
  CNStageIntLLRInputS7xD(25)(3) <= VNStageIntLLROutputS6xD(221)(0);
  CNStageIntLLRInputS7xD(94)(3) <= VNStageIntLLROutputS6xD(221)(1);
  CNStageIntLLRInputS7xD(156)(3) <= VNStageIntLLROutputS6xD(221)(2);
  CNStageIntLLRInputS7xD(190)(3) <= VNStageIntLLROutputS6xD(221)(3);
  CNStageIntLLRInputS7xD(268)(3) <= VNStageIntLLROutputS6xD(221)(4);
  CNStageIntLLRInputS7xD(331)(3) <= VNStageIntLLROutputS6xD(221)(5);
  CNStageIntLLRInputS7xD(342)(3) <= VNStageIntLLROutputS6xD(221)(6);
  CNStageIntLLRInputS7xD(24)(3) <= VNStageIntLLROutputS6xD(222)(0);
  CNStageIntLLRInputS7xD(143)(3) <= VNStageIntLLROutputS6xD(222)(1);
  CNStageIntLLRInputS7xD(241)(3) <= VNStageIntLLROutputS6xD(222)(2);
  CNStageIntLLRInputS7xD(376)(3) <= VNStageIntLLROutputS6xD(222)(3);
  CNStageIntLLRInputS7xD(23)(3) <= VNStageIntLLROutputS6xD(223)(0);
  CNStageIntLLRInputS7xD(76)(3) <= VNStageIntLLROutputS6xD(223)(1);
  CNStageIntLLRInputS7xD(162)(3) <= VNStageIntLLROutputS6xD(223)(2);
  CNStageIntLLRInputS7xD(224)(3) <= VNStageIntLLROutputS6xD(223)(3);
  CNStageIntLLRInputS7xD(229)(3) <= VNStageIntLLROutputS6xD(223)(4);
  CNStageIntLLRInputS7xD(309)(3) <= VNStageIntLLROutputS6xD(223)(5);
  CNStageIntLLRInputS7xD(338)(3) <= VNStageIntLLROutputS6xD(223)(6);
  CNStageIntLLRInputS7xD(22)(3) <= VNStageIntLLROutputS6xD(224)(0);
  CNStageIntLLRInputS7xD(90)(3) <= VNStageIntLLROutputS6xD(224)(1);
  CNStageIntLLRInputS7xD(135)(3) <= VNStageIntLLROutputS6xD(224)(2);
  CNStageIntLLRInputS7xD(193)(3) <= VNStageIntLLROutputS6xD(224)(3);
  CNStageIntLLRInputS7xD(270)(3) <= VNStageIntLLROutputS6xD(224)(4);
  CNStageIntLLRInputS7xD(328)(3) <= VNStageIntLLROutputS6xD(224)(5);
  CNStageIntLLRInputS7xD(366)(3) <= VNStageIntLLROutputS6xD(224)(6);
  CNStageIntLLRInputS7xD(21)(3) <= VNStageIntLLROutputS6xD(225)(0);
  CNStageIntLLRInputS7xD(61)(3) <= VNStageIntLLROutputS6xD(225)(1);
  CNStageIntLLRInputS7xD(132)(3) <= VNStageIntLLROutputS6xD(225)(2);
  CNStageIntLLRInputS7xD(188)(3) <= VNStageIntLLROutputS6xD(225)(3);
  CNStageIntLLRInputS7xD(232)(3) <= VNStageIntLLROutputS6xD(225)(4);
  CNStageIntLLRInputS7xD(301)(3) <= VNStageIntLLROutputS6xD(225)(5);
  CNStageIntLLRInputS7xD(20)(3) <= VNStageIntLLROutputS6xD(226)(0);
  CNStageIntLLRInputS7xD(148)(3) <= VNStageIntLLROutputS6xD(226)(1);
  CNStageIntLLRInputS7xD(378)(3) <= VNStageIntLLROutputS6xD(226)(2);
  CNStageIntLLRInputS7xD(19)(3) <= VNStageIntLLROutputS6xD(227)(0);
  CNStageIntLLRInputS7xD(63)(3) <= VNStageIntLLROutputS6xD(227)(1);
  CNStageIntLLRInputS7xD(140)(3) <= VNStageIntLLROutputS6xD(227)(2);
  CNStageIntLLRInputS7xD(178)(3) <= VNStageIntLLROutputS6xD(227)(3);
  CNStageIntLLRInputS7xD(258)(3) <= VNStageIntLLROutputS6xD(227)(4);
  CNStageIntLLRInputS7xD(314)(3) <= VNStageIntLLROutputS6xD(227)(5);
  CNStageIntLLRInputS7xD(368)(3) <= VNStageIntLLROutputS6xD(227)(6);
  CNStageIntLLRInputS7xD(18)(3) <= VNStageIntLLROutputS6xD(228)(0);
  CNStageIntLLRInputS7xD(78)(3) <= VNStageIntLLROutputS6xD(228)(1);
  CNStageIntLLRInputS7xD(114)(3) <= VNStageIntLLROutputS6xD(228)(2);
  CNStageIntLLRInputS7xD(198)(3) <= VNStageIntLLROutputS6xD(228)(3);
  CNStageIntLLRInputS7xD(253)(3) <= VNStageIntLLROutputS6xD(228)(4);
  CNStageIntLLRInputS7xD(307)(3) <= VNStageIntLLROutputS6xD(228)(5);
  CNStageIntLLRInputS7xD(17)(3) <= VNStageIntLLROutputS6xD(229)(0);
  CNStageIntLLRInputS7xD(74)(3) <= VNStageIntLLROutputS6xD(229)(1);
  CNStageIntLLRInputS7xD(124)(3) <= VNStageIntLLROutputS6xD(229)(2);
  CNStageIntLLRInputS7xD(259)(3) <= VNStageIntLLROutputS6xD(229)(3);
  CNStageIntLLRInputS7xD(374)(3) <= VNStageIntLLROutputS6xD(229)(4);
  CNStageIntLLRInputS7xD(16)(3) <= VNStageIntLLROutputS6xD(230)(0);
  CNStageIntLLRInputS7xD(118)(3) <= VNStageIntLLROutputS6xD(230)(1);
  CNStageIntLLRInputS7xD(176)(3) <= VNStageIntLLROutputS6xD(230)(2);
  CNStageIntLLRInputS7xD(249)(3) <= VNStageIntLLROutputS6xD(230)(3);
  CNStageIntLLRInputS7xD(293)(3) <= VNStageIntLLROutputS6xD(230)(4);
  CNStageIntLLRInputS7xD(347)(3) <= VNStageIntLLROutputS6xD(230)(5);
  CNStageIntLLRInputS7xD(15)(3) <= VNStageIntLLROutputS6xD(231)(0);
  CNStageIntLLRInputS7xD(56)(3) <= VNStageIntLLROutputS6xD(231)(1);
  CNStageIntLLRInputS7xD(209)(3) <= VNStageIntLLROutputS6xD(231)(2);
  CNStageIntLLRInputS7xD(272)(3) <= VNStageIntLLROutputS6xD(231)(3);
  CNStageIntLLRInputS7xD(287)(3) <= VNStageIntLLROutputS6xD(231)(4);
  CNStageIntLLRInputS7xD(344)(3) <= VNStageIntLLROutputS6xD(231)(5);
  CNStageIntLLRInputS7xD(14)(3) <= VNStageIntLLROutputS6xD(232)(0);
  CNStageIntLLRInputS7xD(57)(3) <= VNStageIntLLROutputS6xD(232)(1);
  CNStageIntLLRInputS7xD(212)(3) <= VNStageIntLLROutputS6xD(232)(2);
  CNStageIntLLRInputS7xD(278)(3) <= VNStageIntLLROutputS6xD(232)(3);
  CNStageIntLLRInputS7xD(291)(3) <= VNStageIntLLROutputS6xD(232)(4);
  CNStageIntLLRInputS7xD(359)(3) <= VNStageIntLLROutputS6xD(232)(5);
  CNStageIntLLRInputS7xD(13)(3) <= VNStageIntLLROutputS6xD(233)(0);
  CNStageIntLLRInputS7xD(92)(3) <= VNStageIntLLROutputS6xD(233)(1);
  CNStageIntLLRInputS7xD(149)(3) <= VNStageIntLLROutputS6xD(233)(2);
  CNStageIntLLRInputS7xD(263)(3) <= VNStageIntLLROutputS6xD(233)(3);
  CNStageIntLLRInputS7xD(352)(3) <= VNStageIntLLROutputS6xD(233)(4);
  CNStageIntLLRInputS7xD(12)(3) <= VNStageIntLLROutputS6xD(234)(0);
  CNStageIntLLRInputS7xD(84)(3) <= VNStageIntLLROutputS6xD(234)(1);
  CNStageIntLLRInputS7xD(131)(3) <= VNStageIntLLROutputS6xD(234)(2);
  CNStageIntLLRInputS7xD(177)(3) <= VNStageIntLLROutputS6xD(234)(3);
  CNStageIntLLRInputS7xD(265)(3) <= VNStageIntLLROutputS6xD(234)(4);
  CNStageIntLLRInputS7xD(315)(3) <= VNStageIntLLROutputS6xD(234)(5);
  CNStageIntLLRInputS7xD(100)(3) <= VNStageIntLLROutputS6xD(235)(0);
  CNStageIntLLRInputS7xD(144)(3) <= VNStageIntLLROutputS6xD(235)(1);
  CNStageIntLLRInputS7xD(196)(3) <= VNStageIntLLROutputS6xD(235)(2);
  CNStageIntLLRInputS7xD(235)(3) <= VNStageIntLLROutputS6xD(235)(3);
  CNStageIntLLRInputS7xD(336)(3) <= VNStageIntLLROutputS6xD(235)(4);
  CNStageIntLLRInputS7xD(11)(3) <= VNStageIntLLROutputS6xD(236)(0);
  CNStageIntLLRInputS7xD(104)(3) <= VNStageIntLLROutputS6xD(236)(1);
  CNStageIntLLRInputS7xD(155)(3) <= VNStageIntLLROutputS6xD(236)(2);
  CNStageIntLLRInputS7xD(221)(3) <= VNStageIntLLROutputS6xD(236)(3);
  CNStageIntLLRInputS7xD(271)(3) <= VNStageIntLLROutputS6xD(236)(4);
  CNStageIntLLRInputS7xD(310)(3) <= VNStageIntLLROutputS6xD(236)(5);
  CNStageIntLLRInputS7xD(10)(3) <= VNStageIntLLROutputS6xD(237)(0);
  CNStageIntLLRInputS7xD(110)(3) <= VNStageIntLLROutputS6xD(237)(1);
  CNStageIntLLRInputS7xD(125)(3) <= VNStageIntLLROutputS6xD(237)(2);
  CNStageIntLLRInputS7xD(228)(3) <= VNStageIntLLROutputS6xD(237)(3);
  CNStageIntLLRInputS7xD(322)(3) <= VNStageIntLLROutputS6xD(237)(4);
  CNStageIntLLRInputS7xD(334)(3) <= VNStageIntLLROutputS6xD(237)(5);
  CNStageIntLLRInputS7xD(9)(3) <= VNStageIntLLROutputS6xD(238)(0);
  CNStageIntLLRInputS7xD(103)(3) <= VNStageIntLLROutputS6xD(238)(1);
  CNStageIntLLRInputS7xD(113)(3) <= VNStageIntLLROutputS6xD(238)(2);
  CNStageIntLLRInputS7xD(179)(3) <= VNStageIntLLROutputS6xD(238)(3);
  CNStageIntLLRInputS7xD(236)(3) <= VNStageIntLLROutputS6xD(238)(4);
  CNStageIntLLRInputS7xD(294)(3) <= VNStageIntLLROutputS6xD(238)(5);
  CNStageIntLLRInputS7xD(383)(3) <= VNStageIntLLROutputS6xD(238)(6);
  CNStageIntLLRInputS7xD(8)(3) <= VNStageIntLLROutputS6xD(239)(0);
  CNStageIntLLRInputS7xD(98)(3) <= VNStageIntLLROutputS6xD(239)(1);
  CNStageIntLLRInputS7xD(158)(3) <= VNStageIntLLROutputS6xD(239)(2);
  CNStageIntLLRInputS7xD(223)(3) <= VNStageIntLLROutputS6xD(239)(3);
  CNStageIntLLRInputS7xD(264)(3) <= VNStageIntLLROutputS6xD(239)(4);
  CNStageIntLLRInputS7xD(284)(3) <= VNStageIntLLROutputS6xD(239)(5);
  CNStageIntLLRInputS7xD(360)(3) <= VNStageIntLLROutputS6xD(239)(6);
  CNStageIntLLRInputS7xD(7)(3) <= VNStageIntLLROutputS6xD(240)(0);
  CNStageIntLLRInputS7xD(81)(3) <= VNStageIntLLROutputS6xD(240)(1);
  CNStageIntLLRInputS7xD(116)(3) <= VNStageIntLLROutputS6xD(240)(2);
  CNStageIntLLRInputS7xD(210)(3) <= VNStageIntLLROutputS6xD(240)(3);
  CNStageIntLLRInputS7xD(277)(3) <= VNStageIntLLROutputS6xD(240)(4);
  CNStageIntLLRInputS7xD(324)(3) <= VNStageIntLLROutputS6xD(240)(5);
  CNStageIntLLRInputS7xD(343)(3) <= VNStageIntLLROutputS6xD(240)(6);
  CNStageIntLLRInputS7xD(6)(3) <= VNStageIntLLROutputS6xD(241)(0);
  CNStageIntLLRInputS7xD(88)(3) <= VNStageIntLLROutputS6xD(241)(1);
  CNStageIntLLRInputS7xD(175)(3) <= VNStageIntLLROutputS6xD(241)(2);
  CNStageIntLLRInputS7xD(250)(3) <= VNStageIntLLROutputS6xD(241)(3);
  CNStageIntLLRInputS7xD(285)(3) <= VNStageIntLLROutputS6xD(241)(4);
  CNStageIntLLRInputS7xD(355)(3) <= VNStageIntLLROutputS6xD(241)(5);
  CNStageIntLLRInputS7xD(5)(3) <= VNStageIntLLROutputS6xD(242)(0);
  CNStageIntLLRInputS7xD(108)(3) <= VNStageIntLLROutputS6xD(242)(1);
  CNStageIntLLRInputS7xD(146)(3) <= VNStageIntLLROutputS6xD(242)(2);
  CNStageIntLLRInputS7xD(203)(3) <= VNStageIntLLROutputS6xD(242)(3);
  CNStageIntLLRInputS7xD(231)(3) <= VNStageIntLLROutputS6xD(242)(4);
  CNStageIntLLRInputS7xD(303)(3) <= VNStageIntLLROutputS6xD(242)(5);
  CNStageIntLLRInputS7xD(367)(3) <= VNStageIntLLROutputS6xD(242)(6);
  CNStageIntLLRInputS7xD(4)(3) <= VNStageIntLLROutputS6xD(243)(0);
  CNStageIntLLRInputS7xD(106)(3) <= VNStageIntLLROutputS6xD(243)(1);
  CNStageIntLLRInputS7xD(141)(3) <= VNStageIntLLROutputS6xD(243)(2);
  CNStageIntLLRInputS7xD(200)(3) <= VNStageIntLLROutputS6xD(243)(3);
  CNStageIntLLRInputS7xD(252)(3) <= VNStageIntLLROutputS6xD(243)(4);
  CNStageIntLLRInputS7xD(312)(3) <= VNStageIntLLROutputS6xD(243)(5);
  CNStageIntLLRInputS7xD(337)(3) <= VNStageIntLLROutputS6xD(243)(6);
  CNStageIntLLRInputS7xD(147)(3) <= VNStageIntLLROutputS6xD(244)(0);
  CNStageIntLLRInputS7xD(266)(3) <= VNStageIntLLROutputS6xD(244)(1);
  CNStageIntLLRInputS7xD(3)(3) <= VNStageIntLLROutputS6xD(245)(0);
  CNStageIntLLRInputS7xD(66)(3) <= VNStageIntLLROutputS6xD(245)(1);
  CNStageIntLLRInputS7xD(136)(3) <= VNStageIntLLROutputS6xD(245)(2);
  CNStageIntLLRInputS7xD(207)(3) <= VNStageIntLLROutputS6xD(245)(3);
  CNStageIntLLRInputS7xD(262)(3) <= VNStageIntLLROutputS6xD(245)(4);
  CNStageIntLLRInputS7xD(313)(3) <= VNStageIntLLROutputS6xD(245)(5);
  CNStageIntLLRInputS7xD(370)(3) <= VNStageIntLLROutputS6xD(245)(6);
  CNStageIntLLRInputS7xD(2)(3) <= VNStageIntLLROutputS6xD(246)(0);
  CNStageIntLLRInputS7xD(69)(3) <= VNStageIntLLROutputS6xD(246)(1);
  CNStageIntLLRInputS7xD(161)(3) <= VNStageIntLLROutputS6xD(246)(2);
  CNStageIntLLRInputS7xD(185)(3) <= VNStageIntLLROutputS6xD(246)(3);
  CNStageIntLLRInputS7xD(226)(3) <= VNStageIntLLROutputS6xD(246)(4);
  CNStageIntLLRInputS7xD(302)(3) <= VNStageIntLLROutputS6xD(246)(5);
  CNStageIntLLRInputS7xD(1)(3) <= VNStageIntLLROutputS6xD(247)(0);
  CNStageIntLLRInputS7xD(109)(3) <= VNStageIntLLROutputS6xD(247)(1);
  CNStageIntLLRInputS7xD(168)(3) <= VNStageIntLLROutputS6xD(247)(2);
  CNStageIntLLRInputS7xD(194)(3) <= VNStageIntLLROutputS6xD(247)(3);
  CNStageIntLLRInputS7xD(247)(3) <= VNStageIntLLROutputS6xD(247)(4);
  CNStageIntLLRInputS7xD(327)(3) <= VNStageIntLLROutputS6xD(247)(5);
  CNStageIntLLRInputS7xD(349)(3) <= VNStageIntLLROutputS6xD(247)(6);
  CNStageIntLLRInputS7xD(0)(3) <= VNStageIntLLROutputS6xD(248)(0);
  CNStageIntLLRInputS7xD(87)(3) <= VNStageIntLLROutputS6xD(248)(1);
  CNStageIntLLRInputS7xD(151)(3) <= VNStageIntLLROutputS6xD(248)(2);
  CNStageIntLLRInputS7xD(189)(3) <= VNStageIntLLROutputS6xD(248)(3);
  CNStageIntLLRInputS7xD(248)(3) <= VNStageIntLLROutputS6xD(248)(4);
  CNStageIntLLRInputS7xD(280)(3) <= VNStageIntLLROutputS6xD(248)(5);
  CNStageIntLLRInputS7xD(357)(3) <= VNStageIntLLROutputS6xD(248)(6);
  CNStageIntLLRInputS7xD(152)(3) <= VNStageIntLLROutputS6xD(249)(0);
  CNStageIntLLRInputS7xD(192)(3) <= VNStageIntLLROutputS6xD(249)(1);
  CNStageIntLLRInputS7xD(225)(3) <= VNStageIntLLROutputS6xD(249)(2);
  CNStageIntLLRInputS7xD(317)(3) <= VNStageIntLLROutputS6xD(249)(3);
  CNStageIntLLRInputS7xD(353)(3) <= VNStageIntLLROutputS6xD(249)(4);
  CNStageIntLLRInputS7xD(79)(3) <= VNStageIntLLROutputS6xD(250)(0);
  CNStageIntLLRInputS7xD(120)(3) <= VNStageIntLLROutputS6xD(250)(1);
  CNStageIntLLRInputS7xD(184)(3) <= VNStageIntLLROutputS6xD(250)(2);
  CNStageIntLLRInputS7xD(319)(3) <= VNStageIntLLROutputS6xD(250)(3);
  CNStageIntLLRInputS7xD(358)(3) <= VNStageIntLLROutputS6xD(250)(4);
  CNStageIntLLRInputS7xD(62)(3) <= VNStageIntLLROutputS6xD(251)(0);
  CNStageIntLLRInputS7xD(159)(3) <= VNStageIntLLROutputS6xD(251)(1);
  CNStageIntLLRInputS7xD(215)(3) <= VNStageIntLLROutputS6xD(251)(2);
  CNStageIntLLRInputS7xD(289)(3) <= VNStageIntLLROutputS6xD(251)(3);
  CNStageIntLLRInputS7xD(348)(3) <= VNStageIntLLROutputS6xD(251)(4);
  CNStageIntLLRInputS7xD(89)(3) <= VNStageIntLLROutputS6xD(252)(0);
  CNStageIntLLRInputS7xD(112)(3) <= VNStageIntLLROutputS6xD(252)(1);
  CNStageIntLLRInputS7xD(199)(3) <= VNStageIntLLROutputS6xD(252)(2);
  CNStageIntLLRInputS7xD(239)(3) <= VNStageIntLLROutputS6xD(252)(3);
  CNStageIntLLRInputS7xD(325)(3) <= VNStageIntLLROutputS6xD(252)(4);
  CNStageIntLLRInputS7xD(373)(3) <= VNStageIntLLROutputS6xD(252)(5);
  CNStageIntLLRInputS7xD(80)(3) <= VNStageIntLLROutputS6xD(253)(0);
  CNStageIntLLRInputS7xD(121)(3) <= VNStageIntLLROutputS6xD(253)(1);
  CNStageIntLLRInputS7xD(211)(3) <= VNStageIntLLROutputS6xD(253)(2);
  CNStageIntLLRInputS7xD(279)(3) <= VNStageIntLLROutputS6xD(253)(3);
  CNStageIntLLRInputS7xD(283)(3) <= VNStageIntLLROutputS6xD(253)(4);
  CNStageIntLLRInputS7xD(380)(3) <= VNStageIntLLROutputS6xD(253)(5);
  CNStageIntLLRInputS7xD(67)(3) <= VNStageIntLLROutputS6xD(254)(0);
  CNStageIntLLRInputS7xD(222)(3) <= VNStageIntLLROutputS6xD(254)(1);
  CNStageIntLLRInputS7xD(238)(3) <= VNStageIntLLROutputS6xD(254)(2);
  CNStageIntLLRInputS7xD(290)(3) <= VNStageIntLLROutputS6xD(254)(3);
  CNStageIntLLRInputS7xD(362)(3) <= VNStageIntLLROutputS6xD(254)(4);
  CNStageIntLLRInputS7xD(52)(3) <= VNStageIntLLROutputS6xD(255)(0);
  CNStageIntLLRInputS7xD(86)(3) <= VNStageIntLLROutputS6xD(255)(1);
  CNStageIntLLRInputS7xD(167)(3) <= VNStageIntLLROutputS6xD(255)(2);
  CNStageIntLLRInputS7xD(195)(3) <= VNStageIntLLROutputS6xD(255)(3);
  CNStageIntLLRInputS7xD(233)(3) <= VNStageIntLLROutputS6xD(255)(4);
  CNStageIntLLRInputS7xD(318)(3) <= VNStageIntLLROutputS6xD(255)(5);
  CNStageIntLLRInputS7xD(364)(3) <= VNStageIntLLROutputS6xD(255)(6);
  CNStageIntLLRInputS7xD(53)(4) <= VNStageIntLLROutputS6xD(256)(0);
  CNStageIntLLRInputS7xD(106)(4) <= VNStageIntLLROutputS6xD(256)(1);
  CNStageIntLLRInputS7xD(127)(4) <= VNStageIntLLROutputS6xD(256)(2);
  CNStageIntLLRInputS7xD(242)(4) <= VNStageIntLLROutputS6xD(256)(3);
  CNStageIntLLRInputS7xD(296)(4) <= VNStageIntLLROutputS6xD(256)(4);
  CNStageIntLLRInputS7xD(339)(4) <= VNStageIntLLROutputS6xD(256)(5);
  CNStageIntLLRInputS7xD(51)(4) <= VNStageIntLLROutputS6xD(257)(0);
  CNStageIntLLRInputS7xD(85)(4) <= VNStageIntLLROutputS6xD(257)(1);
  CNStageIntLLRInputS7xD(166)(4) <= VNStageIntLLROutputS6xD(257)(2);
  CNStageIntLLRInputS7xD(194)(4) <= VNStageIntLLROutputS6xD(257)(3);
  CNStageIntLLRInputS7xD(232)(4) <= VNStageIntLLROutputS6xD(257)(4);
  CNStageIntLLRInputS7xD(317)(4) <= VNStageIntLLROutputS6xD(257)(5);
  CNStageIntLLRInputS7xD(363)(4) <= VNStageIntLLROutputS6xD(257)(6);
  CNStageIntLLRInputS7xD(50)(4) <= VNStageIntLLROutputS6xD(258)(0);
  CNStageIntLLRInputS7xD(57)(4) <= VNStageIntLLROutputS6xD(258)(1);
  CNStageIntLLRInputS7xD(331)(4) <= VNStageIntLLROutputS6xD(258)(2);
  CNStageIntLLRInputS7xD(54)(4) <= VNStageIntLLROutputS6xD(259)(0);
  CNStageIntLLRInputS7xD(114)(4) <= VNStageIntLLROutputS6xD(259)(1);
  CNStageIntLLRInputS7xD(274)(4) <= VNStageIntLLROutputS6xD(259)(2);
  CNStageIntLLRInputS7xD(303)(4) <= VNStageIntLLROutputS6xD(259)(3);
  CNStageIntLLRInputS7xD(370)(4) <= VNStageIntLLROutputS6xD(259)(4);
  CNStageIntLLRInputS7xD(49)(4) <= VNStageIntLLROutputS6xD(260)(0);
  CNStageIntLLRInputS7xD(71)(4) <= VNStageIntLLROutputS6xD(260)(1);
  CNStageIntLLRInputS7xD(138)(4) <= VNStageIntLLROutputS6xD(260)(2);
  CNStageIntLLRInputS7xD(186)(4) <= VNStageIntLLROutputS6xD(260)(3);
  CNStageIntLLRInputS7xD(243)(4) <= VNStageIntLLROutputS6xD(260)(4);
  CNStageIntLLRInputS7xD(383)(4) <= VNStageIntLLROutputS6xD(260)(5);
  CNStageIntLLRInputS7xD(48)(4) <= VNStageIntLLROutputS6xD(261)(0);
  CNStageIntLLRInputS7xD(63)(4) <= VNStageIntLLROutputS6xD(261)(1);
  CNStageIntLLRInputS7xD(152)(4) <= VNStageIntLLROutputS6xD(261)(2);
  CNStageIntLLRInputS7xD(204)(4) <= VNStageIntLLROutputS6xD(261)(3);
  CNStageIntLLRInputS7xD(305)(4) <= VNStageIntLLROutputS6xD(261)(4);
  CNStageIntLLRInputS7xD(333)(4) <= VNStageIntLLROutputS6xD(261)(5);
  CNStageIntLLRInputS7xD(47)(4) <= VNStageIntLLROutputS6xD(262)(0);
  CNStageIntLLRInputS7xD(95)(4) <= VNStageIntLLROutputS6xD(262)(1);
  CNStageIntLLRInputS7xD(149)(4) <= VNStageIntLLROutputS6xD(262)(2);
  CNStageIntLLRInputS7xD(212)(4) <= VNStageIntLLROutputS6xD(262)(3);
  CNStageIntLLRInputS7xD(319)(4) <= VNStageIntLLROutputS6xD(262)(4);
  CNStageIntLLRInputS7xD(362)(4) <= VNStageIntLLROutputS6xD(262)(5);
  CNStageIntLLRInputS7xD(46)(4) <= VNStageIntLLROutputS6xD(263)(0);
  CNStageIntLLRInputS7xD(104)(4) <= VNStageIntLLROutputS6xD(263)(1);
  CNStageIntLLRInputS7xD(169)(4) <= VNStageIntLLROutputS6xD(263)(2);
  CNStageIntLLRInputS7xD(207)(4) <= VNStageIntLLROutputS6xD(263)(3);
  CNStageIntLLRInputS7xD(253)(4) <= VNStageIntLLROutputS6xD(263)(4);
  CNStageIntLLRInputS7xD(315)(4) <= VNStageIntLLROutputS6xD(263)(5);
  CNStageIntLLRInputS7xD(378)(4) <= VNStageIntLLROutputS6xD(263)(6);
  CNStageIntLLRInputS7xD(45)(4) <= VNStageIntLLROutputS6xD(264)(0);
  CNStageIntLLRInputS7xD(98)(4) <= VNStageIntLLROutputS6xD(264)(1);
  CNStageIntLLRInputS7xD(132)(4) <= VNStageIntLLROutputS6xD(264)(2);
  CNStageIntLLRInputS7xD(213)(4) <= VNStageIntLLROutputS6xD(264)(3);
  CNStageIntLLRInputS7xD(256)(4) <= VNStageIntLLROutputS6xD(264)(4);
  CNStageIntLLRInputS7xD(281)(4) <= VNStageIntLLROutputS6xD(264)(5);
  CNStageIntLLRInputS7xD(349)(4) <= VNStageIntLLROutputS6xD(264)(6);
  CNStageIntLLRInputS7xD(44)(4) <= VNStageIntLLROutputS6xD(265)(0);
  CNStageIntLLRInputS7xD(133)(4) <= VNStageIntLLROutputS6xD(265)(1);
  CNStageIntLLRInputS7xD(203)(4) <= VNStageIntLLROutputS6xD(265)(2);
  CNStageIntLLRInputS7xD(244)(4) <= VNStageIntLLROutputS6xD(265)(3);
  CNStageIntLLRInputS7xD(43)(4) <= VNStageIntLLROutputS6xD(266)(0);
  CNStageIntLLRInputS7xD(168)(4) <= VNStageIntLLROutputS6xD(266)(1);
  CNStageIntLLRInputS7xD(173)(4) <= VNStageIntLLROutputS6xD(266)(2);
  CNStageIntLLRInputS7xD(273)(4) <= VNStageIntLLROutputS6xD(266)(3);
  CNStageIntLLRInputS7xD(300)(4) <= VNStageIntLLROutputS6xD(266)(4);
  CNStageIntLLRInputS7xD(42)(4) <= VNStageIntLLROutputS6xD(267)(0);
  CNStageIntLLRInputS7xD(72)(4) <= VNStageIntLLROutputS6xD(267)(1);
  CNStageIntLLRInputS7xD(159)(4) <= VNStageIntLLROutputS6xD(267)(2);
  CNStageIntLLRInputS7xD(180)(4) <= VNStageIntLLROutputS6xD(267)(3);
  CNStageIntLLRInputS7xD(241)(4) <= VNStageIntLLROutputS6xD(267)(4);
  CNStageIntLLRInputS7xD(280)(4) <= VNStageIntLLROutputS6xD(267)(5);
  CNStageIntLLRInputS7xD(364)(4) <= VNStageIntLLROutputS6xD(267)(6);
  CNStageIntLLRInputS7xD(41)(4) <= VNStageIntLLROutputS6xD(268)(0);
  CNStageIntLLRInputS7xD(109)(4) <= VNStageIntLLROutputS6xD(268)(1);
  CNStageIntLLRInputS7xD(118)(4) <= VNStageIntLLROutputS6xD(268)(2);
  CNStageIntLLRInputS7xD(216)(4) <= VNStageIntLLROutputS6xD(268)(3);
  CNStageIntLLRInputS7xD(266)(4) <= VNStageIntLLROutputS6xD(268)(4);
  CNStageIntLLRInputS7xD(325)(4) <= VNStageIntLLROutputS6xD(268)(5);
  CNStageIntLLRInputS7xD(360)(4) <= VNStageIntLLROutputS6xD(268)(6);
  CNStageIntLLRInputS7xD(67)(4) <= VNStageIntLLROutputS6xD(269)(0);
  CNStageIntLLRInputS7xD(122)(4) <= VNStageIntLLROutputS6xD(269)(1);
  CNStageIntLLRInputS7xD(218)(4) <= VNStageIntLLROutputS6xD(269)(2);
  CNStageIntLLRInputS7xD(250)(4) <= VNStageIntLLROutputS6xD(269)(3);
  CNStageIntLLRInputS7xD(287)(4) <= VNStageIntLLROutputS6xD(269)(4);
  CNStageIntLLRInputS7xD(381)(4) <= VNStageIntLLROutputS6xD(269)(5);
  CNStageIntLLRInputS7xD(40)(4) <= VNStageIntLLROutputS6xD(270)(0);
  CNStageIntLLRInputS7xD(79)(4) <= VNStageIntLLROutputS6xD(270)(1);
  CNStageIntLLRInputS7xD(170)(4) <= VNStageIntLLROutputS6xD(270)(2);
  CNStageIntLLRInputS7xD(190)(4) <= VNStageIntLLROutputS6xD(270)(3);
  CNStageIntLLRInputS7xD(275)(4) <= VNStageIntLLROutputS6xD(270)(4);
  CNStageIntLLRInputS7xD(292)(4) <= VNStageIntLLROutputS6xD(270)(5);
  CNStageIntLLRInputS7xD(344)(4) <= VNStageIntLLROutputS6xD(270)(6);
  CNStageIntLLRInputS7xD(39)(4) <= VNStageIntLLROutputS6xD(271)(0);
  CNStageIntLLRInputS7xD(105)(4) <= VNStageIntLLROutputS6xD(271)(1);
  CNStageIntLLRInputS7xD(171)(4) <= VNStageIntLLROutputS6xD(271)(2);
  CNStageIntLLRInputS7xD(268)(4) <= VNStageIntLLROutputS6xD(271)(3);
  CNStageIntLLRInputS7xD(332)(4) <= VNStageIntLLROutputS6xD(271)(4);
  CNStageIntLLRInputS7xD(345)(4) <= VNStageIntLLROutputS6xD(271)(5);
  CNStageIntLLRInputS7xD(38)(4) <= VNStageIntLLROutputS6xD(272)(0);
  CNStageIntLLRInputS7xD(94)(4) <= VNStageIntLLROutputS6xD(272)(1);
  CNStageIntLLRInputS7xD(116)(4) <= VNStageIntLLROutputS6xD(272)(2);
  CNStageIntLLRInputS7xD(184)(4) <= VNStageIntLLROutputS6xD(272)(3);
  CNStageIntLLRInputS7xD(254)(4) <= VNStageIntLLROutputS6xD(272)(4);
  CNStageIntLLRInputS7xD(291)(4) <= VNStageIntLLROutputS6xD(272)(5);
  CNStageIntLLRInputS7xD(380)(4) <= VNStageIntLLROutputS6xD(272)(6);
  CNStageIntLLRInputS7xD(37)(4) <= VNStageIntLLROutputS6xD(273)(0);
  CNStageIntLLRInputS7xD(81)(4) <= VNStageIntLLROutputS6xD(273)(1);
  CNStageIntLLRInputS7xD(156)(4) <= VNStageIntLLROutputS6xD(273)(2);
  CNStageIntLLRInputS7xD(272)(4) <= VNStageIntLLROutputS6xD(273)(3);
  CNStageIntLLRInputS7xD(285)(4) <= VNStageIntLLROutputS6xD(273)(4);
  CNStageIntLLRInputS7xD(371)(4) <= VNStageIntLLROutputS6xD(273)(5);
  CNStageIntLLRInputS7xD(36)(4) <= VNStageIntLLROutputS6xD(274)(0);
  CNStageIntLLRInputS7xD(164)(4) <= VNStageIntLLROutputS6xD(274)(1);
  CNStageIntLLRInputS7xD(217)(4) <= VNStageIntLLROutputS6xD(274)(2);
  CNStageIntLLRInputS7xD(248)(4) <= VNStageIntLLROutputS6xD(274)(3);
  CNStageIntLLRInputS7xD(35)(4) <= VNStageIntLLROutputS6xD(275)(0);
  CNStageIntLLRInputS7xD(59)(4) <= VNStageIntLLROutputS6xD(275)(1);
  CNStageIntLLRInputS7xD(128)(4) <= VNStageIntLLROutputS6xD(275)(2);
  CNStageIntLLRInputS7xD(179)(4) <= VNStageIntLLROutputS6xD(275)(3);
  CNStageIntLLRInputS7xD(329)(4) <= VNStageIntLLROutputS6xD(275)(4);
  CNStageIntLLRInputS7xD(34)(4) <= VNStageIntLLROutputS6xD(276)(0);
  CNStageIntLLRInputS7xD(69)(4) <= VNStageIntLLROutputS6xD(276)(1);
  CNStageIntLLRInputS7xD(126)(4) <= VNStageIntLLROutputS6xD(276)(2);
  CNStageIntLLRInputS7xD(205)(4) <= VNStageIntLLROutputS6xD(276)(3);
  CNStageIntLLRInputS7xD(259)(4) <= VNStageIntLLROutputS6xD(276)(4);
  CNStageIntLLRInputS7xD(297)(4) <= VNStageIntLLROutputS6xD(276)(5);
  CNStageIntLLRInputS7xD(33)(4) <= VNStageIntLLROutputS6xD(277)(0);
  CNStageIntLLRInputS7xD(64)(4) <= VNStageIntLLROutputS6xD(277)(1);
  CNStageIntLLRInputS7xD(162)(4) <= VNStageIntLLROutputS6xD(277)(2);
  CNStageIntLLRInputS7xD(185)(4) <= VNStageIntLLROutputS6xD(277)(3);
  CNStageIntLLRInputS7xD(252)(4) <= VNStageIntLLROutputS6xD(277)(4);
  CNStageIntLLRInputS7xD(295)(4) <= VNStageIntLLROutputS6xD(277)(5);
  CNStageIntLLRInputS7xD(334)(4) <= VNStageIntLLROutputS6xD(277)(6);
  CNStageIntLLRInputS7xD(32)(4) <= VNStageIntLLROutputS6xD(278)(0);
  CNStageIntLLRInputS7xD(70)(4) <= VNStageIntLLROutputS6xD(278)(1);
  CNStageIntLLRInputS7xD(141)(4) <= VNStageIntLLROutputS6xD(278)(2);
  CNStageIntLLRInputS7xD(229)(4) <= VNStageIntLLROutputS6xD(278)(3);
  CNStageIntLLRInputS7xD(328)(4) <= VNStageIntLLROutputS6xD(278)(4);
  CNStageIntLLRInputS7xD(31)(4) <= VNStageIntLLROutputS6xD(279)(0);
  CNStageIntLLRInputS7xD(58)(4) <= VNStageIntLLROutputS6xD(279)(1);
  CNStageIntLLRInputS7xD(144)(4) <= VNStageIntLLROutputS6xD(279)(2);
  CNStageIntLLRInputS7xD(219)(4) <= VNStageIntLLROutputS6xD(279)(3);
  CNStageIntLLRInputS7xD(239)(4) <= VNStageIntLLROutputS6xD(279)(4);
  CNStageIntLLRInputS7xD(368)(4) <= VNStageIntLLROutputS6xD(279)(5);
  CNStageIntLLRInputS7xD(30)(4) <= VNStageIntLLROutputS6xD(280)(0);
  CNStageIntLLRInputS7xD(84)(4) <= VNStageIntLLROutputS6xD(280)(1);
  CNStageIntLLRInputS7xD(129)(4) <= VNStageIntLLROutputS6xD(280)(2);
  CNStageIntLLRInputS7xD(215)(4) <= VNStageIntLLROutputS6xD(280)(3);
  CNStageIntLLRInputS7xD(233)(4) <= VNStageIntLLROutputS6xD(280)(4);
  CNStageIntLLRInputS7xD(310)(4) <= VNStageIntLLROutputS6xD(280)(5);
  CNStageIntLLRInputS7xD(376)(4) <= VNStageIntLLROutputS6xD(280)(6);
  CNStageIntLLRInputS7xD(29)(4) <= VNStageIntLLROutputS6xD(281)(0);
  CNStageIntLLRInputS7xD(90)(4) <= VNStageIntLLROutputS6xD(281)(1);
  CNStageIntLLRInputS7xD(163)(4) <= VNStageIntLLROutputS6xD(281)(2);
  CNStageIntLLRInputS7xD(182)(4) <= VNStageIntLLROutputS6xD(281)(3);
  CNStageIntLLRInputS7xD(236)(4) <= VNStageIntLLROutputS6xD(281)(4);
  CNStageIntLLRInputS7xD(298)(4) <= VNStageIntLLROutputS6xD(281)(5);
  CNStageIntLLRInputS7xD(340)(4) <= VNStageIntLLROutputS6xD(281)(6);
  CNStageIntLLRInputS7xD(28)(4) <= VNStageIntLLROutputS6xD(282)(0);
  CNStageIntLLRInputS7xD(74)(4) <= VNStageIntLLROutputS6xD(282)(1);
  CNStageIntLLRInputS7xD(125)(4) <= VNStageIntLLROutputS6xD(282)(2);
  CNStageIntLLRInputS7xD(200)(4) <= VNStageIntLLROutputS6xD(282)(3);
  CNStageIntLLRInputS7xD(226)(4) <= VNStageIntLLROutputS6xD(282)(4);
  CNStageIntLLRInputS7xD(338)(4) <= VNStageIntLLROutputS6xD(282)(5);
  CNStageIntLLRInputS7xD(27)(4) <= VNStageIntLLROutputS6xD(283)(0);
  CNStageIntLLRInputS7xD(76)(4) <= VNStageIntLLROutputS6xD(283)(1);
  CNStageIntLLRInputS7xD(153)(4) <= VNStageIntLLROutputS6xD(283)(2);
  CNStageIntLLRInputS7xD(201)(4) <= VNStageIntLLROutputS6xD(283)(3);
  CNStageIntLLRInputS7xD(260)(4) <= VNStageIntLLROutputS6xD(283)(4);
  CNStageIntLLRInputS7xD(294)(4) <= VNStageIntLLROutputS6xD(283)(5);
  CNStageIntLLRInputS7xD(374)(4) <= VNStageIntLLROutputS6xD(283)(6);
  CNStageIntLLRInputS7xD(26)(4) <= VNStageIntLLROutputS6xD(284)(0);
  CNStageIntLLRInputS7xD(100)(4) <= VNStageIntLLROutputS6xD(284)(1);
  CNStageIntLLRInputS7xD(137)(4) <= VNStageIntLLROutputS6xD(284)(2);
  CNStageIntLLRInputS7xD(181)(4) <= VNStageIntLLROutputS6xD(284)(3);
  CNStageIntLLRInputS7xD(245)(4) <= VNStageIntLLROutputS6xD(284)(4);
  CNStageIntLLRInputS7xD(320)(4) <= VNStageIntLLROutputS6xD(284)(5);
  CNStageIntLLRInputS7xD(353)(4) <= VNStageIntLLROutputS6xD(284)(6);
  CNStageIntLLRInputS7xD(25)(4) <= VNStageIntLLROutputS6xD(285)(0);
  CNStageIntLLRInputS7xD(82)(4) <= VNStageIntLLROutputS6xD(285)(1);
  CNStageIntLLRInputS7xD(165)(4) <= VNStageIntLLROutputS6xD(285)(2);
  CNStageIntLLRInputS7xD(172)(4) <= VNStageIntLLROutputS6xD(285)(3);
  CNStageIntLLRInputS7xD(255)(4) <= VNStageIntLLROutputS6xD(285)(4);
  CNStageIntLLRInputS7xD(304)(4) <= VNStageIntLLROutputS6xD(285)(5);
  CNStageIntLLRInputS7xD(355)(4) <= VNStageIntLLROutputS6xD(285)(6);
  CNStageIntLLRInputS7xD(24)(4) <= VNStageIntLLROutputS6xD(286)(0);
  CNStageIntLLRInputS7xD(93)(4) <= VNStageIntLLROutputS6xD(286)(1);
  CNStageIntLLRInputS7xD(155)(4) <= VNStageIntLLROutputS6xD(286)(2);
  CNStageIntLLRInputS7xD(189)(4) <= VNStageIntLLROutputS6xD(286)(3);
  CNStageIntLLRInputS7xD(267)(4) <= VNStageIntLLROutputS6xD(286)(4);
  CNStageIntLLRInputS7xD(330)(4) <= VNStageIntLLROutputS6xD(286)(5);
  CNStageIntLLRInputS7xD(341)(4) <= VNStageIntLLROutputS6xD(286)(6);
  CNStageIntLLRInputS7xD(23)(4) <= VNStageIntLLROutputS6xD(287)(0);
  CNStageIntLLRInputS7xD(101)(4) <= VNStageIntLLROutputS6xD(287)(1);
  CNStageIntLLRInputS7xD(142)(4) <= VNStageIntLLROutputS6xD(287)(2);
  CNStageIntLLRInputS7xD(193)(4) <= VNStageIntLLROutputS6xD(287)(3);
  CNStageIntLLRInputS7xD(240)(4) <= VNStageIntLLROutputS6xD(287)(4);
  CNStageIntLLRInputS7xD(322)(4) <= VNStageIntLLROutputS6xD(287)(5);
  CNStageIntLLRInputS7xD(375)(4) <= VNStageIntLLROutputS6xD(287)(6);
  CNStageIntLLRInputS7xD(22)(4) <= VNStageIntLLROutputS6xD(288)(0);
  CNStageIntLLRInputS7xD(75)(4) <= VNStageIntLLROutputS6xD(288)(1);
  CNStageIntLLRInputS7xD(161)(4) <= VNStageIntLLROutputS6xD(288)(2);
  CNStageIntLLRInputS7xD(224)(4) <= VNStageIntLLROutputS6xD(288)(3);
  CNStageIntLLRInputS7xD(228)(4) <= VNStageIntLLROutputS6xD(288)(4);
  CNStageIntLLRInputS7xD(308)(4) <= VNStageIntLLROutputS6xD(288)(5);
  CNStageIntLLRInputS7xD(337)(4) <= VNStageIntLLROutputS6xD(288)(6);
  CNStageIntLLRInputS7xD(21)(4) <= VNStageIntLLROutputS6xD(289)(0);
  CNStageIntLLRInputS7xD(89)(4) <= VNStageIntLLROutputS6xD(289)(1);
  CNStageIntLLRInputS7xD(134)(4) <= VNStageIntLLROutputS6xD(289)(2);
  CNStageIntLLRInputS7xD(192)(4) <= VNStageIntLLROutputS6xD(289)(3);
  CNStageIntLLRInputS7xD(269)(4) <= VNStageIntLLROutputS6xD(289)(4);
  CNStageIntLLRInputS7xD(327)(4) <= VNStageIntLLROutputS6xD(289)(5);
  CNStageIntLLRInputS7xD(365)(4) <= VNStageIntLLROutputS6xD(289)(6);
  CNStageIntLLRInputS7xD(20)(4) <= VNStageIntLLROutputS6xD(290)(0);
  CNStageIntLLRInputS7xD(60)(4) <= VNStageIntLLROutputS6xD(290)(1);
  CNStageIntLLRInputS7xD(131)(4) <= VNStageIntLLROutputS6xD(290)(2);
  CNStageIntLLRInputS7xD(187)(4) <= VNStageIntLLROutputS6xD(290)(3);
  CNStageIntLLRInputS7xD(231)(4) <= VNStageIntLLROutputS6xD(290)(4);
  CNStageIntLLRInputS7xD(350)(4) <= VNStageIntLLROutputS6xD(290)(5);
  CNStageIntLLRInputS7xD(19)(4) <= VNStageIntLLROutputS6xD(291)(0);
  CNStageIntLLRInputS7xD(96)(4) <= VNStageIntLLROutputS6xD(291)(1);
  CNStageIntLLRInputS7xD(147)(4) <= VNStageIntLLROutputS6xD(291)(2);
  CNStageIntLLRInputS7xD(223)(4) <= VNStageIntLLROutputS6xD(291)(3);
  CNStageIntLLRInputS7xD(249)(4) <= VNStageIntLLROutputS6xD(291)(4);
  CNStageIntLLRInputS7xD(377)(4) <= VNStageIntLLROutputS6xD(291)(5);
  CNStageIntLLRInputS7xD(18)(4) <= VNStageIntLLROutputS6xD(292)(0);
  CNStageIntLLRInputS7xD(62)(4) <= VNStageIntLLROutputS6xD(292)(1);
  CNStageIntLLRInputS7xD(139)(4) <= VNStageIntLLROutputS6xD(292)(2);
  CNStageIntLLRInputS7xD(177)(4) <= VNStageIntLLROutputS6xD(292)(3);
  CNStageIntLLRInputS7xD(257)(4) <= VNStageIntLLROutputS6xD(292)(4);
  CNStageIntLLRInputS7xD(313)(4) <= VNStageIntLLROutputS6xD(292)(5);
  CNStageIntLLRInputS7xD(367)(4) <= VNStageIntLLROutputS6xD(292)(6);
  CNStageIntLLRInputS7xD(17)(4) <= VNStageIntLLROutputS6xD(293)(0);
  CNStageIntLLRInputS7xD(77)(4) <= VNStageIntLLROutputS6xD(293)(1);
  CNStageIntLLRInputS7xD(113)(4) <= VNStageIntLLROutputS6xD(293)(2);
  CNStageIntLLRInputS7xD(197)(4) <= VNStageIntLLROutputS6xD(293)(3);
  CNStageIntLLRInputS7xD(306)(4) <= VNStageIntLLROutputS6xD(293)(4);
  CNStageIntLLRInputS7xD(354)(4) <= VNStageIntLLROutputS6xD(293)(5);
  CNStageIntLLRInputS7xD(16)(4) <= VNStageIntLLROutputS6xD(294)(0);
  CNStageIntLLRInputS7xD(73)(4) <= VNStageIntLLROutputS6xD(294)(1);
  CNStageIntLLRInputS7xD(123)(4) <= VNStageIntLLROutputS6xD(294)(2);
  CNStageIntLLRInputS7xD(196)(4) <= VNStageIntLLROutputS6xD(294)(3);
  CNStageIntLLRInputS7xD(258)(4) <= VNStageIntLLROutputS6xD(294)(4);
  CNStageIntLLRInputS7xD(284)(4) <= VNStageIntLLROutputS6xD(294)(5);
  CNStageIntLLRInputS7xD(373)(4) <= VNStageIntLLROutputS6xD(294)(6);
  CNStageIntLLRInputS7xD(15)(4) <= VNStageIntLLROutputS6xD(295)(0);
  CNStageIntLLRInputS7xD(92)(4) <= VNStageIntLLROutputS6xD(295)(1);
  CNStageIntLLRInputS7xD(117)(4) <= VNStageIntLLROutputS6xD(295)(2);
  CNStageIntLLRInputS7xD(175)(4) <= VNStageIntLLROutputS6xD(295)(3);
  CNStageIntLLRInputS7xD(346)(4) <= VNStageIntLLROutputS6xD(295)(4);
  CNStageIntLLRInputS7xD(14)(4) <= VNStageIntLLROutputS6xD(296)(0);
  CNStageIntLLRInputS7xD(55)(4) <= VNStageIntLLROutputS6xD(296)(1);
  CNStageIntLLRInputS7xD(121)(4) <= VNStageIntLLROutputS6xD(296)(2);
  CNStageIntLLRInputS7xD(208)(4) <= VNStageIntLLROutputS6xD(296)(3);
  CNStageIntLLRInputS7xD(286)(4) <= VNStageIntLLROutputS6xD(296)(4);
  CNStageIntLLRInputS7xD(343)(4) <= VNStageIntLLROutputS6xD(296)(5);
  CNStageIntLLRInputS7xD(13)(4) <= VNStageIntLLROutputS6xD(297)(0);
  CNStageIntLLRInputS7xD(56)(4) <= VNStageIntLLROutputS6xD(297)(1);
  CNStageIntLLRInputS7xD(111)(4) <= VNStageIntLLROutputS6xD(297)(2);
  CNStageIntLLRInputS7xD(211)(4) <= VNStageIntLLROutputS6xD(297)(3);
  CNStageIntLLRInputS7xD(277)(4) <= VNStageIntLLROutputS6xD(297)(4);
  CNStageIntLLRInputS7xD(290)(4) <= VNStageIntLLROutputS6xD(297)(5);
  CNStageIntLLRInputS7xD(358)(4) <= VNStageIntLLROutputS6xD(297)(6);
  CNStageIntLLRInputS7xD(12)(4) <= VNStageIntLLROutputS6xD(298)(0);
  CNStageIntLLRInputS7xD(91)(4) <= VNStageIntLLROutputS6xD(298)(1);
  CNStageIntLLRInputS7xD(148)(4) <= VNStageIntLLROutputS6xD(298)(2);
  CNStageIntLLRInputS7xD(198)(4) <= VNStageIntLLROutputS6xD(298)(3);
  CNStageIntLLRInputS7xD(262)(4) <= VNStageIntLLROutputS6xD(298)(4);
  CNStageIntLLRInputS7xD(282)(4) <= VNStageIntLLROutputS6xD(298)(5);
  CNStageIntLLRInputS7xD(351)(4) <= VNStageIntLLROutputS6xD(298)(6);
  CNStageIntLLRInputS7xD(83)(4) <= VNStageIntLLROutputS6xD(299)(0);
  CNStageIntLLRInputS7xD(130)(4) <= VNStageIntLLROutputS6xD(299)(1);
  CNStageIntLLRInputS7xD(176)(4) <= VNStageIntLLROutputS6xD(299)(2);
  CNStageIntLLRInputS7xD(264)(4) <= VNStageIntLLROutputS6xD(299)(3);
  CNStageIntLLRInputS7xD(314)(4) <= VNStageIntLLROutputS6xD(299)(4);
  CNStageIntLLRInputS7xD(11)(4) <= VNStageIntLLROutputS6xD(300)(0);
  CNStageIntLLRInputS7xD(99)(4) <= VNStageIntLLROutputS6xD(300)(1);
  CNStageIntLLRInputS7xD(143)(4) <= VNStageIntLLROutputS6xD(300)(2);
  CNStageIntLLRInputS7xD(195)(4) <= VNStageIntLLROutputS6xD(300)(3);
  CNStageIntLLRInputS7xD(299)(4) <= VNStageIntLLROutputS6xD(300)(4);
  CNStageIntLLRInputS7xD(335)(4) <= VNStageIntLLROutputS6xD(300)(5);
  CNStageIntLLRInputS7xD(10)(4) <= VNStageIntLLROutputS6xD(301)(0);
  CNStageIntLLRInputS7xD(103)(4) <= VNStageIntLLROutputS6xD(301)(1);
  CNStageIntLLRInputS7xD(154)(4) <= VNStageIntLLROutputS6xD(301)(2);
  CNStageIntLLRInputS7xD(220)(4) <= VNStageIntLLROutputS6xD(301)(3);
  CNStageIntLLRInputS7xD(270)(4) <= VNStageIntLLROutputS6xD(301)(4);
  CNStageIntLLRInputS7xD(309)(4) <= VNStageIntLLROutputS6xD(301)(5);
  CNStageIntLLRInputS7xD(9)(4) <= VNStageIntLLROutputS6xD(302)(0);
  CNStageIntLLRInputS7xD(110)(4) <= VNStageIntLLROutputS6xD(302)(1);
  CNStageIntLLRInputS7xD(124)(4) <= VNStageIntLLROutputS6xD(302)(2);
  CNStageIntLLRInputS7xD(206)(4) <= VNStageIntLLROutputS6xD(302)(3);
  CNStageIntLLRInputS7xD(227)(4) <= VNStageIntLLROutputS6xD(302)(4);
  CNStageIntLLRInputS7xD(321)(4) <= VNStageIntLLROutputS6xD(302)(5);
  CNStageIntLLRInputS7xD(8)(4) <= VNStageIntLLROutputS6xD(303)(0);
  CNStageIntLLRInputS7xD(102)(4) <= VNStageIntLLROutputS6xD(303)(1);
  CNStageIntLLRInputS7xD(112)(4) <= VNStageIntLLROutputS6xD(303)(2);
  CNStageIntLLRInputS7xD(178)(4) <= VNStageIntLLROutputS6xD(303)(3);
  CNStageIntLLRInputS7xD(235)(4) <= VNStageIntLLROutputS6xD(303)(4);
  CNStageIntLLRInputS7xD(293)(4) <= VNStageIntLLROutputS6xD(303)(5);
  CNStageIntLLRInputS7xD(382)(4) <= VNStageIntLLROutputS6xD(303)(6);
  CNStageIntLLRInputS7xD(7)(4) <= VNStageIntLLROutputS6xD(304)(0);
  CNStageIntLLRInputS7xD(97)(4) <= VNStageIntLLROutputS6xD(304)(1);
  CNStageIntLLRInputS7xD(157)(4) <= VNStageIntLLROutputS6xD(304)(2);
  CNStageIntLLRInputS7xD(222)(4) <= VNStageIntLLROutputS6xD(304)(3);
  CNStageIntLLRInputS7xD(263)(4) <= VNStageIntLLROutputS6xD(304)(4);
  CNStageIntLLRInputS7xD(283)(4) <= VNStageIntLLROutputS6xD(304)(5);
  CNStageIntLLRInputS7xD(359)(4) <= VNStageIntLLROutputS6xD(304)(6);
  CNStageIntLLRInputS7xD(6)(4) <= VNStageIntLLROutputS6xD(305)(0);
  CNStageIntLLRInputS7xD(80)(4) <= VNStageIntLLROutputS6xD(305)(1);
  CNStageIntLLRInputS7xD(115)(4) <= VNStageIntLLROutputS6xD(305)(2);
  CNStageIntLLRInputS7xD(209)(4) <= VNStageIntLLROutputS6xD(305)(3);
  CNStageIntLLRInputS7xD(276)(4) <= VNStageIntLLROutputS6xD(305)(4);
  CNStageIntLLRInputS7xD(323)(4) <= VNStageIntLLROutputS6xD(305)(5);
  CNStageIntLLRInputS7xD(342)(4) <= VNStageIntLLROutputS6xD(305)(6);
  CNStageIntLLRInputS7xD(5)(4) <= VNStageIntLLROutputS6xD(306)(0);
  CNStageIntLLRInputS7xD(87)(4) <= VNStageIntLLROutputS6xD(306)(1);
  CNStageIntLLRInputS7xD(136)(4) <= VNStageIntLLROutputS6xD(306)(2);
  CNStageIntLLRInputS7xD(174)(4) <= VNStageIntLLROutputS6xD(306)(3);
  CNStageIntLLRInputS7xD(4)(4) <= VNStageIntLLROutputS6xD(307)(0);
  CNStageIntLLRInputS7xD(107)(4) <= VNStageIntLLROutputS6xD(307)(1);
  CNStageIntLLRInputS7xD(145)(4) <= VNStageIntLLROutputS6xD(307)(2);
  CNStageIntLLRInputS7xD(202)(4) <= VNStageIntLLROutputS6xD(307)(3);
  CNStageIntLLRInputS7xD(230)(4) <= VNStageIntLLROutputS6xD(307)(4);
  CNStageIntLLRInputS7xD(302)(4) <= VNStageIntLLROutputS6xD(307)(5);
  CNStageIntLLRInputS7xD(366)(4) <= VNStageIntLLROutputS6xD(307)(6);
  CNStageIntLLRInputS7xD(140)(4) <= VNStageIntLLROutputS6xD(308)(0);
  CNStageIntLLRInputS7xD(199)(4) <= VNStageIntLLROutputS6xD(308)(1);
  CNStageIntLLRInputS7xD(251)(4) <= VNStageIntLLROutputS6xD(308)(2);
  CNStageIntLLRInputS7xD(311)(4) <= VNStageIntLLROutputS6xD(308)(3);
  CNStageIntLLRInputS7xD(336)(4) <= VNStageIntLLROutputS6xD(308)(4);
  CNStageIntLLRInputS7xD(3)(4) <= VNStageIntLLROutputS6xD(309)(0);
  CNStageIntLLRInputS7xD(86)(4) <= VNStageIntLLROutputS6xD(309)(1);
  CNStageIntLLRInputS7xD(146)(4) <= VNStageIntLLROutputS6xD(309)(2);
  CNStageIntLLRInputS7xD(214)(4) <= VNStageIntLLROutputS6xD(309)(3);
  CNStageIntLLRInputS7xD(265)(4) <= VNStageIntLLROutputS6xD(309)(4);
  CNStageIntLLRInputS7xD(307)(4) <= VNStageIntLLROutputS6xD(309)(5);
  CNStageIntLLRInputS7xD(2)(4) <= VNStageIntLLROutputS6xD(310)(0);
  CNStageIntLLRInputS7xD(65)(4) <= VNStageIntLLROutputS6xD(310)(1);
  CNStageIntLLRInputS7xD(135)(4) <= VNStageIntLLROutputS6xD(310)(2);
  CNStageIntLLRInputS7xD(261)(4) <= VNStageIntLLROutputS6xD(310)(3);
  CNStageIntLLRInputS7xD(312)(4) <= VNStageIntLLROutputS6xD(310)(4);
  CNStageIntLLRInputS7xD(369)(4) <= VNStageIntLLROutputS6xD(310)(5);
  CNStageIntLLRInputS7xD(1)(4) <= VNStageIntLLROutputS6xD(311)(0);
  CNStageIntLLRInputS7xD(68)(4) <= VNStageIntLLROutputS6xD(311)(1);
  CNStageIntLLRInputS7xD(160)(4) <= VNStageIntLLROutputS6xD(311)(2);
  CNStageIntLLRInputS7xD(225)(4) <= VNStageIntLLROutputS6xD(311)(3);
  CNStageIntLLRInputS7xD(301)(4) <= VNStageIntLLROutputS6xD(311)(4);
  CNStageIntLLRInputS7xD(0)(4) <= VNStageIntLLROutputS6xD(312)(0);
  CNStageIntLLRInputS7xD(108)(4) <= VNStageIntLLROutputS6xD(312)(1);
  CNStageIntLLRInputS7xD(167)(4) <= VNStageIntLLROutputS6xD(312)(2);
  CNStageIntLLRInputS7xD(246)(4) <= VNStageIntLLROutputS6xD(312)(3);
  CNStageIntLLRInputS7xD(326)(4) <= VNStageIntLLROutputS6xD(312)(4);
  CNStageIntLLRInputS7xD(348)(4) <= VNStageIntLLROutputS6xD(312)(5);
  CNStageIntLLRInputS7xD(150)(4) <= VNStageIntLLROutputS6xD(313)(0);
  CNStageIntLLRInputS7xD(188)(4) <= VNStageIntLLROutputS6xD(313)(1);
  CNStageIntLLRInputS7xD(247)(4) <= VNStageIntLLROutputS6xD(313)(2);
  CNStageIntLLRInputS7xD(356)(4) <= VNStageIntLLROutputS6xD(313)(3);
  CNStageIntLLRInputS7xD(191)(4) <= VNStageIntLLROutputS6xD(314)(0);
  CNStageIntLLRInputS7xD(278)(4) <= VNStageIntLLROutputS6xD(314)(1);
  CNStageIntLLRInputS7xD(316)(4) <= VNStageIntLLROutputS6xD(314)(2);
  CNStageIntLLRInputS7xD(352)(4) <= VNStageIntLLROutputS6xD(314)(3);
  CNStageIntLLRInputS7xD(78)(4) <= VNStageIntLLROutputS6xD(315)(0);
  CNStageIntLLRInputS7xD(119)(4) <= VNStageIntLLROutputS6xD(315)(1);
  CNStageIntLLRInputS7xD(183)(4) <= VNStageIntLLROutputS6xD(315)(2);
  CNStageIntLLRInputS7xD(271)(4) <= VNStageIntLLROutputS6xD(315)(3);
  CNStageIntLLRInputS7xD(318)(4) <= VNStageIntLLROutputS6xD(315)(4);
  CNStageIntLLRInputS7xD(357)(4) <= VNStageIntLLROutputS6xD(315)(5);
  CNStageIntLLRInputS7xD(61)(4) <= VNStageIntLLROutputS6xD(316)(0);
  CNStageIntLLRInputS7xD(158)(4) <= VNStageIntLLROutputS6xD(316)(1);
  CNStageIntLLRInputS7xD(234)(4) <= VNStageIntLLROutputS6xD(316)(2);
  CNStageIntLLRInputS7xD(288)(4) <= VNStageIntLLROutputS6xD(316)(3);
  CNStageIntLLRInputS7xD(347)(4) <= VNStageIntLLROutputS6xD(316)(4);
  CNStageIntLLRInputS7xD(88)(4) <= VNStageIntLLROutputS6xD(317)(0);
  CNStageIntLLRInputS7xD(238)(4) <= VNStageIntLLROutputS6xD(317)(1);
  CNStageIntLLRInputS7xD(324)(4) <= VNStageIntLLROutputS6xD(317)(2);
  CNStageIntLLRInputS7xD(372)(4) <= VNStageIntLLROutputS6xD(317)(3);
  CNStageIntLLRInputS7xD(120)(4) <= VNStageIntLLROutputS6xD(318)(0);
  CNStageIntLLRInputS7xD(210)(4) <= VNStageIntLLROutputS6xD(318)(1);
  CNStageIntLLRInputS7xD(279)(4) <= VNStageIntLLROutputS6xD(318)(2);
  CNStageIntLLRInputS7xD(379)(4) <= VNStageIntLLROutputS6xD(318)(3);
  CNStageIntLLRInputS7xD(52)(4) <= VNStageIntLLROutputS6xD(319)(0);
  CNStageIntLLRInputS7xD(66)(4) <= VNStageIntLLROutputS6xD(319)(1);
  CNStageIntLLRInputS7xD(151)(4) <= VNStageIntLLROutputS6xD(319)(2);
  CNStageIntLLRInputS7xD(221)(4) <= VNStageIntLLROutputS6xD(319)(3);
  CNStageIntLLRInputS7xD(237)(4) <= VNStageIntLLROutputS6xD(319)(4);
  CNStageIntLLRInputS7xD(289)(4) <= VNStageIntLLROutputS6xD(319)(5);
  CNStageIntLLRInputS7xD(361)(4) <= VNStageIntLLROutputS6xD(319)(6);
  CNStageIntLLRInputS7xD(53)(5) <= VNStageIntLLROutputS6xD(320)(0);
  CNStageIntLLRInputS7xD(126)(5) <= VNStageIntLLROutputS6xD(320)(1);
  CNStageIntLLRInputS7xD(196)(5) <= VNStageIntLLROutputS6xD(320)(2);
  CNStageIntLLRInputS7xD(295)(5) <= VNStageIntLLROutputS6xD(320)(3);
  CNStageIntLLRInputS7xD(338)(5) <= VNStageIntLLROutputS6xD(320)(4);
  CNStageIntLLRInputS7xD(51)(5) <= VNStageIntLLROutputS6xD(321)(0);
  CNStageIntLLRInputS7xD(65)(5) <= VNStageIntLLROutputS6xD(321)(1);
  CNStageIntLLRInputS7xD(150)(5) <= VNStageIntLLROutputS6xD(321)(2);
  CNStageIntLLRInputS7xD(220)(5) <= VNStageIntLLROutputS6xD(321)(3);
  CNStageIntLLRInputS7xD(236)(5) <= VNStageIntLLROutputS6xD(321)(4);
  CNStageIntLLRInputS7xD(288)(5) <= VNStageIntLLROutputS6xD(321)(5);
  CNStageIntLLRInputS7xD(360)(5) <= VNStageIntLLROutputS6xD(321)(6);
  CNStageIntLLRInputS7xD(50)(5) <= VNStageIntLLROutputS6xD(322)(0);
  CNStageIntLLRInputS7xD(84)(5) <= VNStageIntLLROutputS6xD(322)(1);
  CNStageIntLLRInputS7xD(165)(5) <= VNStageIntLLROutputS6xD(322)(2);
  CNStageIntLLRInputS7xD(231)(5) <= VNStageIntLLROutputS6xD(322)(3);
  CNStageIntLLRInputS7xD(316)(5) <= VNStageIntLLROutputS6xD(322)(4);
  CNStageIntLLRInputS7xD(362)(5) <= VNStageIntLLROutputS6xD(322)(5);
  CNStageIntLLRInputS7xD(56)(5) <= VNStageIntLLROutputS6xD(323)(0);
  CNStageIntLLRInputS7xD(136)(5) <= VNStageIntLLROutputS6xD(323)(1);
  CNStageIntLLRInputS7xD(184)(5) <= VNStageIntLLROutputS6xD(323)(2);
  CNStageIntLLRInputS7xD(268)(5) <= VNStageIntLLROutputS6xD(323)(3);
  CNStageIntLLRInputS7xD(330)(5) <= VNStageIntLLROutputS6xD(323)(4);
  CNStageIntLLRInputS7xD(49)(5) <= VNStageIntLLROutputS6xD(324)(0);
  CNStageIntLLRInputS7xD(109)(5) <= VNStageIntLLROutputS6xD(324)(1);
  CNStageIntLLRInputS7xD(113)(5) <= VNStageIntLLROutputS6xD(324)(2);
  CNStageIntLLRInputS7xD(223)(5) <= VNStageIntLLROutputS6xD(324)(3);
  CNStageIntLLRInputS7xD(273)(5) <= VNStageIntLLROutputS6xD(324)(4);
  CNStageIntLLRInputS7xD(302)(5) <= VNStageIntLLROutputS6xD(324)(5);
  CNStageIntLLRInputS7xD(369)(5) <= VNStageIntLLROutputS6xD(324)(6);
  CNStageIntLLRInputS7xD(48)(5) <= VNStageIntLLROutputS6xD(325)(0);
  CNStageIntLLRInputS7xD(70)(5) <= VNStageIntLLROutputS6xD(325)(1);
  CNStageIntLLRInputS7xD(137)(5) <= VNStageIntLLROutputS6xD(325)(2);
  CNStageIntLLRInputS7xD(185)(5) <= VNStageIntLLROutputS6xD(325)(3);
  CNStageIntLLRInputS7xD(242)(5) <= VNStageIntLLROutputS6xD(325)(4);
  CNStageIntLLRInputS7xD(284)(5) <= VNStageIntLLROutputS6xD(325)(5);
  CNStageIntLLRInputS7xD(382)(5) <= VNStageIntLLROutputS6xD(325)(6);
  CNStageIntLLRInputS7xD(47)(5) <= VNStageIntLLROutputS6xD(326)(0);
  CNStageIntLLRInputS7xD(62)(5) <= VNStageIntLLROutputS6xD(326)(1);
  CNStageIntLLRInputS7xD(203)(5) <= VNStageIntLLROutputS6xD(326)(2);
  CNStageIntLLRInputS7xD(241)(5) <= VNStageIntLLROutputS6xD(326)(3);
  CNStageIntLLRInputS7xD(304)(5) <= VNStageIntLLROutputS6xD(326)(4);
  CNStageIntLLRInputS7xD(46)(5) <= VNStageIntLLROutputS6xD(327)(0);
  CNStageIntLLRInputS7xD(94)(5) <= VNStageIntLLROutputS6xD(327)(1);
  CNStageIntLLRInputS7xD(148)(5) <= VNStageIntLLROutputS6xD(327)(2);
  CNStageIntLLRInputS7xD(211)(5) <= VNStageIntLLROutputS6xD(327)(3);
  CNStageIntLLRInputS7xD(272)(5) <= VNStageIntLLROutputS6xD(327)(4);
  CNStageIntLLRInputS7xD(318)(5) <= VNStageIntLLROutputS6xD(327)(5);
  CNStageIntLLRInputS7xD(361)(5) <= VNStageIntLLROutputS6xD(327)(6);
  CNStageIntLLRInputS7xD(45)(5) <= VNStageIntLLROutputS6xD(328)(0);
  CNStageIntLLRInputS7xD(103)(5) <= VNStageIntLLROutputS6xD(328)(1);
  CNStageIntLLRInputS7xD(168)(5) <= VNStageIntLLROutputS6xD(328)(2);
  CNStageIntLLRInputS7xD(314)(5) <= VNStageIntLLROutputS6xD(328)(3);
  CNStageIntLLRInputS7xD(377)(5) <= VNStageIntLLROutputS6xD(328)(4);
  CNStageIntLLRInputS7xD(44)(5) <= VNStageIntLLROutputS6xD(329)(0);
  CNStageIntLLRInputS7xD(97)(5) <= VNStageIntLLROutputS6xD(329)(1);
  CNStageIntLLRInputS7xD(131)(5) <= VNStageIntLLROutputS6xD(329)(2);
  CNStageIntLLRInputS7xD(212)(5) <= VNStageIntLLROutputS6xD(329)(3);
  CNStageIntLLRInputS7xD(255)(5) <= VNStageIntLLROutputS6xD(329)(4);
  CNStageIntLLRInputS7xD(280)(5) <= VNStageIntLLROutputS6xD(329)(5);
  CNStageIntLLRInputS7xD(348)(5) <= VNStageIntLLROutputS6xD(329)(6);
  CNStageIntLLRInputS7xD(43)(5) <= VNStageIntLLROutputS6xD(330)(0);
  CNStageIntLLRInputS7xD(101)(5) <= VNStageIntLLROutputS6xD(330)(1);
  CNStageIntLLRInputS7xD(132)(5) <= VNStageIntLLROutputS6xD(330)(2);
  CNStageIntLLRInputS7xD(202)(5) <= VNStageIntLLROutputS6xD(330)(3);
  CNStageIntLLRInputS7xD(243)(5) <= VNStageIntLLROutputS6xD(330)(4);
  CNStageIntLLRInputS7xD(42)(5) <= VNStageIntLLROutputS6xD(331)(0);
  CNStageIntLLRInputS7xD(92)(5) <= VNStageIntLLROutputS6xD(331)(1);
  CNStageIntLLRInputS7xD(167)(5) <= VNStageIntLLROutputS6xD(331)(2);
  CNStageIntLLRInputS7xD(172)(5) <= VNStageIntLLROutputS6xD(331)(3);
  CNStageIntLLRInputS7xD(350)(5) <= VNStageIntLLROutputS6xD(331)(4);
  CNStageIntLLRInputS7xD(41)(5) <= VNStageIntLLROutputS6xD(332)(0);
  CNStageIntLLRInputS7xD(71)(5) <= VNStageIntLLROutputS6xD(332)(1);
  CNStageIntLLRInputS7xD(158)(5) <= VNStageIntLLROutputS6xD(332)(2);
  CNStageIntLLRInputS7xD(179)(5) <= VNStageIntLLROutputS6xD(332)(3);
  CNStageIntLLRInputS7xD(240)(5) <= VNStageIntLLROutputS6xD(332)(4);
  CNStageIntLLRInputS7xD(363)(5) <= VNStageIntLLROutputS6xD(332)(5);
  CNStageIntLLRInputS7xD(108)(5) <= VNStageIntLLROutputS6xD(333)(0);
  CNStageIntLLRInputS7xD(117)(5) <= VNStageIntLLROutputS6xD(333)(1);
  CNStageIntLLRInputS7xD(215)(5) <= VNStageIntLLROutputS6xD(333)(2);
  CNStageIntLLRInputS7xD(265)(5) <= VNStageIntLLROutputS6xD(333)(3);
  CNStageIntLLRInputS7xD(324)(5) <= VNStageIntLLROutputS6xD(333)(4);
  CNStageIntLLRInputS7xD(359)(5) <= VNStageIntLLROutputS6xD(333)(5);
  CNStageIntLLRInputS7xD(40)(5) <= VNStageIntLLROutputS6xD(334)(0);
  CNStageIntLLRInputS7xD(66)(5) <= VNStageIntLLROutputS6xD(334)(1);
  CNStageIntLLRInputS7xD(217)(5) <= VNStageIntLLROutputS6xD(334)(2);
  CNStageIntLLRInputS7xD(286)(5) <= VNStageIntLLROutputS6xD(334)(3);
  CNStageIntLLRInputS7xD(380)(5) <= VNStageIntLLROutputS6xD(334)(4);
  CNStageIntLLRInputS7xD(39)(5) <= VNStageIntLLROutputS6xD(335)(0);
  CNStageIntLLRInputS7xD(78)(5) <= VNStageIntLLROutputS6xD(335)(1);
  CNStageIntLLRInputS7xD(170)(5) <= VNStageIntLLROutputS6xD(335)(2);
  CNStageIntLLRInputS7xD(189)(5) <= VNStageIntLLROutputS6xD(335)(3);
  CNStageIntLLRInputS7xD(274)(5) <= VNStageIntLLROutputS6xD(335)(4);
  CNStageIntLLRInputS7xD(291)(5) <= VNStageIntLLROutputS6xD(335)(5);
  CNStageIntLLRInputS7xD(343)(5) <= VNStageIntLLROutputS6xD(335)(6);
  CNStageIntLLRInputS7xD(38)(5) <= VNStageIntLLROutputS6xD(336)(0);
  CNStageIntLLRInputS7xD(104)(5) <= VNStageIntLLROutputS6xD(336)(1);
  CNStageIntLLRInputS7xD(121)(5) <= VNStageIntLLROutputS6xD(336)(2);
  CNStageIntLLRInputS7xD(267)(5) <= VNStageIntLLROutputS6xD(336)(3);
  CNStageIntLLRInputS7xD(332)(5) <= VNStageIntLLROutputS6xD(336)(4);
  CNStageIntLLRInputS7xD(344)(5) <= VNStageIntLLROutputS6xD(336)(5);
  CNStageIntLLRInputS7xD(37)(5) <= VNStageIntLLROutputS6xD(337)(0);
  CNStageIntLLRInputS7xD(93)(5) <= VNStageIntLLROutputS6xD(337)(1);
  CNStageIntLLRInputS7xD(115)(5) <= VNStageIntLLROutputS6xD(337)(2);
  CNStageIntLLRInputS7xD(183)(5) <= VNStageIntLLROutputS6xD(337)(3);
  CNStageIntLLRInputS7xD(253)(5) <= VNStageIntLLROutputS6xD(337)(4);
  CNStageIntLLRInputS7xD(290)(5) <= VNStageIntLLROutputS6xD(337)(5);
  CNStageIntLLRInputS7xD(379)(5) <= VNStageIntLLROutputS6xD(337)(6);
  CNStageIntLLRInputS7xD(36)(5) <= VNStageIntLLROutputS6xD(338)(0);
  CNStageIntLLRInputS7xD(80)(5) <= VNStageIntLLROutputS6xD(338)(1);
  CNStageIntLLRInputS7xD(155)(5) <= VNStageIntLLROutputS6xD(338)(2);
  CNStageIntLLRInputS7xD(190)(5) <= VNStageIntLLROutputS6xD(338)(3);
  CNStageIntLLRInputS7xD(370)(5) <= VNStageIntLLROutputS6xD(338)(4);
  CNStageIntLLRInputS7xD(35)(5) <= VNStageIntLLROutputS6xD(339)(0);
  CNStageIntLLRInputS7xD(96)(5) <= VNStageIntLLROutputS6xD(339)(1);
  CNStageIntLLRInputS7xD(163)(5) <= VNStageIntLLROutputS6xD(339)(2);
  CNStageIntLLRInputS7xD(216)(5) <= VNStageIntLLROutputS6xD(339)(3);
  CNStageIntLLRInputS7xD(247)(5) <= VNStageIntLLROutputS6xD(339)(4);
  CNStageIntLLRInputS7xD(322)(5) <= VNStageIntLLROutputS6xD(339)(5);
  CNStageIntLLRInputS7xD(34)(5) <= VNStageIntLLROutputS6xD(340)(0);
  CNStageIntLLRInputS7xD(58)(5) <= VNStageIntLLROutputS6xD(340)(1);
  CNStageIntLLRInputS7xD(127)(5) <= VNStageIntLLROutputS6xD(340)(2);
  CNStageIntLLRInputS7xD(178)(5) <= VNStageIntLLROutputS6xD(340)(3);
  CNStageIntLLRInputS7xD(245)(5) <= VNStageIntLLROutputS6xD(340)(4);
  CNStageIntLLRInputS7xD(334)(5) <= VNStageIntLLROutputS6xD(340)(5);
  CNStageIntLLRInputS7xD(33)(5) <= VNStageIntLLROutputS6xD(341)(0);
  CNStageIntLLRInputS7xD(68)(5) <= VNStageIntLLROutputS6xD(341)(1);
  CNStageIntLLRInputS7xD(125)(5) <= VNStageIntLLROutputS6xD(341)(2);
  CNStageIntLLRInputS7xD(204)(5) <= VNStageIntLLROutputS6xD(341)(3);
  CNStageIntLLRInputS7xD(258)(5) <= VNStageIntLLROutputS6xD(341)(4);
  CNStageIntLLRInputS7xD(296)(5) <= VNStageIntLLROutputS6xD(341)(5);
  CNStageIntLLRInputS7xD(32)(5) <= VNStageIntLLROutputS6xD(342)(0);
  CNStageIntLLRInputS7xD(63)(5) <= VNStageIntLLROutputS6xD(342)(1);
  CNStageIntLLRInputS7xD(161)(5) <= VNStageIntLLROutputS6xD(342)(2);
  CNStageIntLLRInputS7xD(251)(5) <= VNStageIntLLROutputS6xD(342)(3);
  CNStageIntLLRInputS7xD(294)(5) <= VNStageIntLLROutputS6xD(342)(4);
  CNStageIntLLRInputS7xD(31)(5) <= VNStageIntLLROutputS6xD(343)(0);
  CNStageIntLLRInputS7xD(69)(5) <= VNStageIntLLROutputS6xD(343)(1);
  CNStageIntLLRInputS7xD(140)(5) <= VNStageIntLLROutputS6xD(343)(2);
  CNStageIntLLRInputS7xD(206)(5) <= VNStageIntLLROutputS6xD(343)(3);
  CNStageIntLLRInputS7xD(228)(5) <= VNStageIntLLROutputS6xD(343)(4);
  CNStageIntLLRInputS7xD(327)(5) <= VNStageIntLLROutputS6xD(343)(5);
  CNStageIntLLRInputS7xD(30)(5) <= VNStageIntLLROutputS6xD(344)(0);
  CNStageIntLLRInputS7xD(57)(5) <= VNStageIntLLROutputS6xD(344)(1);
  CNStageIntLLRInputS7xD(143)(5) <= VNStageIntLLROutputS6xD(344)(2);
  CNStageIntLLRInputS7xD(218)(5) <= VNStageIntLLROutputS6xD(344)(3);
  CNStageIntLLRInputS7xD(238)(5) <= VNStageIntLLROutputS6xD(344)(4);
  CNStageIntLLRInputS7xD(307)(5) <= VNStageIntLLROutputS6xD(344)(5);
  CNStageIntLLRInputS7xD(367)(5) <= VNStageIntLLROutputS6xD(344)(6);
  CNStageIntLLRInputS7xD(29)(5) <= VNStageIntLLROutputS6xD(345)(0);
  CNStageIntLLRInputS7xD(83)(5) <= VNStageIntLLROutputS6xD(345)(1);
  CNStageIntLLRInputS7xD(128)(5) <= VNStageIntLLROutputS6xD(345)(2);
  CNStageIntLLRInputS7xD(232)(5) <= VNStageIntLLROutputS6xD(345)(3);
  CNStageIntLLRInputS7xD(309)(5) <= VNStageIntLLROutputS6xD(345)(4);
  CNStageIntLLRInputS7xD(375)(5) <= VNStageIntLLROutputS6xD(345)(5);
  CNStageIntLLRInputS7xD(28)(5) <= VNStageIntLLROutputS6xD(346)(0);
  CNStageIntLLRInputS7xD(89)(5) <= VNStageIntLLROutputS6xD(346)(1);
  CNStageIntLLRInputS7xD(162)(5) <= VNStageIntLLROutputS6xD(346)(2);
  CNStageIntLLRInputS7xD(181)(5) <= VNStageIntLLROutputS6xD(346)(3);
  CNStageIntLLRInputS7xD(235)(5) <= VNStageIntLLROutputS6xD(346)(4);
  CNStageIntLLRInputS7xD(297)(5) <= VNStageIntLLROutputS6xD(346)(5);
  CNStageIntLLRInputS7xD(339)(5) <= VNStageIntLLROutputS6xD(346)(6);
  CNStageIntLLRInputS7xD(27)(5) <= VNStageIntLLROutputS6xD(347)(0);
  CNStageIntLLRInputS7xD(73)(5) <= VNStageIntLLROutputS6xD(347)(1);
  CNStageIntLLRInputS7xD(124)(5) <= VNStageIntLLROutputS6xD(347)(2);
  CNStageIntLLRInputS7xD(199)(5) <= VNStageIntLLROutputS6xD(347)(3);
  CNStageIntLLRInputS7xD(225)(5) <= VNStageIntLLROutputS6xD(347)(4);
  CNStageIntLLRInputS7xD(328)(5) <= VNStageIntLLROutputS6xD(347)(5);
  CNStageIntLLRInputS7xD(337)(5) <= VNStageIntLLROutputS6xD(347)(6);
  CNStageIntLLRInputS7xD(26)(5) <= VNStageIntLLROutputS6xD(348)(0);
  CNStageIntLLRInputS7xD(75)(5) <= VNStageIntLLROutputS6xD(348)(1);
  CNStageIntLLRInputS7xD(152)(5) <= VNStageIntLLROutputS6xD(348)(2);
  CNStageIntLLRInputS7xD(200)(5) <= VNStageIntLLROutputS6xD(348)(3);
  CNStageIntLLRInputS7xD(259)(5) <= VNStageIntLLROutputS6xD(348)(4);
  CNStageIntLLRInputS7xD(293)(5) <= VNStageIntLLROutputS6xD(348)(5);
  CNStageIntLLRInputS7xD(373)(5) <= VNStageIntLLROutputS6xD(348)(6);
  CNStageIntLLRInputS7xD(25)(5) <= VNStageIntLLROutputS6xD(349)(0);
  CNStageIntLLRInputS7xD(99)(5) <= VNStageIntLLROutputS6xD(349)(1);
  CNStageIntLLRInputS7xD(180)(5) <= VNStageIntLLROutputS6xD(349)(2);
  CNStageIntLLRInputS7xD(244)(5) <= VNStageIntLLROutputS6xD(349)(3);
  CNStageIntLLRInputS7xD(319)(5) <= VNStageIntLLROutputS6xD(349)(4);
  CNStageIntLLRInputS7xD(352)(5) <= VNStageIntLLROutputS6xD(349)(5);
  CNStageIntLLRInputS7xD(24)(5) <= VNStageIntLLROutputS6xD(350)(0);
  CNStageIntLLRInputS7xD(81)(5) <= VNStageIntLLROutputS6xD(350)(1);
  CNStageIntLLRInputS7xD(164)(5) <= VNStageIntLLROutputS6xD(350)(2);
  CNStageIntLLRInputS7xD(171)(5) <= VNStageIntLLROutputS6xD(350)(3);
  CNStageIntLLRInputS7xD(254)(5) <= VNStageIntLLROutputS6xD(350)(4);
  CNStageIntLLRInputS7xD(303)(5) <= VNStageIntLLROutputS6xD(350)(5);
  CNStageIntLLRInputS7xD(23)(5) <= VNStageIntLLROutputS6xD(351)(0);
  CNStageIntLLRInputS7xD(154)(5) <= VNStageIntLLROutputS6xD(351)(1);
  CNStageIntLLRInputS7xD(188)(5) <= VNStageIntLLROutputS6xD(351)(2);
  CNStageIntLLRInputS7xD(266)(5) <= VNStageIntLLROutputS6xD(351)(3);
  CNStageIntLLRInputS7xD(329)(5) <= VNStageIntLLROutputS6xD(351)(4);
  CNStageIntLLRInputS7xD(340)(5) <= VNStageIntLLROutputS6xD(351)(5);
  CNStageIntLLRInputS7xD(22)(5) <= VNStageIntLLROutputS6xD(352)(0);
  CNStageIntLLRInputS7xD(100)(5) <= VNStageIntLLROutputS6xD(352)(1);
  CNStageIntLLRInputS7xD(141)(5) <= VNStageIntLLROutputS6xD(352)(2);
  CNStageIntLLRInputS7xD(192)(5) <= VNStageIntLLROutputS6xD(352)(3);
  CNStageIntLLRInputS7xD(239)(5) <= VNStageIntLLROutputS6xD(352)(4);
  CNStageIntLLRInputS7xD(321)(5) <= VNStageIntLLROutputS6xD(352)(5);
  CNStageIntLLRInputS7xD(374)(5) <= VNStageIntLLROutputS6xD(352)(6);
  CNStageIntLLRInputS7xD(21)(5) <= VNStageIntLLROutputS6xD(353)(0);
  CNStageIntLLRInputS7xD(74)(5) <= VNStageIntLLROutputS6xD(353)(1);
  CNStageIntLLRInputS7xD(160)(5) <= VNStageIntLLROutputS6xD(353)(2);
  CNStageIntLLRInputS7xD(224)(5) <= VNStageIntLLROutputS6xD(353)(3);
  CNStageIntLLRInputS7xD(227)(5) <= VNStageIntLLROutputS6xD(353)(4);
  CNStageIntLLRInputS7xD(336)(5) <= VNStageIntLLROutputS6xD(353)(5);
  CNStageIntLLRInputS7xD(20)(5) <= VNStageIntLLROutputS6xD(354)(0);
  CNStageIntLLRInputS7xD(88)(5) <= VNStageIntLLROutputS6xD(354)(1);
  CNStageIntLLRInputS7xD(133)(5) <= VNStageIntLLROutputS6xD(354)(2);
  CNStageIntLLRInputS7xD(191)(5) <= VNStageIntLLROutputS6xD(354)(3);
  CNStageIntLLRInputS7xD(326)(5) <= VNStageIntLLROutputS6xD(354)(4);
  CNStageIntLLRInputS7xD(364)(5) <= VNStageIntLLROutputS6xD(354)(5);
  CNStageIntLLRInputS7xD(19)(5) <= VNStageIntLLROutputS6xD(355)(0);
  CNStageIntLLRInputS7xD(59)(5) <= VNStageIntLLROutputS6xD(355)(1);
  CNStageIntLLRInputS7xD(130)(5) <= VNStageIntLLROutputS6xD(355)(2);
  CNStageIntLLRInputS7xD(186)(5) <= VNStageIntLLROutputS6xD(355)(3);
  CNStageIntLLRInputS7xD(230)(5) <= VNStageIntLLROutputS6xD(355)(4);
  CNStageIntLLRInputS7xD(300)(5) <= VNStageIntLLROutputS6xD(355)(5);
  CNStageIntLLRInputS7xD(349)(5) <= VNStageIntLLROutputS6xD(355)(6);
  CNStageIntLLRInputS7xD(18)(5) <= VNStageIntLLROutputS6xD(356)(0);
  CNStageIntLLRInputS7xD(95)(5) <= VNStageIntLLROutputS6xD(356)(1);
  CNStageIntLLRInputS7xD(146)(5) <= VNStageIntLLROutputS6xD(356)(2);
  CNStageIntLLRInputS7xD(222)(5) <= VNStageIntLLROutputS6xD(356)(3);
  CNStageIntLLRInputS7xD(299)(5) <= VNStageIntLLROutputS6xD(356)(4);
  CNStageIntLLRInputS7xD(376)(5) <= VNStageIntLLROutputS6xD(356)(5);
  CNStageIntLLRInputS7xD(17)(5) <= VNStageIntLLROutputS6xD(357)(0);
  CNStageIntLLRInputS7xD(61)(5) <= VNStageIntLLROutputS6xD(357)(1);
  CNStageIntLLRInputS7xD(138)(5) <= VNStageIntLLROutputS6xD(357)(2);
  CNStageIntLLRInputS7xD(176)(5) <= VNStageIntLLROutputS6xD(357)(3);
  CNStageIntLLRInputS7xD(256)(5) <= VNStageIntLLROutputS6xD(357)(4);
  CNStageIntLLRInputS7xD(312)(5) <= VNStageIntLLROutputS6xD(357)(5);
  CNStageIntLLRInputS7xD(366)(5) <= VNStageIntLLROutputS6xD(357)(6);
  CNStageIntLLRInputS7xD(16)(5) <= VNStageIntLLROutputS6xD(358)(0);
  CNStageIntLLRInputS7xD(76)(5) <= VNStageIntLLROutputS6xD(358)(1);
  CNStageIntLLRInputS7xD(112)(5) <= VNStageIntLLROutputS6xD(358)(2);
  CNStageIntLLRInputS7xD(252)(5) <= VNStageIntLLROutputS6xD(358)(3);
  CNStageIntLLRInputS7xD(305)(5) <= VNStageIntLLROutputS6xD(358)(4);
  CNStageIntLLRInputS7xD(353)(5) <= VNStageIntLLROutputS6xD(358)(5);
  CNStageIntLLRInputS7xD(15)(5) <= VNStageIntLLROutputS6xD(359)(0);
  CNStageIntLLRInputS7xD(72)(5) <= VNStageIntLLROutputS6xD(359)(1);
  CNStageIntLLRInputS7xD(122)(5) <= VNStageIntLLROutputS6xD(359)(2);
  CNStageIntLLRInputS7xD(195)(5) <= VNStageIntLLROutputS6xD(359)(3);
  CNStageIntLLRInputS7xD(257)(5) <= VNStageIntLLROutputS6xD(359)(4);
  CNStageIntLLRInputS7xD(283)(5) <= VNStageIntLLROutputS6xD(359)(5);
  CNStageIntLLRInputS7xD(372)(5) <= VNStageIntLLROutputS6xD(359)(6);
  CNStageIntLLRInputS7xD(14)(5) <= VNStageIntLLROutputS6xD(360)(0);
  CNStageIntLLRInputS7xD(91)(5) <= VNStageIntLLROutputS6xD(360)(1);
  CNStageIntLLRInputS7xD(116)(5) <= VNStageIntLLROutputS6xD(360)(2);
  CNStageIntLLRInputS7xD(174)(5) <= VNStageIntLLROutputS6xD(360)(3);
  CNStageIntLLRInputS7xD(248)(5) <= VNStageIntLLROutputS6xD(360)(4);
  CNStageIntLLRInputS7xD(292)(5) <= VNStageIntLLROutputS6xD(360)(5);
  CNStageIntLLRInputS7xD(345)(5) <= VNStageIntLLROutputS6xD(360)(6);
  CNStageIntLLRInputS7xD(13)(5) <= VNStageIntLLROutputS6xD(361)(0);
  CNStageIntLLRInputS7xD(54)(5) <= VNStageIntLLROutputS6xD(361)(1);
  CNStageIntLLRInputS7xD(120)(5) <= VNStageIntLLROutputS6xD(361)(2);
  CNStageIntLLRInputS7xD(207)(5) <= VNStageIntLLROutputS6xD(361)(3);
  CNStageIntLLRInputS7xD(271)(5) <= VNStageIntLLROutputS6xD(361)(4);
  CNStageIntLLRInputS7xD(285)(5) <= VNStageIntLLROutputS6xD(361)(5);
  CNStageIntLLRInputS7xD(342)(5) <= VNStageIntLLROutputS6xD(361)(6);
  CNStageIntLLRInputS7xD(12)(5) <= VNStageIntLLROutputS6xD(362)(0);
  CNStageIntLLRInputS7xD(55)(5) <= VNStageIntLLROutputS6xD(362)(1);
  CNStageIntLLRInputS7xD(169)(5) <= VNStageIntLLROutputS6xD(362)(2);
  CNStageIntLLRInputS7xD(210)(5) <= VNStageIntLLROutputS6xD(362)(3);
  CNStageIntLLRInputS7xD(276)(5) <= VNStageIntLLROutputS6xD(362)(4);
  CNStageIntLLRInputS7xD(289)(5) <= VNStageIntLLROutputS6xD(362)(5);
  CNStageIntLLRInputS7xD(357)(5) <= VNStageIntLLROutputS6xD(362)(6);
  CNStageIntLLRInputS7xD(90)(5) <= VNStageIntLLROutputS6xD(363)(0);
  CNStageIntLLRInputS7xD(147)(5) <= VNStageIntLLROutputS6xD(363)(1);
  CNStageIntLLRInputS7xD(197)(5) <= VNStageIntLLROutputS6xD(363)(2);
  CNStageIntLLRInputS7xD(261)(5) <= VNStageIntLLROutputS6xD(363)(3);
  CNStageIntLLRInputS7xD(281)(5) <= VNStageIntLLROutputS6xD(363)(4);
  CNStageIntLLRInputS7xD(11)(5) <= VNStageIntLLROutputS6xD(364)(0);
  CNStageIntLLRInputS7xD(82)(5) <= VNStageIntLLROutputS6xD(364)(1);
  CNStageIntLLRInputS7xD(129)(5) <= VNStageIntLLROutputS6xD(364)(2);
  CNStageIntLLRInputS7xD(175)(5) <= VNStageIntLLROutputS6xD(364)(3);
  CNStageIntLLRInputS7xD(263)(5) <= VNStageIntLLROutputS6xD(364)(4);
  CNStageIntLLRInputS7xD(313)(5) <= VNStageIntLLROutputS6xD(364)(5);
  CNStageIntLLRInputS7xD(10)(5) <= VNStageIntLLROutputS6xD(365)(0);
  CNStageIntLLRInputS7xD(98)(5) <= VNStageIntLLROutputS6xD(365)(1);
  CNStageIntLLRInputS7xD(142)(5) <= VNStageIntLLROutputS6xD(365)(2);
  CNStageIntLLRInputS7xD(194)(5) <= VNStageIntLLROutputS6xD(365)(3);
  CNStageIntLLRInputS7xD(234)(5) <= VNStageIntLLROutputS6xD(365)(4);
  CNStageIntLLRInputS7xD(298)(5) <= VNStageIntLLROutputS6xD(365)(5);
  CNStageIntLLRInputS7xD(9)(5) <= VNStageIntLLROutputS6xD(366)(0);
  CNStageIntLLRInputS7xD(102)(5) <= VNStageIntLLROutputS6xD(366)(1);
  CNStageIntLLRInputS7xD(153)(5) <= VNStageIntLLROutputS6xD(366)(2);
  CNStageIntLLRInputS7xD(219)(5) <= VNStageIntLLROutputS6xD(366)(3);
  CNStageIntLLRInputS7xD(269)(5) <= VNStageIntLLROutputS6xD(366)(4);
  CNStageIntLLRInputS7xD(308)(5) <= VNStageIntLLROutputS6xD(366)(5);
  CNStageIntLLRInputS7xD(8)(5) <= VNStageIntLLROutputS6xD(367)(0);
  CNStageIntLLRInputS7xD(110)(5) <= VNStageIntLLROutputS6xD(367)(1);
  CNStageIntLLRInputS7xD(123)(5) <= VNStageIntLLROutputS6xD(367)(2);
  CNStageIntLLRInputS7xD(205)(5) <= VNStageIntLLROutputS6xD(367)(3);
  CNStageIntLLRInputS7xD(226)(5) <= VNStageIntLLROutputS6xD(367)(4);
  CNStageIntLLRInputS7xD(320)(5) <= VNStageIntLLROutputS6xD(367)(5);
  CNStageIntLLRInputS7xD(333)(5) <= VNStageIntLLROutputS6xD(367)(6);
  CNStageIntLLRInputS7xD(7)(5) <= VNStageIntLLROutputS6xD(368)(0);
  CNStageIntLLRInputS7xD(177)(5) <= VNStageIntLLROutputS6xD(368)(1);
  CNStageIntLLRInputS7xD(381)(5) <= VNStageIntLLROutputS6xD(368)(2);
  CNStageIntLLRInputS7xD(6)(5) <= VNStageIntLLROutputS6xD(369)(0);
  CNStageIntLLRInputS7xD(156)(5) <= VNStageIntLLROutputS6xD(369)(1);
  CNStageIntLLRInputS7xD(221)(5) <= VNStageIntLLROutputS6xD(369)(2);
  CNStageIntLLRInputS7xD(262)(5) <= VNStageIntLLROutputS6xD(369)(3);
  CNStageIntLLRInputS7xD(358)(5) <= VNStageIntLLROutputS6xD(369)(4);
  CNStageIntLLRInputS7xD(5)(5) <= VNStageIntLLROutputS6xD(370)(0);
  CNStageIntLLRInputS7xD(114)(5) <= VNStageIntLLROutputS6xD(370)(1);
  CNStageIntLLRInputS7xD(208)(5) <= VNStageIntLLROutputS6xD(370)(2);
  CNStageIntLLRInputS7xD(275)(5) <= VNStageIntLLROutputS6xD(370)(3);
  CNStageIntLLRInputS7xD(341)(5) <= VNStageIntLLROutputS6xD(370)(4);
  CNStageIntLLRInputS7xD(4)(5) <= VNStageIntLLROutputS6xD(371)(0);
  CNStageIntLLRInputS7xD(135)(5) <= VNStageIntLLROutputS6xD(371)(1);
  CNStageIntLLRInputS7xD(173)(5) <= VNStageIntLLROutputS6xD(371)(2);
  CNStageIntLLRInputS7xD(249)(5) <= VNStageIntLLROutputS6xD(371)(3);
  CNStageIntLLRInputS7xD(354)(5) <= VNStageIntLLROutputS6xD(371)(4);
  CNStageIntLLRInputS7xD(106)(5) <= VNStageIntLLROutputS6xD(372)(0);
  CNStageIntLLRInputS7xD(144)(5) <= VNStageIntLLROutputS6xD(372)(1);
  CNStageIntLLRInputS7xD(201)(5) <= VNStageIntLLROutputS6xD(372)(2);
  CNStageIntLLRInputS7xD(229)(5) <= VNStageIntLLROutputS6xD(372)(3);
  CNStageIntLLRInputS7xD(301)(5) <= VNStageIntLLROutputS6xD(372)(4);
  CNStageIntLLRInputS7xD(365)(5) <= VNStageIntLLROutputS6xD(372)(5);
  CNStageIntLLRInputS7xD(3)(5) <= VNStageIntLLROutputS6xD(373)(0);
  CNStageIntLLRInputS7xD(139)(5) <= VNStageIntLLROutputS6xD(373)(1);
  CNStageIntLLRInputS7xD(250)(5) <= VNStageIntLLROutputS6xD(373)(2);
  CNStageIntLLRInputS7xD(310)(5) <= VNStageIntLLROutputS6xD(373)(3);
  CNStageIntLLRInputS7xD(335)(5) <= VNStageIntLLROutputS6xD(373)(4);
  CNStageIntLLRInputS7xD(2)(5) <= VNStageIntLLROutputS6xD(374)(0);
  CNStageIntLLRInputS7xD(85)(5) <= VNStageIntLLROutputS6xD(374)(1);
  CNStageIntLLRInputS7xD(145)(5) <= VNStageIntLLROutputS6xD(374)(2);
  CNStageIntLLRInputS7xD(213)(5) <= VNStageIntLLROutputS6xD(374)(3);
  CNStageIntLLRInputS7xD(264)(5) <= VNStageIntLLROutputS6xD(374)(4);
  CNStageIntLLRInputS7xD(306)(5) <= VNStageIntLLROutputS6xD(374)(5);
  CNStageIntLLRInputS7xD(383)(5) <= VNStageIntLLROutputS6xD(374)(6);
  CNStageIntLLRInputS7xD(1)(5) <= VNStageIntLLROutputS6xD(375)(0);
  CNStageIntLLRInputS7xD(64)(5) <= VNStageIntLLROutputS6xD(375)(1);
  CNStageIntLLRInputS7xD(134)(5) <= VNStageIntLLROutputS6xD(375)(2);
  CNStageIntLLRInputS7xD(260)(5) <= VNStageIntLLROutputS6xD(375)(3);
  CNStageIntLLRInputS7xD(311)(5) <= VNStageIntLLROutputS6xD(375)(4);
  CNStageIntLLRInputS7xD(368)(5) <= VNStageIntLLROutputS6xD(375)(5);
  CNStageIntLLRInputS7xD(0)(5) <= VNStageIntLLROutputS6xD(376)(0);
  CNStageIntLLRInputS7xD(67)(5) <= VNStageIntLLROutputS6xD(376)(1);
  CNStageIntLLRInputS7xD(159)(5) <= VNStageIntLLROutputS6xD(376)(2);
  CNStageIntLLRInputS7xD(278)(5) <= VNStageIntLLROutputS6xD(376)(3);
  CNStageIntLLRInputS7xD(107)(5) <= VNStageIntLLROutputS6xD(377)(0);
  CNStageIntLLRInputS7xD(166)(5) <= VNStageIntLLROutputS6xD(377)(1);
  CNStageIntLLRInputS7xD(193)(5) <= VNStageIntLLROutputS6xD(377)(2);
  CNStageIntLLRInputS7xD(325)(5) <= VNStageIntLLROutputS6xD(377)(3);
  CNStageIntLLRInputS7xD(347)(5) <= VNStageIntLLROutputS6xD(377)(4);
  CNStageIntLLRInputS7xD(86)(5) <= VNStageIntLLROutputS6xD(378)(0);
  CNStageIntLLRInputS7xD(149)(5) <= VNStageIntLLROutputS6xD(378)(1);
  CNStageIntLLRInputS7xD(187)(5) <= VNStageIntLLROutputS6xD(378)(2);
  CNStageIntLLRInputS7xD(246)(5) <= VNStageIntLLROutputS6xD(378)(3);
  CNStageIntLLRInputS7xD(331)(5) <= VNStageIntLLROutputS6xD(378)(4);
  CNStageIntLLRInputS7xD(355)(5) <= VNStageIntLLROutputS6xD(378)(5);
  CNStageIntLLRInputS7xD(105)(5) <= VNStageIntLLROutputS6xD(379)(0);
  CNStageIntLLRInputS7xD(151)(5) <= VNStageIntLLROutputS6xD(379)(1);
  CNStageIntLLRInputS7xD(277)(5) <= VNStageIntLLROutputS6xD(379)(2);
  CNStageIntLLRInputS7xD(315)(5) <= VNStageIntLLROutputS6xD(379)(3);
  CNStageIntLLRInputS7xD(351)(5) <= VNStageIntLLROutputS6xD(379)(4);
  CNStageIntLLRInputS7xD(77)(5) <= VNStageIntLLROutputS6xD(380)(0);
  CNStageIntLLRInputS7xD(118)(5) <= VNStageIntLLROutputS6xD(380)(1);
  CNStageIntLLRInputS7xD(182)(5) <= VNStageIntLLROutputS6xD(380)(2);
  CNStageIntLLRInputS7xD(270)(5) <= VNStageIntLLROutputS6xD(380)(3);
  CNStageIntLLRInputS7xD(317)(5) <= VNStageIntLLROutputS6xD(380)(4);
  CNStageIntLLRInputS7xD(356)(5) <= VNStageIntLLROutputS6xD(380)(5);
  CNStageIntLLRInputS7xD(60)(5) <= VNStageIntLLROutputS6xD(381)(0);
  CNStageIntLLRInputS7xD(157)(5) <= VNStageIntLLROutputS6xD(381)(1);
  CNStageIntLLRInputS7xD(214)(5) <= VNStageIntLLROutputS6xD(381)(2);
  CNStageIntLLRInputS7xD(233)(5) <= VNStageIntLLROutputS6xD(381)(3);
  CNStageIntLLRInputS7xD(287)(5) <= VNStageIntLLROutputS6xD(381)(4);
  CNStageIntLLRInputS7xD(346)(5) <= VNStageIntLLROutputS6xD(381)(5);
  CNStageIntLLRInputS7xD(87)(5) <= VNStageIntLLROutputS6xD(382)(0);
  CNStageIntLLRInputS7xD(111)(5) <= VNStageIntLLROutputS6xD(382)(1);
  CNStageIntLLRInputS7xD(198)(5) <= VNStageIntLLROutputS6xD(382)(2);
  CNStageIntLLRInputS7xD(237)(5) <= VNStageIntLLROutputS6xD(382)(3);
  CNStageIntLLRInputS7xD(323)(5) <= VNStageIntLLROutputS6xD(382)(4);
  CNStageIntLLRInputS7xD(371)(5) <= VNStageIntLLROutputS6xD(382)(5);
  CNStageIntLLRInputS7xD(52)(5) <= VNStageIntLLROutputS6xD(383)(0);
  CNStageIntLLRInputS7xD(79)(5) <= VNStageIntLLROutputS6xD(383)(1);
  CNStageIntLLRInputS7xD(119)(5) <= VNStageIntLLROutputS6xD(383)(2);
  CNStageIntLLRInputS7xD(209)(5) <= VNStageIntLLROutputS6xD(383)(3);
  CNStageIntLLRInputS7xD(279)(5) <= VNStageIntLLROutputS6xD(383)(4);
  CNStageIntLLRInputS7xD(282)(5) <= VNStageIntLLROutputS6xD(383)(5);
  CNStageIntLLRInputS7xD(378)(5) <= VNStageIntLLROutputS6xD(383)(6);

  -- Variable Nodes (Iteration 7)
  VNStageIntLLRInputS7xD(56)(0) <= CNStageIntLLROutputS7xD(0)(0);
  VNStageIntLLRInputS7xD(120)(0) <= CNStageIntLLROutputS7xD(0)(1);
  VNStageIntLLRInputS7xD(184)(0) <= CNStageIntLLROutputS7xD(0)(2);
  VNStageIntLLRInputS7xD(248)(0) <= CNStageIntLLROutputS7xD(0)(3);
  VNStageIntLLRInputS7xD(312)(0) <= CNStageIntLLROutputS7xD(0)(4);
  VNStageIntLLRInputS7xD(376)(0) <= CNStageIntLLROutputS7xD(0)(5);
  VNStageIntLLRInputS7xD(55)(0) <= CNStageIntLLROutputS7xD(1)(0);
  VNStageIntLLRInputS7xD(119)(0) <= CNStageIntLLROutputS7xD(1)(1);
  VNStageIntLLRInputS7xD(183)(0) <= CNStageIntLLROutputS7xD(1)(2);
  VNStageIntLLRInputS7xD(247)(0) <= CNStageIntLLROutputS7xD(1)(3);
  VNStageIntLLRInputS7xD(311)(0) <= CNStageIntLLROutputS7xD(1)(4);
  VNStageIntLLRInputS7xD(375)(0) <= CNStageIntLLROutputS7xD(1)(5);
  VNStageIntLLRInputS7xD(54)(0) <= CNStageIntLLROutputS7xD(2)(0);
  VNStageIntLLRInputS7xD(118)(0) <= CNStageIntLLROutputS7xD(2)(1);
  VNStageIntLLRInputS7xD(182)(0) <= CNStageIntLLROutputS7xD(2)(2);
  VNStageIntLLRInputS7xD(246)(0) <= CNStageIntLLROutputS7xD(2)(3);
  VNStageIntLLRInputS7xD(310)(0) <= CNStageIntLLROutputS7xD(2)(4);
  VNStageIntLLRInputS7xD(374)(0) <= CNStageIntLLROutputS7xD(2)(5);
  VNStageIntLLRInputS7xD(53)(0) <= CNStageIntLLROutputS7xD(3)(0);
  VNStageIntLLRInputS7xD(117)(0) <= CNStageIntLLROutputS7xD(3)(1);
  VNStageIntLLRInputS7xD(181)(0) <= CNStageIntLLROutputS7xD(3)(2);
  VNStageIntLLRInputS7xD(245)(0) <= CNStageIntLLROutputS7xD(3)(3);
  VNStageIntLLRInputS7xD(309)(0) <= CNStageIntLLROutputS7xD(3)(4);
  VNStageIntLLRInputS7xD(373)(0) <= CNStageIntLLROutputS7xD(3)(5);
  VNStageIntLLRInputS7xD(51)(0) <= CNStageIntLLROutputS7xD(4)(0);
  VNStageIntLLRInputS7xD(115)(0) <= CNStageIntLLROutputS7xD(4)(1);
  VNStageIntLLRInputS7xD(179)(0) <= CNStageIntLLROutputS7xD(4)(2);
  VNStageIntLLRInputS7xD(243)(0) <= CNStageIntLLROutputS7xD(4)(3);
  VNStageIntLLRInputS7xD(307)(0) <= CNStageIntLLROutputS7xD(4)(4);
  VNStageIntLLRInputS7xD(371)(0) <= CNStageIntLLROutputS7xD(4)(5);
  VNStageIntLLRInputS7xD(50)(0) <= CNStageIntLLROutputS7xD(5)(0);
  VNStageIntLLRInputS7xD(114)(0) <= CNStageIntLLROutputS7xD(5)(1);
  VNStageIntLLRInputS7xD(178)(0) <= CNStageIntLLROutputS7xD(5)(2);
  VNStageIntLLRInputS7xD(242)(0) <= CNStageIntLLROutputS7xD(5)(3);
  VNStageIntLLRInputS7xD(306)(0) <= CNStageIntLLROutputS7xD(5)(4);
  VNStageIntLLRInputS7xD(370)(0) <= CNStageIntLLROutputS7xD(5)(5);
  VNStageIntLLRInputS7xD(49)(0) <= CNStageIntLLROutputS7xD(6)(0);
  VNStageIntLLRInputS7xD(113)(0) <= CNStageIntLLROutputS7xD(6)(1);
  VNStageIntLLRInputS7xD(177)(0) <= CNStageIntLLROutputS7xD(6)(2);
  VNStageIntLLRInputS7xD(241)(0) <= CNStageIntLLROutputS7xD(6)(3);
  VNStageIntLLRInputS7xD(305)(0) <= CNStageIntLLROutputS7xD(6)(4);
  VNStageIntLLRInputS7xD(369)(0) <= CNStageIntLLROutputS7xD(6)(5);
  VNStageIntLLRInputS7xD(48)(0) <= CNStageIntLLROutputS7xD(7)(0);
  VNStageIntLLRInputS7xD(112)(0) <= CNStageIntLLROutputS7xD(7)(1);
  VNStageIntLLRInputS7xD(176)(0) <= CNStageIntLLROutputS7xD(7)(2);
  VNStageIntLLRInputS7xD(240)(0) <= CNStageIntLLROutputS7xD(7)(3);
  VNStageIntLLRInputS7xD(304)(0) <= CNStageIntLLROutputS7xD(7)(4);
  VNStageIntLLRInputS7xD(368)(0) <= CNStageIntLLROutputS7xD(7)(5);
  VNStageIntLLRInputS7xD(47)(0) <= CNStageIntLLROutputS7xD(8)(0);
  VNStageIntLLRInputS7xD(111)(0) <= CNStageIntLLROutputS7xD(8)(1);
  VNStageIntLLRInputS7xD(175)(0) <= CNStageIntLLROutputS7xD(8)(2);
  VNStageIntLLRInputS7xD(239)(0) <= CNStageIntLLROutputS7xD(8)(3);
  VNStageIntLLRInputS7xD(303)(0) <= CNStageIntLLROutputS7xD(8)(4);
  VNStageIntLLRInputS7xD(367)(0) <= CNStageIntLLROutputS7xD(8)(5);
  VNStageIntLLRInputS7xD(46)(0) <= CNStageIntLLROutputS7xD(9)(0);
  VNStageIntLLRInputS7xD(110)(0) <= CNStageIntLLROutputS7xD(9)(1);
  VNStageIntLLRInputS7xD(174)(0) <= CNStageIntLLROutputS7xD(9)(2);
  VNStageIntLLRInputS7xD(238)(0) <= CNStageIntLLROutputS7xD(9)(3);
  VNStageIntLLRInputS7xD(302)(0) <= CNStageIntLLROutputS7xD(9)(4);
  VNStageIntLLRInputS7xD(366)(0) <= CNStageIntLLROutputS7xD(9)(5);
  VNStageIntLLRInputS7xD(45)(0) <= CNStageIntLLROutputS7xD(10)(0);
  VNStageIntLLRInputS7xD(109)(0) <= CNStageIntLLROutputS7xD(10)(1);
  VNStageIntLLRInputS7xD(173)(0) <= CNStageIntLLROutputS7xD(10)(2);
  VNStageIntLLRInputS7xD(237)(0) <= CNStageIntLLROutputS7xD(10)(3);
  VNStageIntLLRInputS7xD(301)(0) <= CNStageIntLLROutputS7xD(10)(4);
  VNStageIntLLRInputS7xD(365)(0) <= CNStageIntLLROutputS7xD(10)(5);
  VNStageIntLLRInputS7xD(44)(0) <= CNStageIntLLROutputS7xD(11)(0);
  VNStageIntLLRInputS7xD(108)(0) <= CNStageIntLLROutputS7xD(11)(1);
  VNStageIntLLRInputS7xD(172)(0) <= CNStageIntLLROutputS7xD(11)(2);
  VNStageIntLLRInputS7xD(236)(0) <= CNStageIntLLROutputS7xD(11)(3);
  VNStageIntLLRInputS7xD(300)(0) <= CNStageIntLLROutputS7xD(11)(4);
  VNStageIntLLRInputS7xD(364)(0) <= CNStageIntLLROutputS7xD(11)(5);
  VNStageIntLLRInputS7xD(42)(0) <= CNStageIntLLROutputS7xD(12)(0);
  VNStageIntLLRInputS7xD(106)(0) <= CNStageIntLLROutputS7xD(12)(1);
  VNStageIntLLRInputS7xD(170)(0) <= CNStageIntLLROutputS7xD(12)(2);
  VNStageIntLLRInputS7xD(234)(0) <= CNStageIntLLROutputS7xD(12)(3);
  VNStageIntLLRInputS7xD(298)(0) <= CNStageIntLLROutputS7xD(12)(4);
  VNStageIntLLRInputS7xD(362)(0) <= CNStageIntLLROutputS7xD(12)(5);
  VNStageIntLLRInputS7xD(41)(0) <= CNStageIntLLROutputS7xD(13)(0);
  VNStageIntLLRInputS7xD(105)(0) <= CNStageIntLLROutputS7xD(13)(1);
  VNStageIntLLRInputS7xD(169)(0) <= CNStageIntLLROutputS7xD(13)(2);
  VNStageIntLLRInputS7xD(233)(0) <= CNStageIntLLROutputS7xD(13)(3);
  VNStageIntLLRInputS7xD(297)(0) <= CNStageIntLLROutputS7xD(13)(4);
  VNStageIntLLRInputS7xD(361)(0) <= CNStageIntLLROutputS7xD(13)(5);
  VNStageIntLLRInputS7xD(40)(0) <= CNStageIntLLROutputS7xD(14)(0);
  VNStageIntLLRInputS7xD(104)(0) <= CNStageIntLLROutputS7xD(14)(1);
  VNStageIntLLRInputS7xD(168)(0) <= CNStageIntLLROutputS7xD(14)(2);
  VNStageIntLLRInputS7xD(232)(0) <= CNStageIntLLROutputS7xD(14)(3);
  VNStageIntLLRInputS7xD(296)(0) <= CNStageIntLLROutputS7xD(14)(4);
  VNStageIntLLRInputS7xD(360)(0) <= CNStageIntLLROutputS7xD(14)(5);
  VNStageIntLLRInputS7xD(39)(0) <= CNStageIntLLROutputS7xD(15)(0);
  VNStageIntLLRInputS7xD(103)(0) <= CNStageIntLLROutputS7xD(15)(1);
  VNStageIntLLRInputS7xD(167)(0) <= CNStageIntLLROutputS7xD(15)(2);
  VNStageIntLLRInputS7xD(231)(0) <= CNStageIntLLROutputS7xD(15)(3);
  VNStageIntLLRInputS7xD(295)(0) <= CNStageIntLLROutputS7xD(15)(4);
  VNStageIntLLRInputS7xD(359)(0) <= CNStageIntLLROutputS7xD(15)(5);
  VNStageIntLLRInputS7xD(38)(0) <= CNStageIntLLROutputS7xD(16)(0);
  VNStageIntLLRInputS7xD(102)(0) <= CNStageIntLLROutputS7xD(16)(1);
  VNStageIntLLRInputS7xD(166)(0) <= CNStageIntLLROutputS7xD(16)(2);
  VNStageIntLLRInputS7xD(230)(0) <= CNStageIntLLROutputS7xD(16)(3);
  VNStageIntLLRInputS7xD(294)(0) <= CNStageIntLLROutputS7xD(16)(4);
  VNStageIntLLRInputS7xD(358)(0) <= CNStageIntLLROutputS7xD(16)(5);
  VNStageIntLLRInputS7xD(37)(0) <= CNStageIntLLROutputS7xD(17)(0);
  VNStageIntLLRInputS7xD(101)(0) <= CNStageIntLLROutputS7xD(17)(1);
  VNStageIntLLRInputS7xD(165)(0) <= CNStageIntLLROutputS7xD(17)(2);
  VNStageIntLLRInputS7xD(229)(0) <= CNStageIntLLROutputS7xD(17)(3);
  VNStageIntLLRInputS7xD(293)(0) <= CNStageIntLLROutputS7xD(17)(4);
  VNStageIntLLRInputS7xD(357)(0) <= CNStageIntLLROutputS7xD(17)(5);
  VNStageIntLLRInputS7xD(36)(0) <= CNStageIntLLROutputS7xD(18)(0);
  VNStageIntLLRInputS7xD(100)(0) <= CNStageIntLLROutputS7xD(18)(1);
  VNStageIntLLRInputS7xD(164)(0) <= CNStageIntLLROutputS7xD(18)(2);
  VNStageIntLLRInputS7xD(228)(0) <= CNStageIntLLROutputS7xD(18)(3);
  VNStageIntLLRInputS7xD(292)(0) <= CNStageIntLLROutputS7xD(18)(4);
  VNStageIntLLRInputS7xD(356)(0) <= CNStageIntLLROutputS7xD(18)(5);
  VNStageIntLLRInputS7xD(35)(0) <= CNStageIntLLROutputS7xD(19)(0);
  VNStageIntLLRInputS7xD(99)(0) <= CNStageIntLLROutputS7xD(19)(1);
  VNStageIntLLRInputS7xD(163)(0) <= CNStageIntLLROutputS7xD(19)(2);
  VNStageIntLLRInputS7xD(227)(0) <= CNStageIntLLROutputS7xD(19)(3);
  VNStageIntLLRInputS7xD(291)(0) <= CNStageIntLLROutputS7xD(19)(4);
  VNStageIntLLRInputS7xD(355)(0) <= CNStageIntLLROutputS7xD(19)(5);
  VNStageIntLLRInputS7xD(34)(0) <= CNStageIntLLROutputS7xD(20)(0);
  VNStageIntLLRInputS7xD(98)(0) <= CNStageIntLLROutputS7xD(20)(1);
  VNStageIntLLRInputS7xD(162)(0) <= CNStageIntLLROutputS7xD(20)(2);
  VNStageIntLLRInputS7xD(226)(0) <= CNStageIntLLROutputS7xD(20)(3);
  VNStageIntLLRInputS7xD(290)(0) <= CNStageIntLLROutputS7xD(20)(4);
  VNStageIntLLRInputS7xD(354)(0) <= CNStageIntLLROutputS7xD(20)(5);
  VNStageIntLLRInputS7xD(33)(0) <= CNStageIntLLROutputS7xD(21)(0);
  VNStageIntLLRInputS7xD(97)(0) <= CNStageIntLLROutputS7xD(21)(1);
  VNStageIntLLRInputS7xD(161)(0) <= CNStageIntLLROutputS7xD(21)(2);
  VNStageIntLLRInputS7xD(225)(0) <= CNStageIntLLROutputS7xD(21)(3);
  VNStageIntLLRInputS7xD(289)(0) <= CNStageIntLLROutputS7xD(21)(4);
  VNStageIntLLRInputS7xD(353)(0) <= CNStageIntLLROutputS7xD(21)(5);
  VNStageIntLLRInputS7xD(32)(0) <= CNStageIntLLROutputS7xD(22)(0);
  VNStageIntLLRInputS7xD(96)(0) <= CNStageIntLLROutputS7xD(22)(1);
  VNStageIntLLRInputS7xD(160)(0) <= CNStageIntLLROutputS7xD(22)(2);
  VNStageIntLLRInputS7xD(224)(0) <= CNStageIntLLROutputS7xD(22)(3);
  VNStageIntLLRInputS7xD(288)(0) <= CNStageIntLLROutputS7xD(22)(4);
  VNStageIntLLRInputS7xD(352)(0) <= CNStageIntLLROutputS7xD(22)(5);
  VNStageIntLLRInputS7xD(31)(0) <= CNStageIntLLROutputS7xD(23)(0);
  VNStageIntLLRInputS7xD(95)(0) <= CNStageIntLLROutputS7xD(23)(1);
  VNStageIntLLRInputS7xD(159)(0) <= CNStageIntLLROutputS7xD(23)(2);
  VNStageIntLLRInputS7xD(223)(0) <= CNStageIntLLROutputS7xD(23)(3);
  VNStageIntLLRInputS7xD(287)(0) <= CNStageIntLLROutputS7xD(23)(4);
  VNStageIntLLRInputS7xD(351)(0) <= CNStageIntLLROutputS7xD(23)(5);
  VNStageIntLLRInputS7xD(30)(0) <= CNStageIntLLROutputS7xD(24)(0);
  VNStageIntLLRInputS7xD(94)(0) <= CNStageIntLLROutputS7xD(24)(1);
  VNStageIntLLRInputS7xD(158)(0) <= CNStageIntLLROutputS7xD(24)(2);
  VNStageIntLLRInputS7xD(222)(0) <= CNStageIntLLROutputS7xD(24)(3);
  VNStageIntLLRInputS7xD(286)(0) <= CNStageIntLLROutputS7xD(24)(4);
  VNStageIntLLRInputS7xD(350)(0) <= CNStageIntLLROutputS7xD(24)(5);
  VNStageIntLLRInputS7xD(29)(0) <= CNStageIntLLROutputS7xD(25)(0);
  VNStageIntLLRInputS7xD(93)(0) <= CNStageIntLLROutputS7xD(25)(1);
  VNStageIntLLRInputS7xD(157)(0) <= CNStageIntLLROutputS7xD(25)(2);
  VNStageIntLLRInputS7xD(221)(0) <= CNStageIntLLROutputS7xD(25)(3);
  VNStageIntLLRInputS7xD(285)(0) <= CNStageIntLLROutputS7xD(25)(4);
  VNStageIntLLRInputS7xD(349)(0) <= CNStageIntLLROutputS7xD(25)(5);
  VNStageIntLLRInputS7xD(28)(0) <= CNStageIntLLROutputS7xD(26)(0);
  VNStageIntLLRInputS7xD(92)(0) <= CNStageIntLLROutputS7xD(26)(1);
  VNStageIntLLRInputS7xD(156)(0) <= CNStageIntLLROutputS7xD(26)(2);
  VNStageIntLLRInputS7xD(220)(0) <= CNStageIntLLROutputS7xD(26)(3);
  VNStageIntLLRInputS7xD(284)(0) <= CNStageIntLLROutputS7xD(26)(4);
  VNStageIntLLRInputS7xD(348)(0) <= CNStageIntLLROutputS7xD(26)(5);
  VNStageIntLLRInputS7xD(27)(0) <= CNStageIntLLROutputS7xD(27)(0);
  VNStageIntLLRInputS7xD(91)(0) <= CNStageIntLLROutputS7xD(27)(1);
  VNStageIntLLRInputS7xD(155)(0) <= CNStageIntLLROutputS7xD(27)(2);
  VNStageIntLLRInputS7xD(219)(0) <= CNStageIntLLROutputS7xD(27)(3);
  VNStageIntLLRInputS7xD(283)(0) <= CNStageIntLLROutputS7xD(27)(4);
  VNStageIntLLRInputS7xD(347)(0) <= CNStageIntLLROutputS7xD(27)(5);
  VNStageIntLLRInputS7xD(26)(0) <= CNStageIntLLROutputS7xD(28)(0);
  VNStageIntLLRInputS7xD(90)(0) <= CNStageIntLLROutputS7xD(28)(1);
  VNStageIntLLRInputS7xD(154)(0) <= CNStageIntLLROutputS7xD(28)(2);
  VNStageIntLLRInputS7xD(218)(0) <= CNStageIntLLROutputS7xD(28)(3);
  VNStageIntLLRInputS7xD(282)(0) <= CNStageIntLLROutputS7xD(28)(4);
  VNStageIntLLRInputS7xD(346)(0) <= CNStageIntLLROutputS7xD(28)(5);
  VNStageIntLLRInputS7xD(25)(0) <= CNStageIntLLROutputS7xD(29)(0);
  VNStageIntLLRInputS7xD(89)(0) <= CNStageIntLLROutputS7xD(29)(1);
  VNStageIntLLRInputS7xD(153)(0) <= CNStageIntLLROutputS7xD(29)(2);
  VNStageIntLLRInputS7xD(217)(0) <= CNStageIntLLROutputS7xD(29)(3);
  VNStageIntLLRInputS7xD(281)(0) <= CNStageIntLLROutputS7xD(29)(4);
  VNStageIntLLRInputS7xD(345)(0) <= CNStageIntLLROutputS7xD(29)(5);
  VNStageIntLLRInputS7xD(24)(0) <= CNStageIntLLROutputS7xD(30)(0);
  VNStageIntLLRInputS7xD(88)(0) <= CNStageIntLLROutputS7xD(30)(1);
  VNStageIntLLRInputS7xD(152)(0) <= CNStageIntLLROutputS7xD(30)(2);
  VNStageIntLLRInputS7xD(216)(0) <= CNStageIntLLROutputS7xD(30)(3);
  VNStageIntLLRInputS7xD(280)(0) <= CNStageIntLLROutputS7xD(30)(4);
  VNStageIntLLRInputS7xD(344)(0) <= CNStageIntLLROutputS7xD(30)(5);
  VNStageIntLLRInputS7xD(23)(0) <= CNStageIntLLROutputS7xD(31)(0);
  VNStageIntLLRInputS7xD(87)(0) <= CNStageIntLLROutputS7xD(31)(1);
  VNStageIntLLRInputS7xD(151)(0) <= CNStageIntLLROutputS7xD(31)(2);
  VNStageIntLLRInputS7xD(215)(0) <= CNStageIntLLROutputS7xD(31)(3);
  VNStageIntLLRInputS7xD(279)(0) <= CNStageIntLLROutputS7xD(31)(4);
  VNStageIntLLRInputS7xD(343)(0) <= CNStageIntLLROutputS7xD(31)(5);
  VNStageIntLLRInputS7xD(22)(0) <= CNStageIntLLROutputS7xD(32)(0);
  VNStageIntLLRInputS7xD(86)(0) <= CNStageIntLLROutputS7xD(32)(1);
  VNStageIntLLRInputS7xD(150)(0) <= CNStageIntLLROutputS7xD(32)(2);
  VNStageIntLLRInputS7xD(214)(0) <= CNStageIntLLROutputS7xD(32)(3);
  VNStageIntLLRInputS7xD(278)(0) <= CNStageIntLLROutputS7xD(32)(4);
  VNStageIntLLRInputS7xD(342)(0) <= CNStageIntLLROutputS7xD(32)(5);
  VNStageIntLLRInputS7xD(21)(0) <= CNStageIntLLROutputS7xD(33)(0);
  VNStageIntLLRInputS7xD(85)(0) <= CNStageIntLLROutputS7xD(33)(1);
  VNStageIntLLRInputS7xD(149)(0) <= CNStageIntLLROutputS7xD(33)(2);
  VNStageIntLLRInputS7xD(213)(0) <= CNStageIntLLROutputS7xD(33)(3);
  VNStageIntLLRInputS7xD(277)(0) <= CNStageIntLLROutputS7xD(33)(4);
  VNStageIntLLRInputS7xD(341)(0) <= CNStageIntLLROutputS7xD(33)(5);
  VNStageIntLLRInputS7xD(20)(0) <= CNStageIntLLROutputS7xD(34)(0);
  VNStageIntLLRInputS7xD(84)(0) <= CNStageIntLLROutputS7xD(34)(1);
  VNStageIntLLRInputS7xD(148)(0) <= CNStageIntLLROutputS7xD(34)(2);
  VNStageIntLLRInputS7xD(212)(0) <= CNStageIntLLROutputS7xD(34)(3);
  VNStageIntLLRInputS7xD(276)(0) <= CNStageIntLLROutputS7xD(34)(4);
  VNStageIntLLRInputS7xD(340)(0) <= CNStageIntLLROutputS7xD(34)(5);
  VNStageIntLLRInputS7xD(19)(0) <= CNStageIntLLROutputS7xD(35)(0);
  VNStageIntLLRInputS7xD(83)(0) <= CNStageIntLLROutputS7xD(35)(1);
  VNStageIntLLRInputS7xD(147)(0) <= CNStageIntLLROutputS7xD(35)(2);
  VNStageIntLLRInputS7xD(211)(0) <= CNStageIntLLROutputS7xD(35)(3);
  VNStageIntLLRInputS7xD(275)(0) <= CNStageIntLLROutputS7xD(35)(4);
  VNStageIntLLRInputS7xD(339)(0) <= CNStageIntLLROutputS7xD(35)(5);
  VNStageIntLLRInputS7xD(18)(0) <= CNStageIntLLROutputS7xD(36)(0);
  VNStageIntLLRInputS7xD(82)(0) <= CNStageIntLLROutputS7xD(36)(1);
  VNStageIntLLRInputS7xD(146)(0) <= CNStageIntLLROutputS7xD(36)(2);
  VNStageIntLLRInputS7xD(210)(0) <= CNStageIntLLROutputS7xD(36)(3);
  VNStageIntLLRInputS7xD(274)(0) <= CNStageIntLLROutputS7xD(36)(4);
  VNStageIntLLRInputS7xD(338)(0) <= CNStageIntLLROutputS7xD(36)(5);
  VNStageIntLLRInputS7xD(17)(0) <= CNStageIntLLROutputS7xD(37)(0);
  VNStageIntLLRInputS7xD(81)(0) <= CNStageIntLLROutputS7xD(37)(1);
  VNStageIntLLRInputS7xD(145)(0) <= CNStageIntLLROutputS7xD(37)(2);
  VNStageIntLLRInputS7xD(209)(0) <= CNStageIntLLROutputS7xD(37)(3);
  VNStageIntLLRInputS7xD(273)(0) <= CNStageIntLLROutputS7xD(37)(4);
  VNStageIntLLRInputS7xD(337)(0) <= CNStageIntLLROutputS7xD(37)(5);
  VNStageIntLLRInputS7xD(16)(0) <= CNStageIntLLROutputS7xD(38)(0);
  VNStageIntLLRInputS7xD(80)(0) <= CNStageIntLLROutputS7xD(38)(1);
  VNStageIntLLRInputS7xD(144)(0) <= CNStageIntLLROutputS7xD(38)(2);
  VNStageIntLLRInputS7xD(208)(0) <= CNStageIntLLROutputS7xD(38)(3);
  VNStageIntLLRInputS7xD(272)(0) <= CNStageIntLLROutputS7xD(38)(4);
  VNStageIntLLRInputS7xD(336)(0) <= CNStageIntLLROutputS7xD(38)(5);
  VNStageIntLLRInputS7xD(15)(0) <= CNStageIntLLROutputS7xD(39)(0);
  VNStageIntLLRInputS7xD(79)(0) <= CNStageIntLLROutputS7xD(39)(1);
  VNStageIntLLRInputS7xD(143)(0) <= CNStageIntLLROutputS7xD(39)(2);
  VNStageIntLLRInputS7xD(207)(0) <= CNStageIntLLROutputS7xD(39)(3);
  VNStageIntLLRInputS7xD(271)(0) <= CNStageIntLLROutputS7xD(39)(4);
  VNStageIntLLRInputS7xD(335)(0) <= CNStageIntLLROutputS7xD(39)(5);
  VNStageIntLLRInputS7xD(14)(0) <= CNStageIntLLROutputS7xD(40)(0);
  VNStageIntLLRInputS7xD(78)(0) <= CNStageIntLLROutputS7xD(40)(1);
  VNStageIntLLRInputS7xD(142)(0) <= CNStageIntLLROutputS7xD(40)(2);
  VNStageIntLLRInputS7xD(206)(0) <= CNStageIntLLROutputS7xD(40)(3);
  VNStageIntLLRInputS7xD(270)(0) <= CNStageIntLLROutputS7xD(40)(4);
  VNStageIntLLRInputS7xD(334)(0) <= CNStageIntLLROutputS7xD(40)(5);
  VNStageIntLLRInputS7xD(12)(0) <= CNStageIntLLROutputS7xD(41)(0);
  VNStageIntLLRInputS7xD(76)(0) <= CNStageIntLLROutputS7xD(41)(1);
  VNStageIntLLRInputS7xD(140)(0) <= CNStageIntLLROutputS7xD(41)(2);
  VNStageIntLLRInputS7xD(204)(0) <= CNStageIntLLROutputS7xD(41)(3);
  VNStageIntLLRInputS7xD(268)(0) <= CNStageIntLLROutputS7xD(41)(4);
  VNStageIntLLRInputS7xD(332)(0) <= CNStageIntLLROutputS7xD(41)(5);
  VNStageIntLLRInputS7xD(11)(0) <= CNStageIntLLROutputS7xD(42)(0);
  VNStageIntLLRInputS7xD(75)(0) <= CNStageIntLLROutputS7xD(42)(1);
  VNStageIntLLRInputS7xD(139)(0) <= CNStageIntLLROutputS7xD(42)(2);
  VNStageIntLLRInputS7xD(203)(0) <= CNStageIntLLROutputS7xD(42)(3);
  VNStageIntLLRInputS7xD(267)(0) <= CNStageIntLLROutputS7xD(42)(4);
  VNStageIntLLRInputS7xD(331)(0) <= CNStageIntLLROutputS7xD(42)(5);
  VNStageIntLLRInputS7xD(10)(0) <= CNStageIntLLROutputS7xD(43)(0);
  VNStageIntLLRInputS7xD(74)(0) <= CNStageIntLLROutputS7xD(43)(1);
  VNStageIntLLRInputS7xD(138)(0) <= CNStageIntLLROutputS7xD(43)(2);
  VNStageIntLLRInputS7xD(202)(0) <= CNStageIntLLROutputS7xD(43)(3);
  VNStageIntLLRInputS7xD(266)(0) <= CNStageIntLLROutputS7xD(43)(4);
  VNStageIntLLRInputS7xD(330)(0) <= CNStageIntLLROutputS7xD(43)(5);
  VNStageIntLLRInputS7xD(9)(0) <= CNStageIntLLROutputS7xD(44)(0);
  VNStageIntLLRInputS7xD(73)(0) <= CNStageIntLLROutputS7xD(44)(1);
  VNStageIntLLRInputS7xD(137)(0) <= CNStageIntLLROutputS7xD(44)(2);
  VNStageIntLLRInputS7xD(201)(0) <= CNStageIntLLROutputS7xD(44)(3);
  VNStageIntLLRInputS7xD(265)(0) <= CNStageIntLLROutputS7xD(44)(4);
  VNStageIntLLRInputS7xD(329)(0) <= CNStageIntLLROutputS7xD(44)(5);
  VNStageIntLLRInputS7xD(8)(0) <= CNStageIntLLROutputS7xD(45)(0);
  VNStageIntLLRInputS7xD(72)(0) <= CNStageIntLLROutputS7xD(45)(1);
  VNStageIntLLRInputS7xD(136)(0) <= CNStageIntLLROutputS7xD(45)(2);
  VNStageIntLLRInputS7xD(200)(0) <= CNStageIntLLROutputS7xD(45)(3);
  VNStageIntLLRInputS7xD(264)(0) <= CNStageIntLLROutputS7xD(45)(4);
  VNStageIntLLRInputS7xD(328)(0) <= CNStageIntLLROutputS7xD(45)(5);
  VNStageIntLLRInputS7xD(7)(0) <= CNStageIntLLROutputS7xD(46)(0);
  VNStageIntLLRInputS7xD(71)(0) <= CNStageIntLLROutputS7xD(46)(1);
  VNStageIntLLRInputS7xD(135)(0) <= CNStageIntLLROutputS7xD(46)(2);
  VNStageIntLLRInputS7xD(199)(0) <= CNStageIntLLROutputS7xD(46)(3);
  VNStageIntLLRInputS7xD(263)(0) <= CNStageIntLLROutputS7xD(46)(4);
  VNStageIntLLRInputS7xD(327)(0) <= CNStageIntLLROutputS7xD(46)(5);
  VNStageIntLLRInputS7xD(6)(0) <= CNStageIntLLROutputS7xD(47)(0);
  VNStageIntLLRInputS7xD(70)(0) <= CNStageIntLLROutputS7xD(47)(1);
  VNStageIntLLRInputS7xD(134)(0) <= CNStageIntLLROutputS7xD(47)(2);
  VNStageIntLLRInputS7xD(198)(0) <= CNStageIntLLROutputS7xD(47)(3);
  VNStageIntLLRInputS7xD(262)(0) <= CNStageIntLLROutputS7xD(47)(4);
  VNStageIntLLRInputS7xD(326)(0) <= CNStageIntLLROutputS7xD(47)(5);
  VNStageIntLLRInputS7xD(5)(0) <= CNStageIntLLROutputS7xD(48)(0);
  VNStageIntLLRInputS7xD(69)(0) <= CNStageIntLLROutputS7xD(48)(1);
  VNStageIntLLRInputS7xD(133)(0) <= CNStageIntLLROutputS7xD(48)(2);
  VNStageIntLLRInputS7xD(197)(0) <= CNStageIntLLROutputS7xD(48)(3);
  VNStageIntLLRInputS7xD(261)(0) <= CNStageIntLLROutputS7xD(48)(4);
  VNStageIntLLRInputS7xD(325)(0) <= CNStageIntLLROutputS7xD(48)(5);
  VNStageIntLLRInputS7xD(4)(0) <= CNStageIntLLROutputS7xD(49)(0);
  VNStageIntLLRInputS7xD(68)(0) <= CNStageIntLLROutputS7xD(49)(1);
  VNStageIntLLRInputS7xD(132)(0) <= CNStageIntLLROutputS7xD(49)(2);
  VNStageIntLLRInputS7xD(196)(0) <= CNStageIntLLROutputS7xD(49)(3);
  VNStageIntLLRInputS7xD(260)(0) <= CNStageIntLLROutputS7xD(49)(4);
  VNStageIntLLRInputS7xD(324)(0) <= CNStageIntLLROutputS7xD(49)(5);
  VNStageIntLLRInputS7xD(2)(0) <= CNStageIntLLROutputS7xD(50)(0);
  VNStageIntLLRInputS7xD(66)(0) <= CNStageIntLLROutputS7xD(50)(1);
  VNStageIntLLRInputS7xD(130)(0) <= CNStageIntLLROutputS7xD(50)(2);
  VNStageIntLLRInputS7xD(194)(0) <= CNStageIntLLROutputS7xD(50)(3);
  VNStageIntLLRInputS7xD(258)(0) <= CNStageIntLLROutputS7xD(50)(4);
  VNStageIntLLRInputS7xD(322)(0) <= CNStageIntLLROutputS7xD(50)(5);
  VNStageIntLLRInputS7xD(1)(0) <= CNStageIntLLROutputS7xD(51)(0);
  VNStageIntLLRInputS7xD(65)(0) <= CNStageIntLLROutputS7xD(51)(1);
  VNStageIntLLRInputS7xD(129)(0) <= CNStageIntLLROutputS7xD(51)(2);
  VNStageIntLLRInputS7xD(193)(0) <= CNStageIntLLROutputS7xD(51)(3);
  VNStageIntLLRInputS7xD(257)(0) <= CNStageIntLLROutputS7xD(51)(4);
  VNStageIntLLRInputS7xD(321)(0) <= CNStageIntLLROutputS7xD(51)(5);
  VNStageIntLLRInputS7xD(63)(0) <= CNStageIntLLROutputS7xD(52)(0);
  VNStageIntLLRInputS7xD(127)(0) <= CNStageIntLLROutputS7xD(52)(1);
  VNStageIntLLRInputS7xD(191)(0) <= CNStageIntLLROutputS7xD(52)(2);
  VNStageIntLLRInputS7xD(255)(0) <= CNStageIntLLROutputS7xD(52)(3);
  VNStageIntLLRInputS7xD(319)(0) <= CNStageIntLLROutputS7xD(52)(4);
  VNStageIntLLRInputS7xD(383)(0) <= CNStageIntLLROutputS7xD(52)(5);
  VNStageIntLLRInputS7xD(0)(0) <= CNStageIntLLROutputS7xD(53)(0);
  VNStageIntLLRInputS7xD(64)(0) <= CNStageIntLLROutputS7xD(53)(1);
  VNStageIntLLRInputS7xD(128)(0) <= CNStageIntLLROutputS7xD(53)(2);
  VNStageIntLLRInputS7xD(192)(0) <= CNStageIntLLROutputS7xD(53)(3);
  VNStageIntLLRInputS7xD(256)(0) <= CNStageIntLLROutputS7xD(53)(4);
  VNStageIntLLRInputS7xD(320)(0) <= CNStageIntLLROutputS7xD(53)(5);
  VNStageIntLLRInputS7xD(42)(1) <= CNStageIntLLROutputS7xD(54)(0);
  VNStageIntLLRInputS7xD(112)(1) <= CNStageIntLLROutputS7xD(54)(1);
  VNStageIntLLRInputS7xD(182)(1) <= CNStageIntLLROutputS7xD(54)(2);
  VNStageIntLLRInputS7xD(203)(1) <= CNStageIntLLROutputS7xD(54)(3);
  VNStageIntLLRInputS7xD(259)(0) <= CNStageIntLLROutputS7xD(54)(4);
  VNStageIntLLRInputS7xD(361)(1) <= CNStageIntLLROutputS7xD(54)(5);
  VNStageIntLLRInputS7xD(41)(1) <= CNStageIntLLROutputS7xD(55)(0);
  VNStageIntLLRInputS7xD(117)(1) <= CNStageIntLLROutputS7xD(55)(1);
  VNStageIntLLRInputS7xD(138)(1) <= CNStageIntLLROutputS7xD(55)(2);
  VNStageIntLLRInputS7xD(194)(1) <= CNStageIntLLROutputS7xD(55)(3);
  VNStageIntLLRInputS7xD(296)(1) <= CNStageIntLLROutputS7xD(55)(4);
  VNStageIntLLRInputS7xD(362)(1) <= CNStageIntLLROutputS7xD(55)(5);
  VNStageIntLLRInputS7xD(40)(1) <= CNStageIntLLROutputS7xD(56)(0);
  VNStageIntLLRInputS7xD(73)(1) <= CNStageIntLLROutputS7xD(56)(1);
  VNStageIntLLRInputS7xD(129)(1) <= CNStageIntLLROutputS7xD(56)(2);
  VNStageIntLLRInputS7xD(231)(1) <= CNStageIntLLROutputS7xD(56)(3);
  VNStageIntLLRInputS7xD(297)(1) <= CNStageIntLLROutputS7xD(56)(4);
  VNStageIntLLRInputS7xD(323)(0) <= CNStageIntLLROutputS7xD(56)(5);
  VNStageIntLLRInputS7xD(39)(1) <= CNStageIntLLROutputS7xD(57)(0);
  VNStageIntLLRInputS7xD(127)(1) <= CNStageIntLLROutputS7xD(57)(1);
  VNStageIntLLRInputS7xD(166)(1) <= CNStageIntLLROutputS7xD(57)(2);
  VNStageIntLLRInputS7xD(232)(1) <= CNStageIntLLROutputS7xD(57)(3);
  VNStageIntLLRInputS7xD(258)(1) <= CNStageIntLLROutputS7xD(57)(4);
  VNStageIntLLRInputS7xD(344)(1) <= CNStageIntLLROutputS7xD(57)(5);
  VNStageIntLLRInputS7xD(38)(1) <= CNStageIntLLROutputS7xD(58)(0);
  VNStageIntLLRInputS7xD(101)(1) <= CNStageIntLLROutputS7xD(58)(1);
  VNStageIntLLRInputS7xD(167)(1) <= CNStageIntLLROutputS7xD(58)(2);
  VNStageIntLLRInputS7xD(193)(1) <= CNStageIntLLROutputS7xD(58)(3);
  VNStageIntLLRInputS7xD(279)(1) <= CNStageIntLLROutputS7xD(58)(4);
  VNStageIntLLRInputS7xD(340)(1) <= CNStageIntLLROutputS7xD(58)(5);
  VNStageIntLLRInputS7xD(37)(1) <= CNStageIntLLROutputS7xD(59)(0);
  VNStageIntLLRInputS7xD(102)(1) <= CNStageIntLLROutputS7xD(59)(1);
  VNStageIntLLRInputS7xD(191)(1) <= CNStageIntLLROutputS7xD(59)(2);
  VNStageIntLLRInputS7xD(214)(1) <= CNStageIntLLROutputS7xD(59)(3);
  VNStageIntLLRInputS7xD(275)(1) <= CNStageIntLLROutputS7xD(59)(4);
  VNStageIntLLRInputS7xD(355)(1) <= CNStageIntLLROutputS7xD(59)(5);
  VNStageIntLLRInputS7xD(36)(1) <= CNStageIntLLROutputS7xD(60)(0);
  VNStageIntLLRInputS7xD(126)(0) <= CNStageIntLLROutputS7xD(60)(1);
  VNStageIntLLRInputS7xD(149)(1) <= CNStageIntLLROutputS7xD(60)(2);
  VNStageIntLLRInputS7xD(210)(1) <= CNStageIntLLROutputS7xD(60)(3);
  VNStageIntLLRInputS7xD(290)(1) <= CNStageIntLLROutputS7xD(60)(4);
  VNStageIntLLRInputS7xD(381)(0) <= CNStageIntLLROutputS7xD(60)(5);
  VNStageIntLLRInputS7xD(35)(1) <= CNStageIntLLROutputS7xD(61)(0);
  VNStageIntLLRInputS7xD(84)(1) <= CNStageIntLLROutputS7xD(61)(1);
  VNStageIntLLRInputS7xD(145)(1) <= CNStageIntLLROutputS7xD(61)(2);
  VNStageIntLLRInputS7xD(225)(1) <= CNStageIntLLROutputS7xD(61)(3);
  VNStageIntLLRInputS7xD(316)(0) <= CNStageIntLLROutputS7xD(61)(4);
  VNStageIntLLRInputS7xD(357)(1) <= CNStageIntLLROutputS7xD(61)(5);
  VNStageIntLLRInputS7xD(34)(1) <= CNStageIntLLROutputS7xD(62)(0);
  VNStageIntLLRInputS7xD(80)(1) <= CNStageIntLLROutputS7xD(62)(1);
  VNStageIntLLRInputS7xD(160)(1) <= CNStageIntLLROutputS7xD(62)(2);
  VNStageIntLLRInputS7xD(251)(0) <= CNStageIntLLROutputS7xD(62)(3);
  VNStageIntLLRInputS7xD(292)(1) <= CNStageIntLLROutputS7xD(62)(4);
  VNStageIntLLRInputS7xD(326)(1) <= CNStageIntLLROutputS7xD(62)(5);
  VNStageIntLLRInputS7xD(33)(1) <= CNStageIntLLROutputS7xD(63)(0);
  VNStageIntLLRInputS7xD(95)(1) <= CNStageIntLLROutputS7xD(63)(1);
  VNStageIntLLRInputS7xD(186)(0) <= CNStageIntLLROutputS7xD(63)(2);
  VNStageIntLLRInputS7xD(227)(1) <= CNStageIntLLROutputS7xD(63)(3);
  VNStageIntLLRInputS7xD(261)(1) <= CNStageIntLLROutputS7xD(63)(4);
  VNStageIntLLRInputS7xD(342)(1) <= CNStageIntLLROutputS7xD(63)(5);
  VNStageIntLLRInputS7xD(32)(1) <= CNStageIntLLROutputS7xD(64)(0);
  VNStageIntLLRInputS7xD(121)(0) <= CNStageIntLLROutputS7xD(64)(1);
  VNStageIntLLRInputS7xD(162)(1) <= CNStageIntLLROutputS7xD(64)(2);
  VNStageIntLLRInputS7xD(196)(1) <= CNStageIntLLROutputS7xD(64)(3);
  VNStageIntLLRInputS7xD(277)(1) <= CNStageIntLLROutputS7xD(64)(4);
  VNStageIntLLRInputS7xD(375)(1) <= CNStageIntLLROutputS7xD(64)(5);
  VNStageIntLLRInputS7xD(31)(1) <= CNStageIntLLROutputS7xD(65)(0);
  VNStageIntLLRInputS7xD(97)(1) <= CNStageIntLLROutputS7xD(65)(1);
  VNStageIntLLRInputS7xD(131)(0) <= CNStageIntLLROutputS7xD(65)(2);
  VNStageIntLLRInputS7xD(212)(1) <= CNStageIntLLROutputS7xD(65)(3);
  VNStageIntLLRInputS7xD(310)(1) <= CNStageIntLLROutputS7xD(65)(4);
  VNStageIntLLRInputS7xD(321)(1) <= CNStageIntLLROutputS7xD(65)(5);
  VNStageIntLLRInputS7xD(30)(1) <= CNStageIntLLROutputS7xD(66)(0);
  VNStageIntLLRInputS7xD(66)(1) <= CNStageIntLLROutputS7xD(66)(1);
  VNStageIntLLRInputS7xD(147)(1) <= CNStageIntLLROutputS7xD(66)(2);
  VNStageIntLLRInputS7xD(245)(1) <= CNStageIntLLROutputS7xD(66)(3);
  VNStageIntLLRInputS7xD(319)(1) <= CNStageIntLLROutputS7xD(66)(4);
  VNStageIntLLRInputS7xD(334)(1) <= CNStageIntLLROutputS7xD(66)(5);
  VNStageIntLLRInputS7xD(29)(1) <= CNStageIntLLROutputS7xD(67)(0);
  VNStageIntLLRInputS7xD(82)(1) <= CNStageIntLLROutputS7xD(67)(1);
  VNStageIntLLRInputS7xD(180)(0) <= CNStageIntLLROutputS7xD(67)(2);
  VNStageIntLLRInputS7xD(254)(0) <= CNStageIntLLROutputS7xD(67)(3);
  VNStageIntLLRInputS7xD(269)(0) <= CNStageIntLLROutputS7xD(67)(4);
  VNStageIntLLRInputS7xD(376)(1) <= CNStageIntLLROutputS7xD(67)(5);
  VNStageIntLLRInputS7xD(28)(1) <= CNStageIntLLROutputS7xD(68)(0);
  VNStageIntLLRInputS7xD(115)(1) <= CNStageIntLLROutputS7xD(68)(1);
  VNStageIntLLRInputS7xD(189)(0) <= CNStageIntLLROutputS7xD(68)(2);
  VNStageIntLLRInputS7xD(204)(1) <= CNStageIntLLROutputS7xD(68)(3);
  VNStageIntLLRInputS7xD(311)(1) <= CNStageIntLLROutputS7xD(68)(4);
  VNStageIntLLRInputS7xD(341)(1) <= CNStageIntLLROutputS7xD(68)(5);
  VNStageIntLLRInputS7xD(27)(1) <= CNStageIntLLROutputS7xD(69)(0);
  VNStageIntLLRInputS7xD(124)(0) <= CNStageIntLLROutputS7xD(69)(1);
  VNStageIntLLRInputS7xD(139)(1) <= CNStageIntLLROutputS7xD(69)(2);
  VNStageIntLLRInputS7xD(246)(1) <= CNStageIntLLROutputS7xD(69)(3);
  VNStageIntLLRInputS7xD(276)(1) <= CNStageIntLLROutputS7xD(69)(4);
  VNStageIntLLRInputS7xD(343)(1) <= CNStageIntLLROutputS7xD(69)(5);
  VNStageIntLLRInputS7xD(26)(1) <= CNStageIntLLROutputS7xD(70)(0);
  VNStageIntLLRInputS7xD(74)(1) <= CNStageIntLLROutputS7xD(70)(1);
  VNStageIntLLRInputS7xD(181)(1) <= CNStageIntLLROutputS7xD(70)(2);
  VNStageIntLLRInputS7xD(211)(1) <= CNStageIntLLROutputS7xD(70)(3);
  VNStageIntLLRInputS7xD(278)(1) <= CNStageIntLLROutputS7xD(70)(4);
  VNStageIntLLRInputS7xD(325)(1) <= CNStageIntLLROutputS7xD(70)(5);
  VNStageIntLLRInputS7xD(25)(1) <= CNStageIntLLROutputS7xD(71)(0);
  VNStageIntLLRInputS7xD(116)(0) <= CNStageIntLLROutputS7xD(71)(1);
  VNStageIntLLRInputS7xD(146)(1) <= CNStageIntLLROutputS7xD(71)(2);
  VNStageIntLLRInputS7xD(213)(1) <= CNStageIntLLROutputS7xD(71)(3);
  VNStageIntLLRInputS7xD(260)(1) <= CNStageIntLLROutputS7xD(71)(4);
  VNStageIntLLRInputS7xD(332)(1) <= CNStageIntLLROutputS7xD(71)(5);
  VNStageIntLLRInputS7xD(24)(1) <= CNStageIntLLROutputS7xD(72)(0);
  VNStageIntLLRInputS7xD(81)(1) <= CNStageIntLLROutputS7xD(72)(1);
  VNStageIntLLRInputS7xD(148)(1) <= CNStageIntLLROutputS7xD(72)(2);
  VNStageIntLLRInputS7xD(195)(0) <= CNStageIntLLROutputS7xD(72)(3);
  VNStageIntLLRInputS7xD(267)(1) <= CNStageIntLLROutputS7xD(72)(4);
  VNStageIntLLRInputS7xD(359)(1) <= CNStageIntLLROutputS7xD(72)(5);
  VNStageIntLLRInputS7xD(23)(1) <= CNStageIntLLROutputS7xD(73)(0);
  VNStageIntLLRInputS7xD(83)(1) <= CNStageIntLLROutputS7xD(73)(1);
  VNStageIntLLRInputS7xD(130)(1) <= CNStageIntLLROutputS7xD(73)(2);
  VNStageIntLLRInputS7xD(202)(1) <= CNStageIntLLROutputS7xD(73)(3);
  VNStageIntLLRInputS7xD(294)(1) <= CNStageIntLLROutputS7xD(73)(4);
  VNStageIntLLRInputS7xD(347)(1) <= CNStageIntLLROutputS7xD(73)(5);
  VNStageIntLLRInputS7xD(22)(1) <= CNStageIntLLROutputS7xD(74)(0);
  VNStageIntLLRInputS7xD(65)(1) <= CNStageIntLLROutputS7xD(74)(1);
  VNStageIntLLRInputS7xD(137)(1) <= CNStageIntLLROutputS7xD(74)(2);
  VNStageIntLLRInputS7xD(229)(1) <= CNStageIntLLROutputS7xD(74)(3);
  VNStageIntLLRInputS7xD(282)(1) <= CNStageIntLLROutputS7xD(74)(4);
  VNStageIntLLRInputS7xD(353)(1) <= CNStageIntLLROutputS7xD(74)(5);
  VNStageIntLLRInputS7xD(21)(1) <= CNStageIntLLROutputS7xD(75)(0);
  VNStageIntLLRInputS7xD(72)(1) <= CNStageIntLLROutputS7xD(75)(1);
  VNStageIntLLRInputS7xD(164)(1) <= CNStageIntLLROutputS7xD(75)(2);
  VNStageIntLLRInputS7xD(217)(1) <= CNStageIntLLROutputS7xD(75)(3);
  VNStageIntLLRInputS7xD(288)(1) <= CNStageIntLLROutputS7xD(75)(4);
  VNStageIntLLRInputS7xD(348)(1) <= CNStageIntLLROutputS7xD(75)(5);
  VNStageIntLLRInputS7xD(20)(1) <= CNStageIntLLROutputS7xD(76)(0);
  VNStageIntLLRInputS7xD(99)(1) <= CNStageIntLLROutputS7xD(76)(1);
  VNStageIntLLRInputS7xD(152)(1) <= CNStageIntLLROutputS7xD(76)(2);
  VNStageIntLLRInputS7xD(223)(1) <= CNStageIntLLROutputS7xD(76)(3);
  VNStageIntLLRInputS7xD(283)(1) <= CNStageIntLLROutputS7xD(76)(4);
  VNStageIntLLRInputS7xD(358)(1) <= CNStageIntLLROutputS7xD(76)(5);
  VNStageIntLLRInputS7xD(19)(1) <= CNStageIntLLROutputS7xD(77)(0);
  VNStageIntLLRInputS7xD(87)(1) <= CNStageIntLLROutputS7xD(77)(1);
  VNStageIntLLRInputS7xD(158)(1) <= CNStageIntLLROutputS7xD(77)(2);
  VNStageIntLLRInputS7xD(218)(1) <= CNStageIntLLROutputS7xD(77)(3);
  VNStageIntLLRInputS7xD(293)(1) <= CNStageIntLLROutputS7xD(77)(4);
  VNStageIntLLRInputS7xD(380)(0) <= CNStageIntLLROutputS7xD(77)(5);
  VNStageIntLLRInputS7xD(18)(1) <= CNStageIntLLROutputS7xD(78)(0);
  VNStageIntLLRInputS7xD(93)(1) <= CNStageIntLLROutputS7xD(78)(1);
  VNStageIntLLRInputS7xD(153)(1) <= CNStageIntLLROutputS7xD(78)(2);
  VNStageIntLLRInputS7xD(228)(1) <= CNStageIntLLROutputS7xD(78)(3);
  VNStageIntLLRInputS7xD(315)(0) <= CNStageIntLLROutputS7xD(78)(4);
  VNStageIntLLRInputS7xD(335)(1) <= CNStageIntLLROutputS7xD(78)(5);
  VNStageIntLLRInputS7xD(17)(1) <= CNStageIntLLROutputS7xD(79)(0);
  VNStageIntLLRInputS7xD(88)(1) <= CNStageIntLLROutputS7xD(79)(1);
  VNStageIntLLRInputS7xD(163)(1) <= CNStageIntLLROutputS7xD(79)(2);
  VNStageIntLLRInputS7xD(250)(0) <= CNStageIntLLROutputS7xD(79)(3);
  VNStageIntLLRInputS7xD(270)(1) <= CNStageIntLLROutputS7xD(79)(4);
  VNStageIntLLRInputS7xD(383)(1) <= CNStageIntLLROutputS7xD(79)(5);
  VNStageIntLLRInputS7xD(15)(1) <= CNStageIntLLROutputS7xD(80)(0);
  VNStageIntLLRInputS7xD(120)(1) <= CNStageIntLLROutputS7xD(80)(1);
  VNStageIntLLRInputS7xD(140)(1) <= CNStageIntLLROutputS7xD(80)(2);
  VNStageIntLLRInputS7xD(253)(0) <= CNStageIntLLROutputS7xD(80)(3);
  VNStageIntLLRInputS7xD(305)(1) <= CNStageIntLLROutputS7xD(80)(4);
  VNStageIntLLRInputS7xD(338)(1) <= CNStageIntLLROutputS7xD(80)(5);
  VNStageIntLLRInputS7xD(14)(1) <= CNStageIntLLROutputS7xD(81)(0);
  VNStageIntLLRInputS7xD(75)(1) <= CNStageIntLLROutputS7xD(81)(1);
  VNStageIntLLRInputS7xD(188)(0) <= CNStageIntLLROutputS7xD(81)(2);
  VNStageIntLLRInputS7xD(240)(1) <= CNStageIntLLROutputS7xD(81)(3);
  VNStageIntLLRInputS7xD(273)(1) <= CNStageIntLLROutputS7xD(81)(4);
  VNStageIntLLRInputS7xD(350)(1) <= CNStageIntLLROutputS7xD(81)(5);
  VNStageIntLLRInputS7xD(13)(0) <= CNStageIntLLROutputS7xD(82)(0);
  VNStageIntLLRInputS7xD(123)(0) <= CNStageIntLLROutputS7xD(82)(1);
  VNStageIntLLRInputS7xD(175)(1) <= CNStageIntLLROutputS7xD(82)(2);
  VNStageIntLLRInputS7xD(208)(1) <= CNStageIntLLROutputS7xD(82)(3);
  VNStageIntLLRInputS7xD(285)(1) <= CNStageIntLLROutputS7xD(82)(4);
  VNStageIntLLRInputS7xD(364)(1) <= CNStageIntLLROutputS7xD(82)(5);
  VNStageIntLLRInputS7xD(12)(1) <= CNStageIntLLROutputS7xD(83)(0);
  VNStageIntLLRInputS7xD(110)(1) <= CNStageIntLLROutputS7xD(83)(1);
  VNStageIntLLRInputS7xD(143)(1) <= CNStageIntLLROutputS7xD(83)(2);
  VNStageIntLLRInputS7xD(220)(1) <= CNStageIntLLROutputS7xD(83)(3);
  VNStageIntLLRInputS7xD(299)(0) <= CNStageIntLLROutputS7xD(83)(4);
  VNStageIntLLRInputS7xD(345)(1) <= CNStageIntLLROutputS7xD(83)(5);
  VNStageIntLLRInputS7xD(11)(1) <= CNStageIntLLROutputS7xD(84)(0);
  VNStageIntLLRInputS7xD(78)(1) <= CNStageIntLLROutputS7xD(84)(1);
  VNStageIntLLRInputS7xD(155)(1) <= CNStageIntLLROutputS7xD(84)(2);
  VNStageIntLLRInputS7xD(234)(1) <= CNStageIntLLROutputS7xD(84)(3);
  VNStageIntLLRInputS7xD(280)(1) <= CNStageIntLLROutputS7xD(84)(4);
  VNStageIntLLRInputS7xD(322)(1) <= CNStageIntLLROutputS7xD(84)(5);
  VNStageIntLLRInputS7xD(10)(1) <= CNStageIntLLROutputS7xD(85)(0);
  VNStageIntLLRInputS7xD(90)(1) <= CNStageIntLLROutputS7xD(85)(1);
  VNStageIntLLRInputS7xD(169)(1) <= CNStageIntLLROutputS7xD(85)(2);
  VNStageIntLLRInputS7xD(215)(1) <= CNStageIntLLROutputS7xD(85)(3);
  VNStageIntLLRInputS7xD(257)(1) <= CNStageIntLLROutputS7xD(85)(4);
  VNStageIntLLRInputS7xD(374)(1) <= CNStageIntLLROutputS7xD(85)(5);
  VNStageIntLLRInputS7xD(9)(1) <= CNStageIntLLROutputS7xD(86)(0);
  VNStageIntLLRInputS7xD(104)(1) <= CNStageIntLLROutputS7xD(86)(1);
  VNStageIntLLRInputS7xD(150)(1) <= CNStageIntLLROutputS7xD(86)(2);
  VNStageIntLLRInputS7xD(255)(1) <= CNStageIntLLROutputS7xD(86)(3);
  VNStageIntLLRInputS7xD(309)(1) <= CNStageIntLLROutputS7xD(86)(4);
  VNStageIntLLRInputS7xD(378)(0) <= CNStageIntLLROutputS7xD(86)(5);
  VNStageIntLLRInputS7xD(7)(1) <= CNStageIntLLROutputS7xD(87)(0);
  VNStageIntLLRInputS7xD(125)(0) <= CNStageIntLLROutputS7xD(87)(1);
  VNStageIntLLRInputS7xD(179)(1) <= CNStageIntLLROutputS7xD(87)(2);
  VNStageIntLLRInputS7xD(248)(1) <= CNStageIntLLROutputS7xD(87)(3);
  VNStageIntLLRInputS7xD(306)(1) <= CNStageIntLLROutputS7xD(87)(4);
  VNStageIntLLRInputS7xD(382)(0) <= CNStageIntLLROutputS7xD(87)(5);
  VNStageIntLLRInputS7xD(6)(1) <= CNStageIntLLROutputS7xD(88)(0);
  VNStageIntLLRInputS7xD(114)(1) <= CNStageIntLLROutputS7xD(88)(1);
  VNStageIntLLRInputS7xD(183)(1) <= CNStageIntLLROutputS7xD(88)(2);
  VNStageIntLLRInputS7xD(241)(1) <= CNStageIntLLROutputS7xD(88)(3);
  VNStageIntLLRInputS7xD(317)(0) <= CNStageIntLLROutputS7xD(88)(4);
  VNStageIntLLRInputS7xD(354)(1) <= CNStageIntLLROutputS7xD(88)(5);
  VNStageIntLLRInputS7xD(5)(1) <= CNStageIntLLROutputS7xD(89)(0);
  VNStageIntLLRInputS7xD(118)(1) <= CNStageIntLLROutputS7xD(89)(1);
  VNStageIntLLRInputS7xD(176)(1) <= CNStageIntLLROutputS7xD(89)(2);
  VNStageIntLLRInputS7xD(252)(0) <= CNStageIntLLROutputS7xD(89)(3);
  VNStageIntLLRInputS7xD(289)(1) <= CNStageIntLLROutputS7xD(89)(4);
  VNStageIntLLRInputS7xD(346)(1) <= CNStageIntLLROutputS7xD(89)(5);
  VNStageIntLLRInputS7xD(4)(1) <= CNStageIntLLROutputS7xD(90)(0);
  VNStageIntLLRInputS7xD(111)(1) <= CNStageIntLLROutputS7xD(90)(1);
  VNStageIntLLRInputS7xD(187)(0) <= CNStageIntLLROutputS7xD(90)(2);
  VNStageIntLLRInputS7xD(224)(1) <= CNStageIntLLROutputS7xD(90)(3);
  VNStageIntLLRInputS7xD(281)(1) <= CNStageIntLLROutputS7xD(90)(4);
  VNStageIntLLRInputS7xD(363)(0) <= CNStageIntLLROutputS7xD(90)(5);
  VNStageIntLLRInputS7xD(3)(0) <= CNStageIntLLROutputS7xD(91)(0);
  VNStageIntLLRInputS7xD(122)(0) <= CNStageIntLLROutputS7xD(91)(1);
  VNStageIntLLRInputS7xD(159)(1) <= CNStageIntLLROutputS7xD(91)(2);
  VNStageIntLLRInputS7xD(216)(1) <= CNStageIntLLROutputS7xD(91)(3);
  VNStageIntLLRInputS7xD(298)(1) <= CNStageIntLLROutputS7xD(91)(4);
  VNStageIntLLRInputS7xD(360)(1) <= CNStageIntLLROutputS7xD(91)(5);
  VNStageIntLLRInputS7xD(2)(1) <= CNStageIntLLROutputS7xD(92)(0);
  VNStageIntLLRInputS7xD(94)(1) <= CNStageIntLLROutputS7xD(92)(1);
  VNStageIntLLRInputS7xD(151)(1) <= CNStageIntLLROutputS7xD(92)(2);
  VNStageIntLLRInputS7xD(233)(1) <= CNStageIntLLROutputS7xD(92)(3);
  VNStageIntLLRInputS7xD(295)(1) <= CNStageIntLLROutputS7xD(92)(4);
  VNStageIntLLRInputS7xD(331)(1) <= CNStageIntLLROutputS7xD(92)(5);
  VNStageIntLLRInputS7xD(63)(1) <= CNStageIntLLROutputS7xD(93)(0);
  VNStageIntLLRInputS7xD(103)(1) <= CNStageIntLLROutputS7xD(93)(1);
  VNStageIntLLRInputS7xD(165)(1) <= CNStageIntLLROutputS7xD(93)(2);
  VNStageIntLLRInputS7xD(201)(1) <= CNStageIntLLROutputS7xD(93)(3);
  VNStageIntLLRInputS7xD(286)(1) <= CNStageIntLLROutputS7xD(93)(4);
  VNStageIntLLRInputS7xD(337)(1) <= CNStageIntLLROutputS7xD(93)(5);
  VNStageIntLLRInputS7xD(62)(0) <= CNStageIntLLROutputS7xD(94)(0);
  VNStageIntLLRInputS7xD(100)(1) <= CNStageIntLLROutputS7xD(94)(1);
  VNStageIntLLRInputS7xD(136)(1) <= CNStageIntLLROutputS7xD(94)(2);
  VNStageIntLLRInputS7xD(221)(1) <= CNStageIntLLROutputS7xD(94)(3);
  VNStageIntLLRInputS7xD(272)(1) <= CNStageIntLLROutputS7xD(94)(4);
  VNStageIntLLRInputS7xD(327)(1) <= CNStageIntLLROutputS7xD(94)(5);
  VNStageIntLLRInputS7xD(61)(0) <= CNStageIntLLROutputS7xD(95)(0);
  VNStageIntLLRInputS7xD(71)(1) <= CNStageIntLLROutputS7xD(95)(1);
  VNStageIntLLRInputS7xD(156)(1) <= CNStageIntLLROutputS7xD(95)(2);
  VNStageIntLLRInputS7xD(207)(1) <= CNStageIntLLROutputS7xD(95)(3);
  VNStageIntLLRInputS7xD(262)(1) <= CNStageIntLLROutputS7xD(95)(4);
  VNStageIntLLRInputS7xD(356)(1) <= CNStageIntLLROutputS7xD(95)(5);
  VNStageIntLLRInputS7xD(60)(0) <= CNStageIntLLROutputS7xD(96)(0);
  VNStageIntLLRInputS7xD(91)(1) <= CNStageIntLLROutputS7xD(96)(1);
  VNStageIntLLRInputS7xD(142)(1) <= CNStageIntLLROutputS7xD(96)(2);
  VNStageIntLLRInputS7xD(197)(1) <= CNStageIntLLROutputS7xD(96)(3);
  VNStageIntLLRInputS7xD(291)(1) <= CNStageIntLLROutputS7xD(96)(4);
  VNStageIntLLRInputS7xD(339)(1) <= CNStageIntLLROutputS7xD(96)(5);
  VNStageIntLLRInputS7xD(58)(0) <= CNStageIntLLROutputS7xD(97)(0);
  VNStageIntLLRInputS7xD(67)(0) <= CNStageIntLLROutputS7xD(97)(1);
  VNStageIntLLRInputS7xD(161)(1) <= CNStageIntLLROutputS7xD(97)(2);
  VNStageIntLLRInputS7xD(209)(1) <= CNStageIntLLROutputS7xD(97)(3);
  VNStageIntLLRInputS7xD(304)(1) <= CNStageIntLLROutputS7xD(97)(4);
  VNStageIntLLRInputS7xD(329)(1) <= CNStageIntLLROutputS7xD(97)(5);
  VNStageIntLLRInputS7xD(57)(0) <= CNStageIntLLROutputS7xD(98)(0);
  VNStageIntLLRInputS7xD(96)(1) <= CNStageIntLLROutputS7xD(98)(1);
  VNStageIntLLRInputS7xD(144)(1) <= CNStageIntLLROutputS7xD(98)(2);
  VNStageIntLLRInputS7xD(239)(1) <= CNStageIntLLROutputS7xD(98)(3);
  VNStageIntLLRInputS7xD(264)(1) <= CNStageIntLLROutputS7xD(98)(4);
  VNStageIntLLRInputS7xD(365)(1) <= CNStageIntLLROutputS7xD(98)(5);
  VNStageIntLLRInputS7xD(56)(1) <= CNStageIntLLROutputS7xD(99)(0);
  VNStageIntLLRInputS7xD(79)(1) <= CNStageIntLLROutputS7xD(99)(1);
  VNStageIntLLRInputS7xD(174)(1) <= CNStageIntLLROutputS7xD(99)(2);
  VNStageIntLLRInputS7xD(199)(1) <= CNStageIntLLROutputS7xD(99)(3);
  VNStageIntLLRInputS7xD(300)(1) <= CNStageIntLLROutputS7xD(99)(4);
  VNStageIntLLRInputS7xD(349)(1) <= CNStageIntLLROutputS7xD(99)(5);
  VNStageIntLLRInputS7xD(55)(1) <= CNStageIntLLROutputS7xD(100)(0);
  VNStageIntLLRInputS7xD(109)(1) <= CNStageIntLLROutputS7xD(100)(1);
  VNStageIntLLRInputS7xD(134)(1) <= CNStageIntLLROutputS7xD(100)(2);
  VNStageIntLLRInputS7xD(235)(0) <= CNStageIntLLROutputS7xD(100)(3);
  VNStageIntLLRInputS7xD(284)(1) <= CNStageIntLLROutputS7xD(100)(4);
  VNStageIntLLRInputS7xD(352)(1) <= CNStageIntLLROutputS7xD(100)(5);
  VNStageIntLLRInputS7xD(54)(1) <= CNStageIntLLROutputS7xD(101)(0);
  VNStageIntLLRInputS7xD(69)(1) <= CNStageIntLLROutputS7xD(101)(1);
  VNStageIntLLRInputS7xD(170)(1) <= CNStageIntLLROutputS7xD(101)(2);
  VNStageIntLLRInputS7xD(219)(1) <= CNStageIntLLROutputS7xD(101)(3);
  VNStageIntLLRInputS7xD(287)(1) <= CNStageIntLLROutputS7xD(101)(4);
  VNStageIntLLRInputS7xD(330)(1) <= CNStageIntLLROutputS7xD(101)(5);
  VNStageIntLLRInputS7xD(52)(0) <= CNStageIntLLROutputS7xD(102)(0);
  VNStageIntLLRInputS7xD(89)(1) <= CNStageIntLLROutputS7xD(102)(1);
  VNStageIntLLRInputS7xD(157)(1) <= CNStageIntLLROutputS7xD(102)(2);
  VNStageIntLLRInputS7xD(200)(1) <= CNStageIntLLROutputS7xD(102)(3);
  VNStageIntLLRInputS7xD(303)(1) <= CNStageIntLLROutputS7xD(102)(4);
  VNStageIntLLRInputS7xD(366)(1) <= CNStageIntLLROutputS7xD(102)(5);
  VNStageIntLLRInputS7xD(51)(1) <= CNStageIntLLROutputS7xD(103)(0);
  VNStageIntLLRInputS7xD(92)(1) <= CNStageIntLLROutputS7xD(103)(1);
  VNStageIntLLRInputS7xD(135)(1) <= CNStageIntLLROutputS7xD(103)(2);
  VNStageIntLLRInputS7xD(238)(1) <= CNStageIntLLROutputS7xD(103)(3);
  VNStageIntLLRInputS7xD(301)(1) <= CNStageIntLLROutputS7xD(103)(4);
  VNStageIntLLRInputS7xD(328)(1) <= CNStageIntLLROutputS7xD(103)(5);
  VNStageIntLLRInputS7xD(50)(1) <= CNStageIntLLROutputS7xD(104)(0);
  VNStageIntLLRInputS7xD(70)(1) <= CNStageIntLLROutputS7xD(104)(1);
  VNStageIntLLRInputS7xD(173)(1) <= CNStageIntLLROutputS7xD(104)(2);
  VNStageIntLLRInputS7xD(236)(1) <= CNStageIntLLROutputS7xD(104)(3);
  VNStageIntLLRInputS7xD(263)(1) <= CNStageIntLLROutputS7xD(104)(4);
  VNStageIntLLRInputS7xD(336)(1) <= CNStageIntLLROutputS7xD(104)(5);
  VNStageIntLLRInputS7xD(49)(1) <= CNStageIntLLROutputS7xD(105)(0);
  VNStageIntLLRInputS7xD(108)(1) <= CNStageIntLLROutputS7xD(105)(1);
  VNStageIntLLRInputS7xD(171)(0) <= CNStageIntLLROutputS7xD(105)(2);
  VNStageIntLLRInputS7xD(198)(1) <= CNStageIntLLROutputS7xD(105)(3);
  VNStageIntLLRInputS7xD(271)(1) <= CNStageIntLLROutputS7xD(105)(4);
  VNStageIntLLRInputS7xD(379)(0) <= CNStageIntLLROutputS7xD(105)(5);
  VNStageIntLLRInputS7xD(46)(1) <= CNStageIntLLROutputS7xD(106)(0);
  VNStageIntLLRInputS7xD(76)(1) <= CNStageIntLLROutputS7xD(106)(1);
  VNStageIntLLRInputS7xD(184)(1) <= CNStageIntLLROutputS7xD(106)(2);
  VNStageIntLLRInputS7xD(243)(1) <= CNStageIntLLROutputS7xD(106)(3);
  VNStageIntLLRInputS7xD(256)(1) <= CNStageIntLLROutputS7xD(106)(4);
  VNStageIntLLRInputS7xD(372)(0) <= CNStageIntLLROutputS7xD(106)(5);
  VNStageIntLLRInputS7xD(45)(1) <= CNStageIntLLROutputS7xD(107)(0);
  VNStageIntLLRInputS7xD(119)(1) <= CNStageIntLLROutputS7xD(107)(1);
  VNStageIntLLRInputS7xD(178)(1) <= CNStageIntLLROutputS7xD(107)(2);
  VNStageIntLLRInputS7xD(192)(1) <= CNStageIntLLROutputS7xD(107)(3);
  VNStageIntLLRInputS7xD(307)(1) <= CNStageIntLLROutputS7xD(107)(4);
  VNStageIntLLRInputS7xD(377)(0) <= CNStageIntLLROutputS7xD(107)(5);
  VNStageIntLLRInputS7xD(44)(1) <= CNStageIntLLROutputS7xD(108)(0);
  VNStageIntLLRInputS7xD(113)(1) <= CNStageIntLLROutputS7xD(108)(1);
  VNStageIntLLRInputS7xD(128)(1) <= CNStageIntLLROutputS7xD(108)(2);
  VNStageIntLLRInputS7xD(242)(1) <= CNStageIntLLROutputS7xD(108)(3);
  VNStageIntLLRInputS7xD(312)(1) <= CNStageIntLLROutputS7xD(108)(4);
  VNStageIntLLRInputS7xD(333)(0) <= CNStageIntLLROutputS7xD(108)(5);
  VNStageIntLLRInputS7xD(43)(0) <= CNStageIntLLROutputS7xD(109)(0);
  VNStageIntLLRInputS7xD(64)(1) <= CNStageIntLLROutputS7xD(109)(1);
  VNStageIntLLRInputS7xD(177)(1) <= CNStageIntLLROutputS7xD(109)(2);
  VNStageIntLLRInputS7xD(247)(1) <= CNStageIntLLROutputS7xD(109)(3);
  VNStageIntLLRInputS7xD(268)(1) <= CNStageIntLLROutputS7xD(109)(4);
  VNStageIntLLRInputS7xD(324)(1) <= CNStageIntLLROutputS7xD(109)(5);
  VNStageIntLLRInputS7xD(0)(1) <= CNStageIntLLROutputS7xD(110)(0);
  VNStageIntLLRInputS7xD(107)(0) <= CNStageIntLLROutputS7xD(110)(1);
  VNStageIntLLRInputS7xD(172)(1) <= CNStageIntLLROutputS7xD(110)(2);
  VNStageIntLLRInputS7xD(237)(1) <= CNStageIntLLROutputS7xD(110)(3);
  VNStageIntLLRInputS7xD(302)(1) <= CNStageIntLLROutputS7xD(110)(4);
  VNStageIntLLRInputS7xD(367)(1) <= CNStageIntLLROutputS7xD(110)(5);
  VNStageIntLLRInputS7xD(32)(2) <= CNStageIntLLROutputS7xD(111)(0);
  VNStageIntLLRInputS7xD(117)(2) <= CNStageIntLLROutputS7xD(111)(1);
  VNStageIntLLRInputS7xD(136)(2) <= CNStageIntLLROutputS7xD(111)(2);
  VNStageIntLLRInputS7xD(198)(2) <= CNStageIntLLROutputS7xD(111)(3);
  VNStageIntLLRInputS7xD(297)(2) <= CNStageIntLLROutputS7xD(111)(4);
  VNStageIntLLRInputS7xD(382)(1) <= CNStageIntLLROutputS7xD(111)(5);
  VNStageIntLLRInputS7xD(30)(2) <= CNStageIntLLROutputS7xD(112)(0);
  VNStageIntLLRInputS7xD(68)(1) <= CNStageIntLLROutputS7xD(112)(1);
  VNStageIntLLRInputS7xD(167)(2) <= CNStageIntLLROutputS7xD(112)(2);
  VNStageIntLLRInputS7xD(252)(1) <= CNStageIntLLROutputS7xD(112)(3);
  VNStageIntLLRInputS7xD(303)(2) <= CNStageIntLLROutputS7xD(112)(4);
  VNStageIntLLRInputS7xD(358)(2) <= CNStageIntLLROutputS7xD(112)(5);
  VNStageIntLLRInputS7xD(29)(2) <= CNStageIntLLROutputS7xD(113)(0);
  VNStageIntLLRInputS7xD(102)(2) <= CNStageIntLLROutputS7xD(113)(1);
  VNStageIntLLRInputS7xD(187)(1) <= CNStageIntLLROutputS7xD(113)(2);
  VNStageIntLLRInputS7xD(238)(2) <= CNStageIntLLROutputS7xD(113)(3);
  VNStageIntLLRInputS7xD(293)(2) <= CNStageIntLLROutputS7xD(113)(4);
  VNStageIntLLRInputS7xD(324)(2) <= CNStageIntLLROutputS7xD(113)(5);
  VNStageIntLLRInputS7xD(28)(2) <= CNStageIntLLROutputS7xD(114)(0);
  VNStageIntLLRInputS7xD(122)(1) <= CNStageIntLLROutputS7xD(114)(1);
  VNStageIntLLRInputS7xD(173)(2) <= CNStageIntLLROutputS7xD(114)(2);
  VNStageIntLLRInputS7xD(228)(2) <= CNStageIntLLROutputS7xD(114)(3);
  VNStageIntLLRInputS7xD(259)(1) <= CNStageIntLLROutputS7xD(114)(4);
  VNStageIntLLRInputS7xD(370)(1) <= CNStageIntLLROutputS7xD(114)(5);
  VNStageIntLLRInputS7xD(27)(2) <= CNStageIntLLROutputS7xD(115)(0);
  VNStageIntLLRInputS7xD(108)(2) <= CNStageIntLLROutputS7xD(115)(1);
  VNStageIntLLRInputS7xD(163)(2) <= CNStageIntLLROutputS7xD(115)(2);
  VNStageIntLLRInputS7xD(194)(2) <= CNStageIntLLROutputS7xD(115)(3);
  VNStageIntLLRInputS7xD(305)(2) <= CNStageIntLLROutputS7xD(115)(4);
  VNStageIntLLRInputS7xD(337)(2) <= CNStageIntLLROutputS7xD(115)(5);
  VNStageIntLLRInputS7xD(26)(2) <= CNStageIntLLROutputS7xD(116)(0);
  VNStageIntLLRInputS7xD(98)(1) <= CNStageIntLLROutputS7xD(116)(1);
  VNStageIntLLRInputS7xD(129)(2) <= CNStageIntLLROutputS7xD(116)(2);
  VNStageIntLLRInputS7xD(240)(2) <= CNStageIntLLROutputS7xD(116)(3);
  VNStageIntLLRInputS7xD(272)(2) <= CNStageIntLLROutputS7xD(116)(4);
  VNStageIntLLRInputS7xD(360)(2) <= CNStageIntLLROutputS7xD(116)(5);
  VNStageIntLLRInputS7xD(25)(2) <= CNStageIntLLROutputS7xD(117)(0);
  VNStageIntLLRInputS7xD(127)(2) <= CNStageIntLLROutputS7xD(117)(1);
  VNStageIntLLRInputS7xD(175)(2) <= CNStageIntLLROutputS7xD(117)(2);
  VNStageIntLLRInputS7xD(207)(2) <= CNStageIntLLROutputS7xD(117)(3);
  VNStageIntLLRInputS7xD(295)(2) <= CNStageIntLLROutputS7xD(117)(4);
  VNStageIntLLRInputS7xD(333)(1) <= CNStageIntLLROutputS7xD(117)(5);
  VNStageIntLLRInputS7xD(24)(2) <= CNStageIntLLROutputS7xD(118)(0);
  VNStageIntLLRInputS7xD(110)(2) <= CNStageIntLLROutputS7xD(118)(1);
  VNStageIntLLRInputS7xD(142)(2) <= CNStageIntLLROutputS7xD(118)(2);
  VNStageIntLLRInputS7xD(230)(1) <= CNStageIntLLROutputS7xD(118)(3);
  VNStageIntLLRInputS7xD(268)(2) <= CNStageIntLLROutputS7xD(118)(4);
  VNStageIntLLRInputS7xD(380)(1) <= CNStageIntLLROutputS7xD(118)(5);
  VNStageIntLLRInputS7xD(23)(2) <= CNStageIntLLROutputS7xD(119)(0);
  VNStageIntLLRInputS7xD(77)(0) <= CNStageIntLLROutputS7xD(119)(1);
  VNStageIntLLRInputS7xD(165)(2) <= CNStageIntLLROutputS7xD(119)(2);
  VNStageIntLLRInputS7xD(203)(2) <= CNStageIntLLROutputS7xD(119)(3);
  VNStageIntLLRInputS7xD(315)(1) <= CNStageIntLLROutputS7xD(119)(4);
  VNStageIntLLRInputS7xD(383)(2) <= CNStageIntLLROutputS7xD(119)(5);
  VNStageIntLLRInputS7xD(22)(2) <= CNStageIntLLROutputS7xD(120)(0);
  VNStageIntLLRInputS7xD(100)(2) <= CNStageIntLLROutputS7xD(120)(1);
  VNStageIntLLRInputS7xD(138)(2) <= CNStageIntLLROutputS7xD(120)(2);
  VNStageIntLLRInputS7xD(250)(1) <= CNStageIntLLROutputS7xD(120)(3);
  VNStageIntLLRInputS7xD(318)(0) <= CNStageIntLLROutputS7xD(120)(4);
  VNStageIntLLRInputS7xD(361)(2) <= CNStageIntLLROutputS7xD(120)(5);
  VNStageIntLLRInputS7xD(21)(2) <= CNStageIntLLROutputS7xD(121)(0);
  VNStageIntLLRInputS7xD(73)(2) <= CNStageIntLLROutputS7xD(121)(1);
  VNStageIntLLRInputS7xD(185)(0) <= CNStageIntLLROutputS7xD(121)(2);
  VNStageIntLLRInputS7xD(253)(1) <= CNStageIntLLROutputS7xD(121)(3);
  VNStageIntLLRInputS7xD(296)(2) <= CNStageIntLLROutputS7xD(121)(4);
  VNStageIntLLRInputS7xD(336)(2) <= CNStageIntLLROutputS7xD(121)(5);
  VNStageIntLLRInputS7xD(19)(2) <= CNStageIntLLROutputS7xD(122)(0);
  VNStageIntLLRInputS7xD(123)(1) <= CNStageIntLLROutputS7xD(122)(1);
  VNStageIntLLRInputS7xD(166)(2) <= CNStageIntLLROutputS7xD(122)(2);
  VNStageIntLLRInputS7xD(206)(1) <= CNStageIntLLROutputS7xD(122)(3);
  VNStageIntLLRInputS7xD(269)(1) <= CNStageIntLLROutputS7xD(122)(4);
  VNStageIntLLRInputS7xD(359)(2) <= CNStageIntLLROutputS7xD(122)(5);
  VNStageIntLLRInputS7xD(18)(2) <= CNStageIntLLROutputS7xD(123)(0);
  VNStageIntLLRInputS7xD(101)(2) <= CNStageIntLLROutputS7xD(123)(1);
  VNStageIntLLRInputS7xD(141)(0) <= CNStageIntLLROutputS7xD(123)(2);
  VNStageIntLLRInputS7xD(204)(2) <= CNStageIntLLROutputS7xD(123)(3);
  VNStageIntLLRInputS7xD(294)(2) <= CNStageIntLLROutputS7xD(123)(4);
  VNStageIntLLRInputS7xD(367)(2) <= CNStageIntLLROutputS7xD(123)(5);
  VNStageIntLLRInputS7xD(17)(2) <= CNStageIntLLROutputS7xD(124)(0);
  VNStageIntLLRInputS7xD(76)(2) <= CNStageIntLLROutputS7xD(124)(1);
  VNStageIntLLRInputS7xD(139)(2) <= CNStageIntLLROutputS7xD(124)(2);
  VNStageIntLLRInputS7xD(229)(2) <= CNStageIntLLROutputS7xD(124)(3);
  VNStageIntLLRInputS7xD(302)(2) <= CNStageIntLLROutputS7xD(124)(4);
  VNStageIntLLRInputS7xD(347)(2) <= CNStageIntLLROutputS7xD(124)(5);
  VNStageIntLLRInputS7xD(16)(1) <= CNStageIntLLROutputS7xD(125)(0);
  VNStageIntLLRInputS7xD(74)(2) <= CNStageIntLLROutputS7xD(125)(1);
  VNStageIntLLRInputS7xD(164)(2) <= CNStageIntLLROutputS7xD(125)(2);
  VNStageIntLLRInputS7xD(237)(2) <= CNStageIntLLROutputS7xD(125)(3);
  VNStageIntLLRInputS7xD(282)(2) <= CNStageIntLLROutputS7xD(125)(4);
  VNStageIntLLRInputS7xD(341)(2) <= CNStageIntLLROutputS7xD(125)(5);
  VNStageIntLLRInputS7xD(15)(2) <= CNStageIntLLROutputS7xD(126)(0);
  VNStageIntLLRInputS7xD(99)(2) <= CNStageIntLLROutputS7xD(126)(1);
  VNStageIntLLRInputS7xD(172)(2) <= CNStageIntLLROutputS7xD(126)(2);
  VNStageIntLLRInputS7xD(217)(2) <= CNStageIntLLROutputS7xD(126)(3);
  VNStageIntLLRInputS7xD(276)(2) <= CNStageIntLLROutputS7xD(126)(4);
  VNStageIntLLRInputS7xD(320)(1) <= CNStageIntLLROutputS7xD(126)(5);
  VNStageIntLLRInputS7xD(14)(2) <= CNStageIntLLROutputS7xD(127)(0);
  VNStageIntLLRInputS7xD(107)(1) <= CNStageIntLLROutputS7xD(127)(1);
  VNStageIntLLRInputS7xD(152)(2) <= CNStageIntLLROutputS7xD(127)(2);
  VNStageIntLLRInputS7xD(211)(2) <= CNStageIntLLROutputS7xD(127)(3);
  VNStageIntLLRInputS7xD(256)(2) <= CNStageIntLLROutputS7xD(127)(4);
  VNStageIntLLRInputS7xD(340)(2) <= CNStageIntLLROutputS7xD(127)(5);
  VNStageIntLLRInputS7xD(13)(1) <= CNStageIntLLROutputS7xD(128)(0);
  VNStageIntLLRInputS7xD(87)(2) <= CNStageIntLLROutputS7xD(128)(1);
  VNStageIntLLRInputS7xD(146)(2) <= CNStageIntLLROutputS7xD(128)(2);
  VNStageIntLLRInputS7xD(192)(2) <= CNStageIntLLROutputS7xD(128)(3);
  VNStageIntLLRInputS7xD(275)(2) <= CNStageIntLLROutputS7xD(128)(4);
  VNStageIntLLRInputS7xD(345)(2) <= CNStageIntLLROutputS7xD(128)(5);
  VNStageIntLLRInputS7xD(12)(2) <= CNStageIntLLROutputS7xD(129)(0);
  VNStageIntLLRInputS7xD(81)(2) <= CNStageIntLLROutputS7xD(129)(1);
  VNStageIntLLRInputS7xD(128)(2) <= CNStageIntLLROutputS7xD(129)(2);
  VNStageIntLLRInputS7xD(210)(2) <= CNStageIntLLROutputS7xD(129)(3);
  VNStageIntLLRInputS7xD(280)(2) <= CNStageIntLLROutputS7xD(129)(4);
  VNStageIntLLRInputS7xD(364)(2) <= CNStageIntLLROutputS7xD(129)(5);
  VNStageIntLLRInputS7xD(11)(2) <= CNStageIntLLROutputS7xD(130)(0);
  VNStageIntLLRInputS7xD(64)(2) <= CNStageIntLLROutputS7xD(130)(1);
  VNStageIntLLRInputS7xD(145)(2) <= CNStageIntLLROutputS7xD(130)(2);
  VNStageIntLLRInputS7xD(215)(2) <= CNStageIntLLROutputS7xD(130)(3);
  VNStageIntLLRInputS7xD(299)(1) <= CNStageIntLLROutputS7xD(130)(4);
  VNStageIntLLRInputS7xD(355)(2) <= CNStageIntLLROutputS7xD(130)(5);
  VNStageIntLLRInputS7xD(10)(2) <= CNStageIntLLROutputS7xD(131)(0);
  VNStageIntLLRInputS7xD(80)(2) <= CNStageIntLLROutputS7xD(131)(1);
  VNStageIntLLRInputS7xD(150)(2) <= CNStageIntLLROutputS7xD(131)(2);
  VNStageIntLLRInputS7xD(234)(2) <= CNStageIntLLROutputS7xD(131)(3);
  VNStageIntLLRInputS7xD(290)(2) <= CNStageIntLLROutputS7xD(131)(4);
  VNStageIntLLRInputS7xD(329)(2) <= CNStageIntLLROutputS7xD(131)(5);
  VNStageIntLLRInputS7xD(9)(2) <= CNStageIntLLROutputS7xD(132)(0);
  VNStageIntLLRInputS7xD(85)(1) <= CNStageIntLLROutputS7xD(132)(1);
  VNStageIntLLRInputS7xD(169)(2) <= CNStageIntLLROutputS7xD(132)(2);
  VNStageIntLLRInputS7xD(225)(2) <= CNStageIntLLROutputS7xD(132)(3);
  VNStageIntLLRInputS7xD(264)(2) <= CNStageIntLLROutputS7xD(132)(4);
  VNStageIntLLRInputS7xD(330)(2) <= CNStageIntLLROutputS7xD(132)(5);
  VNStageIntLLRInputS7xD(8)(1) <= CNStageIntLLROutputS7xD(133)(0);
  VNStageIntLLRInputS7xD(104)(2) <= CNStageIntLLROutputS7xD(133)(1);
  VNStageIntLLRInputS7xD(160)(2) <= CNStageIntLLROutputS7xD(133)(2);
  VNStageIntLLRInputS7xD(199)(2) <= CNStageIntLLROutputS7xD(133)(3);
  VNStageIntLLRInputS7xD(265)(1) <= CNStageIntLLROutputS7xD(133)(4);
  VNStageIntLLRInputS7xD(354)(2) <= CNStageIntLLROutputS7xD(133)(5);
  VNStageIntLLRInputS7xD(7)(2) <= CNStageIntLLROutputS7xD(134)(0);
  VNStageIntLLRInputS7xD(95)(2) <= CNStageIntLLROutputS7xD(134)(1);
  VNStageIntLLRInputS7xD(134)(2) <= CNStageIntLLROutputS7xD(134)(2);
  VNStageIntLLRInputS7xD(200)(2) <= CNStageIntLLROutputS7xD(134)(3);
  VNStageIntLLRInputS7xD(289)(2) <= CNStageIntLLROutputS7xD(134)(4);
  VNStageIntLLRInputS7xD(375)(2) <= CNStageIntLLROutputS7xD(134)(5);
  VNStageIntLLRInputS7xD(6)(2) <= CNStageIntLLROutputS7xD(135)(0);
  VNStageIntLLRInputS7xD(69)(2) <= CNStageIntLLROutputS7xD(135)(1);
  VNStageIntLLRInputS7xD(135)(2) <= CNStageIntLLROutputS7xD(135)(2);
  VNStageIntLLRInputS7xD(224)(2) <= CNStageIntLLROutputS7xD(135)(3);
  VNStageIntLLRInputS7xD(310)(2) <= CNStageIntLLROutputS7xD(135)(4);
  VNStageIntLLRInputS7xD(371)(1) <= CNStageIntLLROutputS7xD(135)(5);
  VNStageIntLLRInputS7xD(5)(2) <= CNStageIntLLROutputS7xD(136)(0);
  VNStageIntLLRInputS7xD(70)(2) <= CNStageIntLLROutputS7xD(136)(1);
  VNStageIntLLRInputS7xD(159)(2) <= CNStageIntLLROutputS7xD(136)(2);
  VNStageIntLLRInputS7xD(245)(2) <= CNStageIntLLROutputS7xD(136)(3);
  VNStageIntLLRInputS7xD(306)(2) <= CNStageIntLLROutputS7xD(136)(4);
  VNStageIntLLRInputS7xD(323)(1) <= CNStageIntLLROutputS7xD(136)(5);
  VNStageIntLLRInputS7xD(3)(1) <= CNStageIntLLROutputS7xD(137)(0);
  VNStageIntLLRInputS7xD(115)(2) <= CNStageIntLLROutputS7xD(137)(1);
  VNStageIntLLRInputS7xD(176)(2) <= CNStageIntLLROutputS7xD(137)(2);
  VNStageIntLLRInputS7xD(193)(2) <= CNStageIntLLROutputS7xD(137)(3);
  VNStageIntLLRInputS7xD(284)(2) <= CNStageIntLLROutputS7xD(137)(4);
  VNStageIntLLRInputS7xD(325)(2) <= CNStageIntLLROutputS7xD(137)(5);
  VNStageIntLLRInputS7xD(2)(2) <= CNStageIntLLROutputS7xD(138)(0);
  VNStageIntLLRInputS7xD(111)(2) <= CNStageIntLLROutputS7xD(138)(1);
  VNStageIntLLRInputS7xD(191)(2) <= CNStageIntLLROutputS7xD(138)(2);
  VNStageIntLLRInputS7xD(219)(2) <= CNStageIntLLROutputS7xD(138)(3);
  VNStageIntLLRInputS7xD(260)(2) <= CNStageIntLLROutputS7xD(138)(4);
  VNStageIntLLRInputS7xD(357)(2) <= CNStageIntLLROutputS7xD(138)(5);
  VNStageIntLLRInputS7xD(1)(1) <= CNStageIntLLROutputS7xD(139)(0);
  VNStageIntLLRInputS7xD(126)(1) <= CNStageIntLLROutputS7xD(139)(1);
  VNStageIntLLRInputS7xD(154)(1) <= CNStageIntLLROutputS7xD(139)(2);
  VNStageIntLLRInputS7xD(195)(1) <= CNStageIntLLROutputS7xD(139)(3);
  VNStageIntLLRInputS7xD(292)(2) <= CNStageIntLLROutputS7xD(139)(4);
  VNStageIntLLRInputS7xD(373)(1) <= CNStageIntLLROutputS7xD(139)(5);
  VNStageIntLLRInputS7xD(63)(2) <= CNStageIntLLROutputS7xD(140)(0);
  VNStageIntLLRInputS7xD(89)(2) <= CNStageIntLLROutputS7xD(140)(1);
  VNStageIntLLRInputS7xD(130)(2) <= CNStageIntLLROutputS7xD(140)(2);
  VNStageIntLLRInputS7xD(227)(2) <= CNStageIntLLROutputS7xD(140)(3);
  VNStageIntLLRInputS7xD(308)(0) <= CNStageIntLLROutputS7xD(140)(4);
  VNStageIntLLRInputS7xD(343)(2) <= CNStageIntLLROutputS7xD(140)(5);
  VNStageIntLLRInputS7xD(62)(1) <= CNStageIntLLROutputS7xD(141)(0);
  VNStageIntLLRInputS7xD(65)(2) <= CNStageIntLLROutputS7xD(141)(1);
  VNStageIntLLRInputS7xD(162)(2) <= CNStageIntLLROutputS7xD(141)(2);
  VNStageIntLLRInputS7xD(243)(2) <= CNStageIntLLROutputS7xD(141)(3);
  VNStageIntLLRInputS7xD(278)(2) <= CNStageIntLLROutputS7xD(141)(4);
  VNStageIntLLRInputS7xD(352)(2) <= CNStageIntLLROutputS7xD(141)(5);
  VNStageIntLLRInputS7xD(61)(1) <= CNStageIntLLROutputS7xD(142)(0);
  VNStageIntLLRInputS7xD(97)(2) <= CNStageIntLLROutputS7xD(142)(1);
  VNStageIntLLRInputS7xD(178)(2) <= CNStageIntLLROutputS7xD(142)(2);
  VNStageIntLLRInputS7xD(213)(2) <= CNStageIntLLROutputS7xD(142)(3);
  VNStageIntLLRInputS7xD(287)(2) <= CNStageIntLLROutputS7xD(142)(4);
  VNStageIntLLRInputS7xD(365)(2) <= CNStageIntLLROutputS7xD(142)(5);
  VNStageIntLLRInputS7xD(60)(1) <= CNStageIntLLROutputS7xD(143)(0);
  VNStageIntLLRInputS7xD(113)(2) <= CNStageIntLLROutputS7xD(143)(1);
  VNStageIntLLRInputS7xD(148)(2) <= CNStageIntLLROutputS7xD(143)(2);
  VNStageIntLLRInputS7xD(222)(1) <= CNStageIntLLROutputS7xD(143)(3);
  VNStageIntLLRInputS7xD(300)(2) <= CNStageIntLLROutputS7xD(143)(4);
  VNStageIntLLRInputS7xD(344)(2) <= CNStageIntLLROutputS7xD(143)(5);
  VNStageIntLLRInputS7xD(59)(0) <= CNStageIntLLROutputS7xD(144)(0);
  VNStageIntLLRInputS7xD(83)(2) <= CNStageIntLLROutputS7xD(144)(1);
  VNStageIntLLRInputS7xD(157)(2) <= CNStageIntLLROutputS7xD(144)(2);
  VNStageIntLLRInputS7xD(235)(1) <= CNStageIntLLROutputS7xD(144)(3);
  VNStageIntLLRInputS7xD(279)(2) <= CNStageIntLLROutputS7xD(144)(4);
  VNStageIntLLRInputS7xD(372)(1) <= CNStageIntLLROutputS7xD(144)(5);
  VNStageIntLLRInputS7xD(58)(1) <= CNStageIntLLROutputS7xD(145)(0);
  VNStageIntLLRInputS7xD(92)(2) <= CNStageIntLLROutputS7xD(145)(1);
  VNStageIntLLRInputS7xD(170)(2) <= CNStageIntLLROutputS7xD(145)(2);
  VNStageIntLLRInputS7xD(214)(2) <= CNStageIntLLROutputS7xD(145)(3);
  VNStageIntLLRInputS7xD(307)(2) <= CNStageIntLLROutputS7xD(145)(4);
  VNStageIntLLRInputS7xD(374)(2) <= CNStageIntLLROutputS7xD(145)(5);
  VNStageIntLLRInputS7xD(57)(1) <= CNStageIntLLROutputS7xD(146)(0);
  VNStageIntLLRInputS7xD(105)(1) <= CNStageIntLLROutputS7xD(146)(1);
  VNStageIntLLRInputS7xD(149)(2) <= CNStageIntLLROutputS7xD(146)(2);
  VNStageIntLLRInputS7xD(242)(2) <= CNStageIntLLROutputS7xD(146)(3);
  VNStageIntLLRInputS7xD(309)(2) <= CNStageIntLLROutputS7xD(146)(4);
  VNStageIntLLRInputS7xD(356)(2) <= CNStageIntLLROutputS7xD(146)(5);
  VNStageIntLLRInputS7xD(56)(2) <= CNStageIntLLROutputS7xD(147)(0);
  VNStageIntLLRInputS7xD(84)(2) <= CNStageIntLLROutputS7xD(147)(1);
  VNStageIntLLRInputS7xD(177)(2) <= CNStageIntLLROutputS7xD(147)(2);
  VNStageIntLLRInputS7xD(244)(0) <= CNStageIntLLROutputS7xD(147)(3);
  VNStageIntLLRInputS7xD(291)(2) <= CNStageIntLLROutputS7xD(147)(4);
  VNStageIntLLRInputS7xD(363)(1) <= CNStageIntLLROutputS7xD(147)(5);
  VNStageIntLLRInputS7xD(55)(2) <= CNStageIntLLROutputS7xD(148)(0);
  VNStageIntLLRInputS7xD(112)(2) <= CNStageIntLLROutputS7xD(148)(1);
  VNStageIntLLRInputS7xD(179)(2) <= CNStageIntLLROutputS7xD(148)(2);
  VNStageIntLLRInputS7xD(226)(1) <= CNStageIntLLROutputS7xD(148)(3);
  VNStageIntLLRInputS7xD(298)(2) <= CNStageIntLLROutputS7xD(148)(4);
  VNStageIntLLRInputS7xD(327)(2) <= CNStageIntLLROutputS7xD(148)(5);
  VNStageIntLLRInputS7xD(54)(2) <= CNStageIntLLROutputS7xD(149)(0);
  VNStageIntLLRInputS7xD(114)(2) <= CNStageIntLLROutputS7xD(149)(1);
  VNStageIntLLRInputS7xD(161)(2) <= CNStageIntLLROutputS7xD(149)(2);
  VNStageIntLLRInputS7xD(233)(2) <= CNStageIntLLROutputS7xD(149)(3);
  VNStageIntLLRInputS7xD(262)(2) <= CNStageIntLLROutputS7xD(149)(4);
  VNStageIntLLRInputS7xD(378)(1) <= CNStageIntLLROutputS7xD(149)(5);
  VNStageIntLLRInputS7xD(53)(1) <= CNStageIntLLROutputS7xD(150)(0);
  VNStageIntLLRInputS7xD(96)(2) <= CNStageIntLLROutputS7xD(150)(1);
  VNStageIntLLRInputS7xD(168)(1) <= CNStageIntLLROutputS7xD(150)(2);
  VNStageIntLLRInputS7xD(197)(2) <= CNStageIntLLROutputS7xD(150)(3);
  VNStageIntLLRInputS7xD(313)(0) <= CNStageIntLLROutputS7xD(150)(4);
  VNStageIntLLRInputS7xD(321)(2) <= CNStageIntLLROutputS7xD(150)(5);
  VNStageIntLLRInputS7xD(52)(1) <= CNStageIntLLROutputS7xD(151)(0);
  VNStageIntLLRInputS7xD(103)(2) <= CNStageIntLLROutputS7xD(151)(1);
  VNStageIntLLRInputS7xD(132)(1) <= CNStageIntLLROutputS7xD(151)(2);
  VNStageIntLLRInputS7xD(248)(2) <= CNStageIntLLROutputS7xD(151)(3);
  VNStageIntLLRInputS7xD(319)(2) <= CNStageIntLLROutputS7xD(151)(4);
  VNStageIntLLRInputS7xD(379)(1) <= CNStageIntLLROutputS7xD(151)(5);
  VNStageIntLLRInputS7xD(50)(2) <= CNStageIntLLROutputS7xD(152)(0);
  VNStageIntLLRInputS7xD(118)(2) <= CNStageIntLLROutputS7xD(152)(1);
  VNStageIntLLRInputS7xD(189)(1) <= CNStageIntLLROutputS7xD(152)(2);
  VNStageIntLLRInputS7xD(249)(0) <= CNStageIntLLROutputS7xD(152)(3);
  VNStageIntLLRInputS7xD(261)(2) <= CNStageIntLLROutputS7xD(152)(4);
  VNStageIntLLRInputS7xD(348)(2) <= CNStageIntLLROutputS7xD(152)(5);
  VNStageIntLLRInputS7xD(49)(2) <= CNStageIntLLROutputS7xD(153)(0);
  VNStageIntLLRInputS7xD(124)(1) <= CNStageIntLLROutputS7xD(153)(1);
  VNStageIntLLRInputS7xD(184)(2) <= CNStageIntLLROutputS7xD(153)(2);
  VNStageIntLLRInputS7xD(196)(2) <= CNStageIntLLROutputS7xD(153)(3);
  VNStageIntLLRInputS7xD(283)(2) <= CNStageIntLLROutputS7xD(153)(4);
  VNStageIntLLRInputS7xD(366)(2) <= CNStageIntLLROutputS7xD(153)(5);
  VNStageIntLLRInputS7xD(48)(1) <= CNStageIntLLROutputS7xD(154)(0);
  VNStageIntLLRInputS7xD(119)(2) <= CNStageIntLLROutputS7xD(154)(1);
  VNStageIntLLRInputS7xD(131)(1) <= CNStageIntLLROutputS7xD(154)(2);
  VNStageIntLLRInputS7xD(218)(2) <= CNStageIntLLROutputS7xD(154)(3);
  VNStageIntLLRInputS7xD(301)(2) <= CNStageIntLLROutputS7xD(154)(4);
  VNStageIntLLRInputS7xD(351)(1) <= CNStageIntLLROutputS7xD(154)(5);
  VNStageIntLLRInputS7xD(47)(1) <= CNStageIntLLROutputS7xD(155)(0);
  VNStageIntLLRInputS7xD(66)(2) <= CNStageIntLLROutputS7xD(155)(1);
  VNStageIntLLRInputS7xD(153)(2) <= CNStageIntLLROutputS7xD(155)(2);
  VNStageIntLLRInputS7xD(236)(2) <= CNStageIntLLROutputS7xD(155)(3);
  VNStageIntLLRInputS7xD(286)(2) <= CNStageIntLLROutputS7xD(155)(4);
  VNStageIntLLRInputS7xD(338)(2) <= CNStageIntLLROutputS7xD(155)(5);
  VNStageIntLLRInputS7xD(46)(2) <= CNStageIntLLROutputS7xD(156)(0);
  VNStageIntLLRInputS7xD(88)(2) <= CNStageIntLLROutputS7xD(156)(1);
  VNStageIntLLRInputS7xD(171)(1) <= CNStageIntLLROutputS7xD(156)(2);
  VNStageIntLLRInputS7xD(221)(2) <= CNStageIntLLROutputS7xD(156)(3);
  VNStageIntLLRInputS7xD(273)(2) <= CNStageIntLLROutputS7xD(156)(4);
  VNStageIntLLRInputS7xD(369)(1) <= CNStageIntLLROutputS7xD(156)(5);
  VNStageIntLLRInputS7xD(45)(2) <= CNStageIntLLROutputS7xD(157)(0);
  VNStageIntLLRInputS7xD(106)(1) <= CNStageIntLLROutputS7xD(157)(1);
  VNStageIntLLRInputS7xD(156)(2) <= CNStageIntLLROutputS7xD(157)(2);
  VNStageIntLLRInputS7xD(208)(2) <= CNStageIntLLROutputS7xD(157)(3);
  VNStageIntLLRInputS7xD(304)(2) <= CNStageIntLLROutputS7xD(157)(4);
  VNStageIntLLRInputS7xD(381)(1) <= CNStageIntLLROutputS7xD(157)(5);
  VNStageIntLLRInputS7xD(44)(2) <= CNStageIntLLROutputS7xD(158)(0);
  VNStageIntLLRInputS7xD(91)(2) <= CNStageIntLLROutputS7xD(158)(1);
  VNStageIntLLRInputS7xD(143)(2) <= CNStageIntLLROutputS7xD(158)(2);
  VNStageIntLLRInputS7xD(239)(2) <= CNStageIntLLROutputS7xD(158)(3);
  VNStageIntLLRInputS7xD(316)(1) <= CNStageIntLLROutputS7xD(158)(4);
  VNStageIntLLRInputS7xD(332)(2) <= CNStageIntLLROutputS7xD(158)(5);
  VNStageIntLLRInputS7xD(43)(1) <= CNStageIntLLROutputS7xD(159)(0);
  VNStageIntLLRInputS7xD(78)(2) <= CNStageIntLLROutputS7xD(159)(1);
  VNStageIntLLRInputS7xD(174)(2) <= CNStageIntLLROutputS7xD(159)(2);
  VNStageIntLLRInputS7xD(251)(1) <= CNStageIntLLROutputS7xD(159)(3);
  VNStageIntLLRInputS7xD(267)(2) <= CNStageIntLLROutputS7xD(159)(4);
  VNStageIntLLRInputS7xD(376)(2) <= CNStageIntLLROutputS7xD(159)(5);
  VNStageIntLLRInputS7xD(42)(2) <= CNStageIntLLROutputS7xD(160)(0);
  VNStageIntLLRInputS7xD(109)(2) <= CNStageIntLLROutputS7xD(160)(1);
  VNStageIntLLRInputS7xD(186)(1) <= CNStageIntLLROutputS7xD(160)(2);
  VNStageIntLLRInputS7xD(202)(2) <= CNStageIntLLROutputS7xD(160)(3);
  VNStageIntLLRInputS7xD(311)(2) <= CNStageIntLLROutputS7xD(160)(4);
  VNStageIntLLRInputS7xD(353)(2) <= CNStageIntLLROutputS7xD(160)(5);
  VNStageIntLLRInputS7xD(41)(2) <= CNStageIntLLROutputS7xD(161)(0);
  VNStageIntLLRInputS7xD(121)(1) <= CNStageIntLLROutputS7xD(161)(1);
  VNStageIntLLRInputS7xD(137)(2) <= CNStageIntLLROutputS7xD(161)(2);
  VNStageIntLLRInputS7xD(246)(2) <= CNStageIntLLROutputS7xD(161)(3);
  VNStageIntLLRInputS7xD(288)(2) <= CNStageIntLLROutputS7xD(161)(4);
  VNStageIntLLRInputS7xD(342)(2) <= CNStageIntLLROutputS7xD(161)(5);
  VNStageIntLLRInputS7xD(40)(2) <= CNStageIntLLROutputS7xD(162)(0);
  VNStageIntLLRInputS7xD(72)(2) <= CNStageIntLLROutputS7xD(162)(1);
  VNStageIntLLRInputS7xD(181)(2) <= CNStageIntLLROutputS7xD(162)(2);
  VNStageIntLLRInputS7xD(223)(2) <= CNStageIntLLROutputS7xD(162)(3);
  VNStageIntLLRInputS7xD(277)(2) <= CNStageIntLLROutputS7xD(162)(4);
  VNStageIntLLRInputS7xD(346)(2) <= CNStageIntLLROutputS7xD(162)(5);
  VNStageIntLLRInputS7xD(39)(2) <= CNStageIntLLROutputS7xD(163)(0);
  VNStageIntLLRInputS7xD(116)(1) <= CNStageIntLLROutputS7xD(163)(1);
  VNStageIntLLRInputS7xD(158)(2) <= CNStageIntLLROutputS7xD(163)(2);
  VNStageIntLLRInputS7xD(212)(2) <= CNStageIntLLROutputS7xD(163)(3);
  VNStageIntLLRInputS7xD(281)(2) <= CNStageIntLLROutputS7xD(163)(4);
  VNStageIntLLRInputS7xD(339)(2) <= CNStageIntLLROutputS7xD(163)(5);
  VNStageIntLLRInputS7xD(38)(2) <= CNStageIntLLROutputS7xD(164)(0);
  VNStageIntLLRInputS7xD(93)(2) <= CNStageIntLLROutputS7xD(164)(1);
  VNStageIntLLRInputS7xD(147)(2) <= CNStageIntLLROutputS7xD(164)(2);
  VNStageIntLLRInputS7xD(216)(2) <= CNStageIntLLROutputS7xD(164)(3);
  VNStageIntLLRInputS7xD(274)(1) <= CNStageIntLLROutputS7xD(164)(4);
  VNStageIntLLRInputS7xD(350)(2) <= CNStageIntLLROutputS7xD(164)(5);
  VNStageIntLLRInputS7xD(37)(2) <= CNStageIntLLROutputS7xD(165)(0);
  VNStageIntLLRInputS7xD(82)(2) <= CNStageIntLLROutputS7xD(165)(1);
  VNStageIntLLRInputS7xD(151)(2) <= CNStageIntLLROutputS7xD(165)(2);
  VNStageIntLLRInputS7xD(209)(2) <= CNStageIntLLROutputS7xD(165)(3);
  VNStageIntLLRInputS7xD(285)(2) <= CNStageIntLLROutputS7xD(165)(4);
  VNStageIntLLRInputS7xD(322)(2) <= CNStageIntLLROutputS7xD(165)(5);
  VNStageIntLLRInputS7xD(36)(2) <= CNStageIntLLROutputS7xD(166)(0);
  VNStageIntLLRInputS7xD(86)(1) <= CNStageIntLLROutputS7xD(166)(1);
  VNStageIntLLRInputS7xD(144)(2) <= CNStageIntLLROutputS7xD(166)(2);
  VNStageIntLLRInputS7xD(220)(2) <= CNStageIntLLROutputS7xD(166)(3);
  VNStageIntLLRInputS7xD(257)(2) <= CNStageIntLLROutputS7xD(166)(4);
  VNStageIntLLRInputS7xD(377)(1) <= CNStageIntLLROutputS7xD(166)(5);
  VNStageIntLLRInputS7xD(35)(2) <= CNStageIntLLROutputS7xD(167)(0);
  VNStageIntLLRInputS7xD(79)(2) <= CNStageIntLLROutputS7xD(167)(1);
  VNStageIntLLRInputS7xD(155)(2) <= CNStageIntLLROutputS7xD(167)(2);
  VNStageIntLLRInputS7xD(255)(2) <= CNStageIntLLROutputS7xD(167)(3);
  VNStageIntLLRInputS7xD(312)(2) <= CNStageIntLLROutputS7xD(167)(4);
  VNStageIntLLRInputS7xD(331)(2) <= CNStageIntLLROutputS7xD(167)(5);
  VNStageIntLLRInputS7xD(34)(2) <= CNStageIntLLROutputS7xD(168)(0);
  VNStageIntLLRInputS7xD(90)(2) <= CNStageIntLLROutputS7xD(168)(1);
  VNStageIntLLRInputS7xD(190)(0) <= CNStageIntLLROutputS7xD(168)(2);
  VNStageIntLLRInputS7xD(247)(2) <= CNStageIntLLROutputS7xD(168)(3);
  VNStageIntLLRInputS7xD(266)(1) <= CNStageIntLLROutputS7xD(168)(4);
  VNStageIntLLRInputS7xD(328)(2) <= CNStageIntLLROutputS7xD(168)(5);
  VNStageIntLLRInputS7xD(33)(2) <= CNStageIntLLROutputS7xD(169)(0);
  VNStageIntLLRInputS7xD(125)(1) <= CNStageIntLLROutputS7xD(169)(1);
  VNStageIntLLRInputS7xD(182)(2) <= CNStageIntLLROutputS7xD(169)(2);
  VNStageIntLLRInputS7xD(201)(2) <= CNStageIntLLROutputS7xD(169)(3);
  VNStageIntLLRInputS7xD(263)(2) <= CNStageIntLLROutputS7xD(169)(4);
  VNStageIntLLRInputS7xD(362)(2) <= CNStageIntLLROutputS7xD(169)(5);
  VNStageIntLLRInputS7xD(0)(2) <= CNStageIntLLROutputS7xD(170)(0);
  VNStageIntLLRInputS7xD(75)(2) <= CNStageIntLLROutputS7xD(170)(1);
  VNStageIntLLRInputS7xD(140)(2) <= CNStageIntLLROutputS7xD(170)(2);
  VNStageIntLLRInputS7xD(205)(0) <= CNStageIntLLROutputS7xD(170)(3);
  VNStageIntLLRInputS7xD(270)(2) <= CNStageIntLLROutputS7xD(170)(4);
  VNStageIntLLRInputS7xD(335)(2) <= CNStageIntLLROutputS7xD(170)(5);
  VNStageIntLLRInputS7xD(62)(2) <= CNStageIntLLROutputS7xD(171)(0);
  VNStageIntLLRInputS7xD(109)(3) <= CNStageIntLLROutputS7xD(171)(1);
  VNStageIntLLRInputS7xD(161)(3) <= CNStageIntLLROutputS7xD(171)(2);
  VNStageIntLLRInputS7xD(194)(3) <= CNStageIntLLROutputS7xD(171)(3);
  VNStageIntLLRInputS7xD(271)(2) <= CNStageIntLLROutputS7xD(171)(4);
  VNStageIntLLRInputS7xD(350)(3) <= CNStageIntLLROutputS7xD(171)(5);
  VNStageIntLLRInputS7xD(61)(2) <= CNStageIntLLROutputS7xD(172)(0);
  VNStageIntLLRInputS7xD(96)(3) <= CNStageIntLLROutputS7xD(172)(1);
  VNStageIntLLRInputS7xD(129)(3) <= CNStageIntLLROutputS7xD(172)(2);
  VNStageIntLLRInputS7xD(206)(2) <= CNStageIntLLROutputS7xD(172)(3);
  VNStageIntLLRInputS7xD(285)(3) <= CNStageIntLLROutputS7xD(172)(4);
  VNStageIntLLRInputS7xD(331)(3) <= CNStageIntLLROutputS7xD(172)(5);
  VNStageIntLLRInputS7xD(60)(2) <= CNStageIntLLROutputS7xD(173)(0);
  VNStageIntLLRInputS7xD(127)(3) <= CNStageIntLLROutputS7xD(173)(1);
  VNStageIntLLRInputS7xD(141)(1) <= CNStageIntLLROutputS7xD(173)(2);
  VNStageIntLLRInputS7xD(220)(3) <= CNStageIntLLROutputS7xD(173)(3);
  VNStageIntLLRInputS7xD(266)(2) <= CNStageIntLLROutputS7xD(173)(4);
  VNStageIntLLRInputS7xD(371)(2) <= CNStageIntLLROutputS7xD(173)(5);
  VNStageIntLLRInputS7xD(59)(1) <= CNStageIntLLROutputS7xD(174)(0);
  VNStageIntLLRInputS7xD(76)(3) <= CNStageIntLLROutputS7xD(174)(1);
  VNStageIntLLRInputS7xD(155)(3) <= CNStageIntLLROutputS7xD(174)(2);
  VNStageIntLLRInputS7xD(201)(3) <= CNStageIntLLROutputS7xD(174)(3);
  VNStageIntLLRInputS7xD(306)(3) <= CNStageIntLLROutputS7xD(174)(4);
  VNStageIntLLRInputS7xD(360)(3) <= CNStageIntLLROutputS7xD(174)(5);
  VNStageIntLLRInputS7xD(58)(2) <= CNStageIntLLROutputS7xD(175)(0);
  VNStageIntLLRInputS7xD(90)(3) <= CNStageIntLLROutputS7xD(175)(1);
  VNStageIntLLRInputS7xD(136)(3) <= CNStageIntLLROutputS7xD(175)(2);
  VNStageIntLLRInputS7xD(241)(2) <= CNStageIntLLROutputS7xD(175)(3);
  VNStageIntLLRInputS7xD(295)(3) <= CNStageIntLLROutputS7xD(175)(4);
  VNStageIntLLRInputS7xD(364)(3) <= CNStageIntLLROutputS7xD(175)(5);
  VNStageIntLLRInputS7xD(57)(2) <= CNStageIntLLROutputS7xD(176)(0);
  VNStageIntLLRInputS7xD(71)(2) <= CNStageIntLLROutputS7xD(176)(1);
  VNStageIntLLRInputS7xD(176)(3) <= CNStageIntLLROutputS7xD(176)(2);
  VNStageIntLLRInputS7xD(230)(2) <= CNStageIntLLROutputS7xD(176)(3);
  VNStageIntLLRInputS7xD(299)(2) <= CNStageIntLLROutputS7xD(176)(4);
  VNStageIntLLRInputS7xD(357)(3) <= CNStageIntLLROutputS7xD(176)(5);
  VNStageIntLLRInputS7xD(56)(3) <= CNStageIntLLROutputS7xD(177)(0);
  VNStageIntLLRInputS7xD(111)(3) <= CNStageIntLLROutputS7xD(177)(1);
  VNStageIntLLRInputS7xD(165)(3) <= CNStageIntLLROutputS7xD(177)(2);
  VNStageIntLLRInputS7xD(234)(3) <= CNStageIntLLROutputS7xD(177)(3);
  VNStageIntLLRInputS7xD(292)(3) <= CNStageIntLLROutputS7xD(177)(4);
  VNStageIntLLRInputS7xD(368)(1) <= CNStageIntLLROutputS7xD(177)(5);
  VNStageIntLLRInputS7xD(55)(3) <= CNStageIntLLROutputS7xD(178)(0);
  VNStageIntLLRInputS7xD(100)(3) <= CNStageIntLLROutputS7xD(178)(1);
  VNStageIntLLRInputS7xD(169)(3) <= CNStageIntLLROutputS7xD(178)(2);
  VNStageIntLLRInputS7xD(227)(3) <= CNStageIntLLROutputS7xD(178)(3);
  VNStageIntLLRInputS7xD(303)(3) <= CNStageIntLLROutputS7xD(178)(4);
  VNStageIntLLRInputS7xD(340)(3) <= CNStageIntLLROutputS7xD(178)(5);
  VNStageIntLLRInputS7xD(54)(3) <= CNStageIntLLROutputS7xD(179)(0);
  VNStageIntLLRInputS7xD(104)(3) <= CNStageIntLLROutputS7xD(179)(1);
  VNStageIntLLRInputS7xD(162)(3) <= CNStageIntLLROutputS7xD(179)(2);
  VNStageIntLLRInputS7xD(238)(3) <= CNStageIntLLROutputS7xD(179)(3);
  VNStageIntLLRInputS7xD(275)(3) <= CNStageIntLLROutputS7xD(179)(4);
  VNStageIntLLRInputS7xD(332)(3) <= CNStageIntLLROutputS7xD(179)(5);
  VNStageIntLLRInputS7xD(53)(2) <= CNStageIntLLROutputS7xD(180)(0);
  VNStageIntLLRInputS7xD(97)(3) <= CNStageIntLLROutputS7xD(180)(1);
  VNStageIntLLRInputS7xD(173)(3) <= CNStageIntLLROutputS7xD(180)(2);
  VNStageIntLLRInputS7xD(210)(3) <= CNStageIntLLROutputS7xD(180)(3);
  VNStageIntLLRInputS7xD(267)(3) <= CNStageIntLLROutputS7xD(180)(4);
  VNStageIntLLRInputS7xD(349)(2) <= CNStageIntLLROutputS7xD(180)(5);
  VNStageIntLLRInputS7xD(52)(2) <= CNStageIntLLROutputS7xD(181)(0);
  VNStageIntLLRInputS7xD(108)(3) <= CNStageIntLLROutputS7xD(181)(1);
  VNStageIntLLRInputS7xD(145)(3) <= CNStageIntLLROutputS7xD(181)(2);
  VNStageIntLLRInputS7xD(202)(3) <= CNStageIntLLROutputS7xD(181)(3);
  VNStageIntLLRInputS7xD(284)(3) <= CNStageIntLLROutputS7xD(181)(4);
  VNStageIntLLRInputS7xD(346)(3) <= CNStageIntLLROutputS7xD(181)(5);
  VNStageIntLLRInputS7xD(51)(2) <= CNStageIntLLROutputS7xD(182)(0);
  VNStageIntLLRInputS7xD(80)(3) <= CNStageIntLLROutputS7xD(182)(1);
  VNStageIntLLRInputS7xD(137)(3) <= CNStageIntLLROutputS7xD(182)(2);
  VNStageIntLLRInputS7xD(219)(3) <= CNStageIntLLROutputS7xD(182)(3);
  VNStageIntLLRInputS7xD(281)(3) <= CNStageIntLLROutputS7xD(182)(4);
  VNStageIntLLRInputS7xD(380)(2) <= CNStageIntLLROutputS7xD(182)(5);
  VNStageIntLLRInputS7xD(50)(3) <= CNStageIntLLROutputS7xD(183)(0);
  VNStageIntLLRInputS7xD(72)(3) <= CNStageIntLLROutputS7xD(183)(1);
  VNStageIntLLRInputS7xD(154)(2) <= CNStageIntLLROutputS7xD(183)(2);
  VNStageIntLLRInputS7xD(216)(3) <= CNStageIntLLROutputS7xD(183)(3);
  VNStageIntLLRInputS7xD(315)(2) <= CNStageIntLLROutputS7xD(183)(4);
  VNStageIntLLRInputS7xD(337)(3) <= CNStageIntLLROutputS7xD(183)(5);
  VNStageIntLLRInputS7xD(49)(3) <= CNStageIntLLROutputS7xD(184)(0);
  VNStageIntLLRInputS7xD(89)(3) <= CNStageIntLLROutputS7xD(184)(1);
  VNStageIntLLRInputS7xD(151)(3) <= CNStageIntLLROutputS7xD(184)(2);
  VNStageIntLLRInputS7xD(250)(2) <= CNStageIntLLROutputS7xD(184)(3);
  VNStageIntLLRInputS7xD(272)(3) <= CNStageIntLLROutputS7xD(184)(4);
  VNStageIntLLRInputS7xD(323)(2) <= CNStageIntLLROutputS7xD(184)(5);
  VNStageIntLLRInputS7xD(46)(3) <= CNStageIntLLROutputS7xD(185)(0);
  VNStageIntLLRInputS7xD(77)(1) <= CNStageIntLLROutputS7xD(185)(1);
  VNStageIntLLRInputS7xD(191)(3) <= CNStageIntLLROutputS7xD(185)(2);
  VNStageIntLLRInputS7xD(246)(3) <= CNStageIntLLROutputS7xD(185)(3);
  VNStageIntLLRInputS7xD(277)(3) <= CNStageIntLLROutputS7xD(185)(4);
  VNStageIntLLRInputS7xD(325)(3) <= CNStageIntLLROutputS7xD(185)(5);
  VNStageIntLLRInputS7xD(45)(3) <= CNStageIntLLROutputS7xD(186)(0);
  VNStageIntLLRInputS7xD(126)(2) <= CNStageIntLLROutputS7xD(186)(1);
  VNStageIntLLRInputS7xD(181)(3) <= CNStageIntLLROutputS7xD(186)(2);
  VNStageIntLLRInputS7xD(212)(3) <= CNStageIntLLROutputS7xD(186)(3);
  VNStageIntLLRInputS7xD(260)(3) <= CNStageIntLLROutputS7xD(186)(4);
  VNStageIntLLRInputS7xD(355)(3) <= CNStageIntLLROutputS7xD(186)(5);
  VNStageIntLLRInputS7xD(44)(3) <= CNStageIntLLROutputS7xD(187)(0);
  VNStageIntLLRInputS7xD(116)(2) <= CNStageIntLLROutputS7xD(187)(1);
  VNStageIntLLRInputS7xD(147)(3) <= CNStageIntLLROutputS7xD(187)(2);
  VNStageIntLLRInputS7xD(195)(2) <= CNStageIntLLROutputS7xD(187)(3);
  VNStageIntLLRInputS7xD(290)(3) <= CNStageIntLLROutputS7xD(187)(4);
  VNStageIntLLRInputS7xD(378)(2) <= CNStageIntLLROutputS7xD(187)(5);
  VNStageIntLLRInputS7xD(43)(2) <= CNStageIntLLROutputS7xD(188)(0);
  VNStageIntLLRInputS7xD(82)(3) <= CNStageIntLLROutputS7xD(188)(1);
  VNStageIntLLRInputS7xD(130)(3) <= CNStageIntLLROutputS7xD(188)(2);
  VNStageIntLLRInputS7xD(225)(3) <= CNStageIntLLROutputS7xD(188)(3);
  VNStageIntLLRInputS7xD(313)(1) <= CNStageIntLLROutputS7xD(188)(4);
  VNStageIntLLRInputS7xD(351)(2) <= CNStageIntLLROutputS7xD(188)(5);
  VNStageIntLLRInputS7xD(42)(3) <= CNStageIntLLROutputS7xD(189)(0);
  VNStageIntLLRInputS7xD(65)(3) <= CNStageIntLLROutputS7xD(189)(1);
  VNStageIntLLRInputS7xD(160)(3) <= CNStageIntLLROutputS7xD(189)(2);
  VNStageIntLLRInputS7xD(248)(3) <= CNStageIntLLROutputS7xD(189)(3);
  VNStageIntLLRInputS7xD(286)(3) <= CNStageIntLLROutputS7xD(189)(4);
  VNStageIntLLRInputS7xD(335)(3) <= CNStageIntLLROutputS7xD(189)(5);
  VNStageIntLLRInputS7xD(41)(3) <= CNStageIntLLROutputS7xD(190)(0);
  VNStageIntLLRInputS7xD(95)(3) <= CNStageIntLLROutputS7xD(190)(1);
  VNStageIntLLRInputS7xD(183)(2) <= CNStageIntLLROutputS7xD(190)(2);
  VNStageIntLLRInputS7xD(221)(3) <= CNStageIntLLROutputS7xD(190)(3);
  VNStageIntLLRInputS7xD(270)(3) <= CNStageIntLLROutputS7xD(190)(4);
  VNStageIntLLRInputS7xD(338)(3) <= CNStageIntLLROutputS7xD(190)(5);
  VNStageIntLLRInputS7xD(39)(3) <= CNStageIntLLROutputS7xD(191)(0);
  VNStageIntLLRInputS7xD(91)(3) <= CNStageIntLLROutputS7xD(191)(1);
  VNStageIntLLRInputS7xD(140)(3) <= CNStageIntLLROutputS7xD(191)(2);
  VNStageIntLLRInputS7xD(208)(3) <= CNStageIntLLROutputS7xD(191)(3);
  VNStageIntLLRInputS7xD(314)(0) <= CNStageIntLLROutputS7xD(191)(4);
  VNStageIntLLRInputS7xD(354)(3) <= CNStageIntLLROutputS7xD(191)(5);
  VNStageIntLLRInputS7xD(38)(3) <= CNStageIntLLROutputS7xD(192)(0);
  VNStageIntLLRInputS7xD(75)(3) <= CNStageIntLLROutputS7xD(192)(1);
  VNStageIntLLRInputS7xD(143)(3) <= CNStageIntLLROutputS7xD(192)(2);
  VNStageIntLLRInputS7xD(249)(1) <= CNStageIntLLROutputS7xD(192)(3);
  VNStageIntLLRInputS7xD(289)(3) <= CNStageIntLLROutputS7xD(192)(4);
  VNStageIntLLRInputS7xD(352)(3) <= CNStageIntLLROutputS7xD(192)(5);
  VNStageIntLLRInputS7xD(37)(3) <= CNStageIntLLROutputS7xD(193)(0);
  VNStageIntLLRInputS7xD(78)(3) <= CNStageIntLLROutputS7xD(193)(1);
  VNStageIntLLRInputS7xD(184)(3) <= CNStageIntLLROutputS7xD(193)(2);
  VNStageIntLLRInputS7xD(224)(3) <= CNStageIntLLROutputS7xD(193)(3);
  VNStageIntLLRInputS7xD(287)(3) <= CNStageIntLLROutputS7xD(193)(4);
  VNStageIntLLRInputS7xD(377)(2) <= CNStageIntLLROutputS7xD(193)(5);
  VNStageIntLLRInputS7xD(35)(3) <= CNStageIntLLROutputS7xD(194)(0);
  VNStageIntLLRInputS7xD(94)(2) <= CNStageIntLLROutputS7xD(194)(1);
  VNStageIntLLRInputS7xD(157)(3) <= CNStageIntLLROutputS7xD(194)(2);
  VNStageIntLLRInputS7xD(247)(3) <= CNStageIntLLROutputS7xD(194)(3);
  VNStageIntLLRInputS7xD(257)(3) <= CNStageIntLLROutputS7xD(194)(4);
  VNStageIntLLRInputS7xD(365)(3) <= CNStageIntLLROutputS7xD(194)(5);
  VNStageIntLLRInputS7xD(34)(3) <= CNStageIntLLROutputS7xD(195)(0);
  VNStageIntLLRInputS7xD(92)(3) <= CNStageIntLLROutputS7xD(195)(1);
  VNStageIntLLRInputS7xD(182)(3) <= CNStageIntLLROutputS7xD(195)(2);
  VNStageIntLLRInputS7xD(255)(3) <= CNStageIntLLROutputS7xD(195)(3);
  VNStageIntLLRInputS7xD(300)(3) <= CNStageIntLLROutputS7xD(195)(4);
  VNStageIntLLRInputS7xD(359)(3) <= CNStageIntLLROutputS7xD(195)(5);
  VNStageIntLLRInputS7xD(33)(3) <= CNStageIntLLROutputS7xD(196)(0);
  VNStageIntLLRInputS7xD(117)(3) <= CNStageIntLLROutputS7xD(196)(1);
  VNStageIntLLRInputS7xD(190)(1) <= CNStageIntLLROutputS7xD(196)(2);
  VNStageIntLLRInputS7xD(235)(2) <= CNStageIntLLROutputS7xD(196)(3);
  VNStageIntLLRInputS7xD(294)(3) <= CNStageIntLLROutputS7xD(196)(4);
  VNStageIntLLRInputS7xD(320)(2) <= CNStageIntLLROutputS7xD(196)(5);
  VNStageIntLLRInputS7xD(31)(2) <= CNStageIntLLROutputS7xD(197)(0);
  VNStageIntLLRInputS7xD(105)(2) <= CNStageIntLLROutputS7xD(197)(1);
  VNStageIntLLRInputS7xD(164)(3) <= CNStageIntLLROutputS7xD(197)(2);
  VNStageIntLLRInputS7xD(192)(3) <= CNStageIntLLROutputS7xD(197)(3);
  VNStageIntLLRInputS7xD(293)(3) <= CNStageIntLLROutputS7xD(197)(4);
  VNStageIntLLRInputS7xD(363)(2) <= CNStageIntLLROutputS7xD(197)(5);
  VNStageIntLLRInputS7xD(30)(3) <= CNStageIntLLROutputS7xD(198)(0);
  VNStageIntLLRInputS7xD(99)(3) <= CNStageIntLLROutputS7xD(198)(1);
  VNStageIntLLRInputS7xD(128)(3) <= CNStageIntLLROutputS7xD(198)(2);
  VNStageIntLLRInputS7xD(228)(3) <= CNStageIntLLROutputS7xD(198)(3);
  VNStageIntLLRInputS7xD(298)(3) <= CNStageIntLLROutputS7xD(198)(4);
  VNStageIntLLRInputS7xD(382)(2) <= CNStageIntLLROutputS7xD(198)(5);
  VNStageIntLLRInputS7xD(28)(3) <= CNStageIntLLROutputS7xD(199)(0);
  VNStageIntLLRInputS7xD(98)(2) <= CNStageIntLLROutputS7xD(199)(1);
  VNStageIntLLRInputS7xD(168)(2) <= CNStageIntLLROutputS7xD(199)(2);
  VNStageIntLLRInputS7xD(252)(2) <= CNStageIntLLROutputS7xD(199)(3);
  VNStageIntLLRInputS7xD(308)(1) <= CNStageIntLLROutputS7xD(199)(4);
  VNStageIntLLRInputS7xD(347)(3) <= CNStageIntLLROutputS7xD(199)(5);
  VNStageIntLLRInputS7xD(27)(3) <= CNStageIntLLROutputS7xD(200)(0);
  VNStageIntLLRInputS7xD(103)(3) <= CNStageIntLLROutputS7xD(200)(1);
  VNStageIntLLRInputS7xD(187)(2) <= CNStageIntLLROutputS7xD(200)(2);
  VNStageIntLLRInputS7xD(243)(3) <= CNStageIntLLROutputS7xD(200)(3);
  VNStageIntLLRInputS7xD(282)(3) <= CNStageIntLLROutputS7xD(200)(4);
  VNStageIntLLRInputS7xD(348)(3) <= CNStageIntLLROutputS7xD(200)(5);
  VNStageIntLLRInputS7xD(26)(3) <= CNStageIntLLROutputS7xD(201)(0);
  VNStageIntLLRInputS7xD(122)(2) <= CNStageIntLLROutputS7xD(201)(1);
  VNStageIntLLRInputS7xD(178)(3) <= CNStageIntLLROutputS7xD(201)(2);
  VNStageIntLLRInputS7xD(217)(3) <= CNStageIntLLROutputS7xD(201)(3);
  VNStageIntLLRInputS7xD(283)(3) <= CNStageIntLLROutputS7xD(201)(4);
  VNStageIntLLRInputS7xD(372)(2) <= CNStageIntLLROutputS7xD(201)(5);
  VNStageIntLLRInputS7xD(25)(3) <= CNStageIntLLROutputS7xD(202)(0);
  VNStageIntLLRInputS7xD(113)(3) <= CNStageIntLLROutputS7xD(202)(1);
  VNStageIntLLRInputS7xD(152)(3) <= CNStageIntLLROutputS7xD(202)(2);
  VNStageIntLLRInputS7xD(218)(3) <= CNStageIntLLROutputS7xD(202)(3);
  VNStageIntLLRInputS7xD(307)(3) <= CNStageIntLLROutputS7xD(202)(4);
  VNStageIntLLRInputS7xD(330)(3) <= CNStageIntLLROutputS7xD(202)(5);
  VNStageIntLLRInputS7xD(24)(3) <= CNStageIntLLROutputS7xD(203)(0);
  VNStageIntLLRInputS7xD(87)(3) <= CNStageIntLLROutputS7xD(203)(1);
  VNStageIntLLRInputS7xD(153)(3) <= CNStageIntLLROutputS7xD(203)(2);
  VNStageIntLLRInputS7xD(242)(3) <= CNStageIntLLROutputS7xD(203)(3);
  VNStageIntLLRInputS7xD(265)(2) <= CNStageIntLLROutputS7xD(203)(4);
  VNStageIntLLRInputS7xD(326)(2) <= CNStageIntLLROutputS7xD(203)(5);
  VNStageIntLLRInputS7xD(23)(3) <= CNStageIntLLROutputS7xD(204)(0);
  VNStageIntLLRInputS7xD(88)(3) <= CNStageIntLLROutputS7xD(204)(1);
  VNStageIntLLRInputS7xD(177)(3) <= CNStageIntLLROutputS7xD(204)(2);
  VNStageIntLLRInputS7xD(200)(3) <= CNStageIntLLROutputS7xD(204)(3);
  VNStageIntLLRInputS7xD(261)(3) <= CNStageIntLLROutputS7xD(204)(4);
  VNStageIntLLRInputS7xD(341)(3) <= CNStageIntLLROutputS7xD(204)(5);
  VNStageIntLLRInputS7xD(22)(3) <= CNStageIntLLROutputS7xD(205)(0);
  VNStageIntLLRInputS7xD(112)(3) <= CNStageIntLLROutputS7xD(205)(1);
  VNStageIntLLRInputS7xD(135)(3) <= CNStageIntLLROutputS7xD(205)(2);
  VNStageIntLLRInputS7xD(196)(3) <= CNStageIntLLROutputS7xD(205)(3);
  VNStageIntLLRInputS7xD(276)(3) <= CNStageIntLLROutputS7xD(205)(4);
  VNStageIntLLRInputS7xD(367)(3) <= CNStageIntLLROutputS7xD(205)(5);
  VNStageIntLLRInputS7xD(21)(3) <= CNStageIntLLROutputS7xD(206)(0);
  VNStageIntLLRInputS7xD(70)(3) <= CNStageIntLLROutputS7xD(206)(1);
  VNStageIntLLRInputS7xD(131)(2) <= CNStageIntLLROutputS7xD(206)(2);
  VNStageIntLLRInputS7xD(211)(3) <= CNStageIntLLROutputS7xD(206)(3);
  VNStageIntLLRInputS7xD(302)(3) <= CNStageIntLLROutputS7xD(206)(4);
  VNStageIntLLRInputS7xD(343)(3) <= CNStageIntLLROutputS7xD(206)(5);
  VNStageIntLLRInputS7xD(18)(3) <= CNStageIntLLROutputS7xD(207)(0);
  VNStageIntLLRInputS7xD(107)(2) <= CNStageIntLLROutputS7xD(207)(1);
  VNStageIntLLRInputS7xD(148)(3) <= CNStageIntLLROutputS7xD(207)(2);
  VNStageIntLLRInputS7xD(245)(3) <= CNStageIntLLROutputS7xD(207)(3);
  VNStageIntLLRInputS7xD(263)(3) <= CNStageIntLLROutputS7xD(207)(4);
  VNStageIntLLRInputS7xD(361)(3) <= CNStageIntLLROutputS7xD(207)(5);
  VNStageIntLLRInputS7xD(17)(3) <= CNStageIntLLROutputS7xD(208)(0);
  VNStageIntLLRInputS7xD(83)(3) <= CNStageIntLLROutputS7xD(208)(1);
  VNStageIntLLRInputS7xD(180)(1) <= CNStageIntLLROutputS7xD(208)(2);
  VNStageIntLLRInputS7xD(198)(3) <= CNStageIntLLROutputS7xD(208)(3);
  VNStageIntLLRInputS7xD(296)(3) <= CNStageIntLLROutputS7xD(208)(4);
  VNStageIntLLRInputS7xD(370)(2) <= CNStageIntLLROutputS7xD(208)(5);
  VNStageIntLLRInputS7xD(16)(2) <= CNStageIntLLROutputS7xD(209)(0);
  VNStageIntLLRInputS7xD(115)(3) <= CNStageIntLLROutputS7xD(209)(1);
  VNStageIntLLRInputS7xD(133)(1) <= CNStageIntLLROutputS7xD(209)(2);
  VNStageIntLLRInputS7xD(231)(2) <= CNStageIntLLROutputS7xD(209)(3);
  VNStageIntLLRInputS7xD(305)(3) <= CNStageIntLLROutputS7xD(209)(4);
  VNStageIntLLRInputS7xD(383)(3) <= CNStageIntLLROutputS7xD(209)(5);
  VNStageIntLLRInputS7xD(15)(3) <= CNStageIntLLROutputS7xD(210)(0);
  VNStageIntLLRInputS7xD(68)(2) <= CNStageIntLLROutputS7xD(210)(1);
  VNStageIntLLRInputS7xD(166)(3) <= CNStageIntLLROutputS7xD(210)(2);
  VNStageIntLLRInputS7xD(240)(3) <= CNStageIntLLROutputS7xD(210)(3);
  VNStageIntLLRInputS7xD(318)(1) <= CNStageIntLLROutputS7xD(210)(4);
  VNStageIntLLRInputS7xD(362)(3) <= CNStageIntLLROutputS7xD(210)(5);
  VNStageIntLLRInputS7xD(14)(3) <= CNStageIntLLROutputS7xD(211)(0);
  VNStageIntLLRInputS7xD(101)(3) <= CNStageIntLLROutputS7xD(211)(1);
  VNStageIntLLRInputS7xD(175)(3) <= CNStageIntLLROutputS7xD(211)(2);
  VNStageIntLLRInputS7xD(253)(2) <= CNStageIntLLROutputS7xD(211)(3);
  VNStageIntLLRInputS7xD(297)(3) <= CNStageIntLLROutputS7xD(211)(4);
  VNStageIntLLRInputS7xD(327)(3) <= CNStageIntLLROutputS7xD(211)(5);
  VNStageIntLLRInputS7xD(13)(2) <= CNStageIntLLROutputS7xD(212)(0);
  VNStageIntLLRInputS7xD(110)(3) <= CNStageIntLLROutputS7xD(212)(1);
  VNStageIntLLRInputS7xD(188)(1) <= CNStageIntLLROutputS7xD(212)(2);
  VNStageIntLLRInputS7xD(232)(2) <= CNStageIntLLROutputS7xD(212)(3);
  VNStageIntLLRInputS7xD(262)(3) <= CNStageIntLLROutputS7xD(212)(4);
  VNStageIntLLRInputS7xD(329)(3) <= CNStageIntLLROutputS7xD(212)(5);
  VNStageIntLLRInputS7xD(12)(3) <= CNStageIntLLROutputS7xD(213)(0);
  VNStageIntLLRInputS7xD(123)(2) <= CNStageIntLLROutputS7xD(213)(1);
  VNStageIntLLRInputS7xD(167)(3) <= CNStageIntLLROutputS7xD(213)(2);
  VNStageIntLLRInputS7xD(197)(3) <= CNStageIntLLROutputS7xD(213)(3);
  VNStageIntLLRInputS7xD(264)(3) <= CNStageIntLLROutputS7xD(213)(4);
  VNStageIntLLRInputS7xD(374)(3) <= CNStageIntLLROutputS7xD(213)(5);
  VNStageIntLLRInputS7xD(11)(3) <= CNStageIntLLROutputS7xD(214)(0);
  VNStageIntLLRInputS7xD(102)(3) <= CNStageIntLLROutputS7xD(214)(1);
  VNStageIntLLRInputS7xD(132)(2) <= CNStageIntLLROutputS7xD(214)(2);
  VNStageIntLLRInputS7xD(199)(3) <= CNStageIntLLROutputS7xD(214)(3);
  VNStageIntLLRInputS7xD(309)(3) <= CNStageIntLLROutputS7xD(214)(4);
  VNStageIntLLRInputS7xD(381)(2) <= CNStageIntLLROutputS7xD(214)(5);
  VNStageIntLLRInputS7xD(9)(3) <= CNStageIntLLROutputS7xD(215)(0);
  VNStageIntLLRInputS7xD(69)(3) <= CNStageIntLLROutputS7xD(215)(1);
  VNStageIntLLRInputS7xD(179)(3) <= CNStageIntLLROutputS7xD(215)(2);
  VNStageIntLLRInputS7xD(251)(2) <= CNStageIntLLROutputS7xD(215)(3);
  VNStageIntLLRInputS7xD(280)(3) <= CNStageIntLLROutputS7xD(215)(4);
  VNStageIntLLRInputS7xD(333)(2) <= CNStageIntLLROutputS7xD(215)(5);
  VNStageIntLLRInputS7xD(8)(2) <= CNStageIntLLROutputS7xD(216)(0);
  VNStageIntLLRInputS7xD(114)(3) <= CNStageIntLLROutputS7xD(216)(1);
  VNStageIntLLRInputS7xD(186)(2) <= CNStageIntLLROutputS7xD(216)(2);
  VNStageIntLLRInputS7xD(215)(3) <= CNStageIntLLROutputS7xD(216)(3);
  VNStageIntLLRInputS7xD(268)(3) <= CNStageIntLLROutputS7xD(216)(4);
  VNStageIntLLRInputS7xD(339)(3) <= CNStageIntLLROutputS7xD(216)(5);
  VNStageIntLLRInputS7xD(7)(3) <= CNStageIntLLROutputS7xD(217)(0);
  VNStageIntLLRInputS7xD(121)(2) <= CNStageIntLLROutputS7xD(217)(1);
  VNStageIntLLRInputS7xD(150)(3) <= CNStageIntLLROutputS7xD(217)(2);
  VNStageIntLLRInputS7xD(203)(3) <= CNStageIntLLROutputS7xD(217)(3);
  VNStageIntLLRInputS7xD(274)(2) <= CNStageIntLLROutputS7xD(217)(4);
  VNStageIntLLRInputS7xD(334)(2) <= CNStageIntLLROutputS7xD(217)(5);
  VNStageIntLLRInputS7xD(6)(3) <= CNStageIntLLROutputS7xD(218)(0);
  VNStageIntLLRInputS7xD(85)(2) <= CNStageIntLLROutputS7xD(218)(1);
  VNStageIntLLRInputS7xD(138)(3) <= CNStageIntLLROutputS7xD(218)(2);
  VNStageIntLLRInputS7xD(209)(3) <= CNStageIntLLROutputS7xD(218)(3);
  VNStageIntLLRInputS7xD(269)(2) <= CNStageIntLLROutputS7xD(218)(4);
  VNStageIntLLRInputS7xD(344)(3) <= CNStageIntLLROutputS7xD(218)(5);
  VNStageIntLLRInputS7xD(5)(3) <= CNStageIntLLROutputS7xD(219)(0);
  VNStageIntLLRInputS7xD(73)(3) <= CNStageIntLLROutputS7xD(219)(1);
  VNStageIntLLRInputS7xD(144)(3) <= CNStageIntLLROutputS7xD(219)(2);
  VNStageIntLLRInputS7xD(204)(3) <= CNStageIntLLROutputS7xD(219)(3);
  VNStageIntLLRInputS7xD(279)(3) <= CNStageIntLLROutputS7xD(219)(4);
  VNStageIntLLRInputS7xD(366)(3) <= CNStageIntLLROutputS7xD(219)(5);
  VNStageIntLLRInputS7xD(4)(2) <= CNStageIntLLROutputS7xD(220)(0);
  VNStageIntLLRInputS7xD(79)(3) <= CNStageIntLLROutputS7xD(220)(1);
  VNStageIntLLRInputS7xD(139)(3) <= CNStageIntLLROutputS7xD(220)(2);
  VNStageIntLLRInputS7xD(214)(3) <= CNStageIntLLROutputS7xD(220)(3);
  VNStageIntLLRInputS7xD(301)(3) <= CNStageIntLLROutputS7xD(220)(4);
  VNStageIntLLRInputS7xD(321)(3) <= CNStageIntLLROutputS7xD(220)(5);
  VNStageIntLLRInputS7xD(3)(2) <= CNStageIntLLROutputS7xD(221)(0);
  VNStageIntLLRInputS7xD(74)(3) <= CNStageIntLLROutputS7xD(221)(1);
  VNStageIntLLRInputS7xD(149)(3) <= CNStageIntLLROutputS7xD(221)(2);
  VNStageIntLLRInputS7xD(236)(3) <= CNStageIntLLROutputS7xD(221)(3);
  VNStageIntLLRInputS7xD(319)(3) <= CNStageIntLLROutputS7xD(221)(4);
  VNStageIntLLRInputS7xD(369)(2) <= CNStageIntLLROutputS7xD(221)(5);
  VNStageIntLLRInputS7xD(2)(3) <= CNStageIntLLROutputS7xD(222)(0);
  VNStageIntLLRInputS7xD(84)(3) <= CNStageIntLLROutputS7xD(222)(1);
  VNStageIntLLRInputS7xD(171)(2) <= CNStageIntLLROutputS7xD(222)(2);
  VNStageIntLLRInputS7xD(254)(1) <= CNStageIntLLROutputS7xD(222)(3);
  VNStageIntLLRInputS7xD(304)(3) <= CNStageIntLLROutputS7xD(222)(4);
  VNStageIntLLRInputS7xD(356)(3) <= CNStageIntLLROutputS7xD(222)(5);
  VNStageIntLLRInputS7xD(1)(2) <= CNStageIntLLROutputS7xD(223)(0);
  VNStageIntLLRInputS7xD(106)(2) <= CNStageIntLLROutputS7xD(223)(1);
  VNStageIntLLRInputS7xD(189)(2) <= CNStageIntLLROutputS7xD(223)(2);
  VNStageIntLLRInputS7xD(239)(3) <= CNStageIntLLROutputS7xD(223)(3);
  VNStageIntLLRInputS7xD(291)(3) <= CNStageIntLLROutputS7xD(223)(4);
  VNStageIntLLRInputS7xD(324)(3) <= CNStageIntLLROutputS7xD(223)(5);
  VNStageIntLLRInputS7xD(0)(3) <= CNStageIntLLROutputS7xD(224)(0);
  VNStageIntLLRInputS7xD(93)(3) <= CNStageIntLLROutputS7xD(224)(1);
  VNStageIntLLRInputS7xD(158)(3) <= CNStageIntLLROutputS7xD(224)(2);
  VNStageIntLLRInputS7xD(223)(3) <= CNStageIntLLROutputS7xD(224)(3);
  VNStageIntLLRInputS7xD(288)(3) <= CNStageIntLLROutputS7xD(224)(4);
  VNStageIntLLRInputS7xD(353)(3) <= CNStageIntLLROutputS7xD(224)(5);
  VNStageIntLLRInputS7xD(18)(4) <= CNStageIntLLROutputS7xD(225)(0);
  VNStageIntLLRInputS7xD(110)(4) <= CNStageIntLLROutputS7xD(225)(1);
  VNStageIntLLRInputS7xD(167)(4) <= CNStageIntLLROutputS7xD(225)(2);
  VNStageIntLLRInputS7xD(249)(2) <= CNStageIntLLROutputS7xD(225)(3);
  VNStageIntLLRInputS7xD(311)(3) <= CNStageIntLLROutputS7xD(225)(4);
  VNStageIntLLRInputS7xD(347)(4) <= CNStageIntLLROutputS7xD(225)(5);
  VNStageIntLLRInputS7xD(17)(4) <= CNStageIntLLROutputS7xD(226)(0);
  VNStageIntLLRInputS7xD(102)(4) <= CNStageIntLLROutputS7xD(226)(1);
  VNStageIntLLRInputS7xD(184)(4) <= CNStageIntLLROutputS7xD(226)(2);
  VNStageIntLLRInputS7xD(246)(4) <= CNStageIntLLROutputS7xD(226)(3);
  VNStageIntLLRInputS7xD(282)(4) <= CNStageIntLLROutputS7xD(226)(4);
  VNStageIntLLRInputS7xD(367)(4) <= CNStageIntLLROutputS7xD(226)(5);
  VNStageIntLLRInputS7xD(16)(3) <= CNStageIntLLROutputS7xD(227)(0);
  VNStageIntLLRInputS7xD(119)(3) <= CNStageIntLLROutputS7xD(227)(1);
  VNStageIntLLRInputS7xD(181)(4) <= CNStageIntLLROutputS7xD(227)(2);
  VNStageIntLLRInputS7xD(217)(4) <= CNStageIntLLROutputS7xD(227)(3);
  VNStageIntLLRInputS7xD(302)(4) <= CNStageIntLLROutputS7xD(227)(4);
  VNStageIntLLRInputS7xD(353)(4) <= CNStageIntLLROutputS7xD(227)(5);
  VNStageIntLLRInputS7xD(15)(4) <= CNStageIntLLROutputS7xD(228)(0);
  VNStageIntLLRInputS7xD(116)(3) <= CNStageIntLLROutputS7xD(228)(1);
  VNStageIntLLRInputS7xD(152)(4) <= CNStageIntLLROutputS7xD(228)(2);
  VNStageIntLLRInputS7xD(237)(3) <= CNStageIntLLROutputS7xD(228)(3);
  VNStageIntLLRInputS7xD(288)(4) <= CNStageIntLLROutputS7xD(228)(4);
  VNStageIntLLRInputS7xD(343)(4) <= CNStageIntLLROutputS7xD(228)(5);
  VNStageIntLLRInputS7xD(14)(4) <= CNStageIntLLROutputS7xD(229)(0);
  VNStageIntLLRInputS7xD(87)(4) <= CNStageIntLLROutputS7xD(229)(1);
  VNStageIntLLRInputS7xD(172)(3) <= CNStageIntLLROutputS7xD(229)(2);
  VNStageIntLLRInputS7xD(223)(4) <= CNStageIntLLROutputS7xD(229)(3);
  VNStageIntLLRInputS7xD(278)(3) <= CNStageIntLLROutputS7xD(229)(4);
  VNStageIntLLRInputS7xD(372)(3) <= CNStageIntLLROutputS7xD(229)(5);
  VNStageIntLLRInputS7xD(13)(3) <= CNStageIntLLROutputS7xD(230)(0);
  VNStageIntLLRInputS7xD(107)(3) <= CNStageIntLLROutputS7xD(230)(1);
  VNStageIntLLRInputS7xD(158)(4) <= CNStageIntLLROutputS7xD(230)(2);
  VNStageIntLLRInputS7xD(213)(3) <= CNStageIntLLROutputS7xD(230)(3);
  VNStageIntLLRInputS7xD(307)(4) <= CNStageIntLLROutputS7xD(230)(4);
  VNStageIntLLRInputS7xD(355)(4) <= CNStageIntLLROutputS7xD(230)(5);
  VNStageIntLLRInputS7xD(12)(4) <= CNStageIntLLROutputS7xD(231)(0);
  VNStageIntLLRInputS7xD(93)(4) <= CNStageIntLLROutputS7xD(231)(1);
  VNStageIntLLRInputS7xD(148)(4) <= CNStageIntLLROutputS7xD(231)(2);
  VNStageIntLLRInputS7xD(242)(4) <= CNStageIntLLROutputS7xD(231)(3);
  VNStageIntLLRInputS7xD(290)(4) <= CNStageIntLLROutputS7xD(231)(4);
  VNStageIntLLRInputS7xD(322)(3) <= CNStageIntLLROutputS7xD(231)(5);
  VNStageIntLLRInputS7xD(11)(4) <= CNStageIntLLROutputS7xD(232)(0);
  VNStageIntLLRInputS7xD(83)(4) <= CNStageIntLLROutputS7xD(232)(1);
  VNStageIntLLRInputS7xD(177)(4) <= CNStageIntLLROutputS7xD(232)(2);
  VNStageIntLLRInputS7xD(225)(4) <= CNStageIntLLROutputS7xD(232)(3);
  VNStageIntLLRInputS7xD(257)(4) <= CNStageIntLLROutputS7xD(232)(4);
  VNStageIntLLRInputS7xD(345)(3) <= CNStageIntLLROutputS7xD(232)(5);
  VNStageIntLLRInputS7xD(10)(3) <= CNStageIntLLROutputS7xD(233)(0);
  VNStageIntLLRInputS7xD(112)(4) <= CNStageIntLLROutputS7xD(233)(1);
  VNStageIntLLRInputS7xD(160)(4) <= CNStageIntLLROutputS7xD(233)(2);
  VNStageIntLLRInputS7xD(255)(4) <= CNStageIntLLROutputS7xD(233)(3);
  VNStageIntLLRInputS7xD(280)(4) <= CNStageIntLLROutputS7xD(233)(4);
  VNStageIntLLRInputS7xD(381)(3) <= CNStageIntLLROutputS7xD(233)(5);
  VNStageIntLLRInputS7xD(9)(4) <= CNStageIntLLROutputS7xD(234)(0);
  VNStageIntLLRInputS7xD(95)(4) <= CNStageIntLLROutputS7xD(234)(1);
  VNStageIntLLRInputS7xD(190)(2) <= CNStageIntLLROutputS7xD(234)(2);
  VNStageIntLLRInputS7xD(215)(4) <= CNStageIntLLROutputS7xD(234)(3);
  VNStageIntLLRInputS7xD(316)(2) <= CNStageIntLLROutputS7xD(234)(4);
  VNStageIntLLRInputS7xD(365)(4) <= CNStageIntLLROutputS7xD(234)(5);
  VNStageIntLLRInputS7xD(7)(4) <= CNStageIntLLROutputS7xD(235)(0);
  VNStageIntLLRInputS7xD(85)(3) <= CNStageIntLLROutputS7xD(235)(1);
  VNStageIntLLRInputS7xD(186)(3) <= CNStageIntLLROutputS7xD(235)(2);
  VNStageIntLLRInputS7xD(235)(3) <= CNStageIntLLROutputS7xD(235)(3);
  VNStageIntLLRInputS7xD(303)(4) <= CNStageIntLLROutputS7xD(235)(4);
  VNStageIntLLRInputS7xD(346)(4) <= CNStageIntLLROutputS7xD(235)(5);
  VNStageIntLLRInputS7xD(6)(4) <= CNStageIntLLROutputS7xD(236)(0);
  VNStageIntLLRInputS7xD(121)(3) <= CNStageIntLLROutputS7xD(236)(1);
  VNStageIntLLRInputS7xD(170)(3) <= CNStageIntLLROutputS7xD(236)(2);
  VNStageIntLLRInputS7xD(238)(4) <= CNStageIntLLROutputS7xD(236)(3);
  VNStageIntLLRInputS7xD(281)(4) <= CNStageIntLLROutputS7xD(236)(4);
  VNStageIntLLRInputS7xD(321)(4) <= CNStageIntLLROutputS7xD(236)(5);
  VNStageIntLLRInputS7xD(5)(4) <= CNStageIntLLROutputS7xD(237)(0);
  VNStageIntLLRInputS7xD(105)(3) <= CNStageIntLLROutputS7xD(237)(1);
  VNStageIntLLRInputS7xD(173)(4) <= CNStageIntLLROutputS7xD(237)(2);
  VNStageIntLLRInputS7xD(216)(4) <= CNStageIntLLROutputS7xD(237)(3);
  VNStageIntLLRInputS7xD(319)(4) <= CNStageIntLLROutputS7xD(237)(4);
  VNStageIntLLRInputS7xD(382)(3) <= CNStageIntLLROutputS7xD(237)(5);
  VNStageIntLLRInputS7xD(4)(3) <= CNStageIntLLROutputS7xD(238)(0);
  VNStageIntLLRInputS7xD(108)(4) <= CNStageIntLLROutputS7xD(238)(1);
  VNStageIntLLRInputS7xD(151)(4) <= CNStageIntLLROutputS7xD(238)(2);
  VNStageIntLLRInputS7xD(254)(2) <= CNStageIntLLROutputS7xD(238)(3);
  VNStageIntLLRInputS7xD(317)(1) <= CNStageIntLLROutputS7xD(238)(4);
  VNStageIntLLRInputS7xD(344)(4) <= CNStageIntLLROutputS7xD(238)(5);
  VNStageIntLLRInputS7xD(3)(3) <= CNStageIntLLROutputS7xD(239)(0);
  VNStageIntLLRInputS7xD(86)(2) <= CNStageIntLLROutputS7xD(239)(1);
  VNStageIntLLRInputS7xD(189)(3) <= CNStageIntLLROutputS7xD(239)(2);
  VNStageIntLLRInputS7xD(252)(3) <= CNStageIntLLROutputS7xD(239)(3);
  VNStageIntLLRInputS7xD(279)(4) <= CNStageIntLLROutputS7xD(239)(4);
  VNStageIntLLRInputS7xD(352)(4) <= CNStageIntLLROutputS7xD(239)(5);
  VNStageIntLLRInputS7xD(2)(4) <= CNStageIntLLROutputS7xD(240)(0);
  VNStageIntLLRInputS7xD(124)(2) <= CNStageIntLLROutputS7xD(240)(1);
  VNStageIntLLRInputS7xD(187)(3) <= CNStageIntLLROutputS7xD(240)(2);
  VNStageIntLLRInputS7xD(214)(4) <= CNStageIntLLROutputS7xD(240)(3);
  VNStageIntLLRInputS7xD(287)(4) <= CNStageIntLLROutputS7xD(240)(4);
  VNStageIntLLRInputS7xD(332)(4) <= CNStageIntLLROutputS7xD(240)(5);
  VNStageIntLLRInputS7xD(1)(3) <= CNStageIntLLROutputS7xD(241)(0);
  VNStageIntLLRInputS7xD(122)(3) <= CNStageIntLLROutputS7xD(241)(1);
  VNStageIntLLRInputS7xD(149)(4) <= CNStageIntLLROutputS7xD(241)(2);
  VNStageIntLLRInputS7xD(222)(2) <= CNStageIntLLROutputS7xD(241)(3);
  VNStageIntLLRInputS7xD(267)(4) <= CNStageIntLLROutputS7xD(241)(4);
  VNStageIntLLRInputS7xD(326)(3) <= CNStageIntLLROutputS7xD(241)(5);
  VNStageIntLLRInputS7xD(62)(3) <= CNStageIntLLROutputS7xD(242)(0);
  VNStageIntLLRInputS7xD(92)(4) <= CNStageIntLLROutputS7xD(242)(1);
  VNStageIntLLRInputS7xD(137)(4) <= CNStageIntLLROutputS7xD(242)(2);
  VNStageIntLLRInputS7xD(196)(4) <= CNStageIntLLROutputS7xD(242)(3);
  VNStageIntLLRInputS7xD(256)(3) <= CNStageIntLLROutputS7xD(242)(4);
  VNStageIntLLRInputS7xD(325)(4) <= CNStageIntLLROutputS7xD(242)(5);
  VNStageIntLLRInputS7xD(61)(3) <= CNStageIntLLROutputS7xD(243)(0);
  VNStageIntLLRInputS7xD(72)(4) <= CNStageIntLLROutputS7xD(243)(1);
  VNStageIntLLRInputS7xD(131)(3) <= CNStageIntLLROutputS7xD(243)(2);
  VNStageIntLLRInputS7xD(192)(4) <= CNStageIntLLROutputS7xD(243)(3);
  VNStageIntLLRInputS7xD(260)(4) <= CNStageIntLLROutputS7xD(243)(4);
  VNStageIntLLRInputS7xD(330)(4) <= CNStageIntLLROutputS7xD(243)(5);
  VNStageIntLLRInputS7xD(60)(3) <= CNStageIntLLROutputS7xD(244)(0);
  VNStageIntLLRInputS7xD(66)(3) <= CNStageIntLLROutputS7xD(244)(1);
  VNStageIntLLRInputS7xD(128)(4) <= CNStageIntLLROutputS7xD(244)(2);
  VNStageIntLLRInputS7xD(195)(3) <= CNStageIntLLROutputS7xD(244)(3);
  VNStageIntLLRInputS7xD(265)(3) <= CNStageIntLLROutputS7xD(244)(4);
  VNStageIntLLRInputS7xD(349)(3) <= CNStageIntLLROutputS7xD(244)(5);
  VNStageIntLLRInputS7xD(59)(2) <= CNStageIntLLROutputS7xD(245)(0);
  VNStageIntLLRInputS7xD(64)(3) <= CNStageIntLLROutputS7xD(245)(1);
  VNStageIntLLRInputS7xD(130)(4) <= CNStageIntLLROutputS7xD(245)(2);
  VNStageIntLLRInputS7xD(200)(4) <= CNStageIntLLROutputS7xD(245)(3);
  VNStageIntLLRInputS7xD(284)(4) <= CNStageIntLLROutputS7xD(245)(4);
  VNStageIntLLRInputS7xD(340)(4) <= CNStageIntLLROutputS7xD(245)(5);
  VNStageIntLLRInputS7xD(57)(3) <= CNStageIntLLROutputS7xD(246)(0);
  VNStageIntLLRInputS7xD(70)(4) <= CNStageIntLLROutputS7xD(246)(1);
  VNStageIntLLRInputS7xD(154)(3) <= CNStageIntLLROutputS7xD(246)(2);
  VNStageIntLLRInputS7xD(210)(4) <= CNStageIntLLROutputS7xD(246)(3);
  VNStageIntLLRInputS7xD(312)(3) <= CNStageIntLLROutputS7xD(246)(4);
  VNStageIntLLRInputS7xD(378)(3) <= CNStageIntLLROutputS7xD(246)(5);
  VNStageIntLLRInputS7xD(56)(4) <= CNStageIntLLROutputS7xD(247)(0);
  VNStageIntLLRInputS7xD(89)(4) <= CNStageIntLLROutputS7xD(247)(1);
  VNStageIntLLRInputS7xD(145)(4) <= CNStageIntLLROutputS7xD(247)(2);
  VNStageIntLLRInputS7xD(247)(4) <= CNStageIntLLROutputS7xD(247)(3);
  VNStageIntLLRInputS7xD(313)(2) <= CNStageIntLLROutputS7xD(247)(4);
  VNStageIntLLRInputS7xD(339)(4) <= CNStageIntLLROutputS7xD(247)(5);
  VNStageIntLLRInputS7xD(55)(4) <= CNStageIntLLROutputS7xD(248)(0);
  VNStageIntLLRInputS7xD(80)(4) <= CNStageIntLLROutputS7xD(248)(1);
  VNStageIntLLRInputS7xD(182)(4) <= CNStageIntLLROutputS7xD(248)(2);
  VNStageIntLLRInputS7xD(248)(4) <= CNStageIntLLROutputS7xD(248)(3);
  VNStageIntLLRInputS7xD(274)(3) <= CNStageIntLLROutputS7xD(248)(4);
  VNStageIntLLRInputS7xD(360)(4) <= CNStageIntLLROutputS7xD(248)(5);
  VNStageIntLLRInputS7xD(53)(3) <= CNStageIntLLROutputS7xD(249)(0);
  VNStageIntLLRInputS7xD(118)(3) <= CNStageIntLLROutputS7xD(249)(1);
  VNStageIntLLRInputS7xD(144)(4) <= CNStageIntLLROutputS7xD(249)(2);
  VNStageIntLLRInputS7xD(230)(3) <= CNStageIntLLROutputS7xD(249)(3);
  VNStageIntLLRInputS7xD(291)(4) <= CNStageIntLLROutputS7xD(249)(4);
  VNStageIntLLRInputS7xD(371)(3) <= CNStageIntLLROutputS7xD(249)(5);
  VNStageIntLLRInputS7xD(51)(3) <= CNStageIntLLROutputS7xD(250)(0);
  VNStageIntLLRInputS7xD(100)(4) <= CNStageIntLLROutputS7xD(250)(1);
  VNStageIntLLRInputS7xD(161)(4) <= CNStageIntLLROutputS7xD(250)(2);
  VNStageIntLLRInputS7xD(241)(3) <= CNStageIntLLROutputS7xD(250)(3);
  VNStageIntLLRInputS7xD(269)(3) <= CNStageIntLLROutputS7xD(250)(4);
  VNStageIntLLRInputS7xD(373)(2) <= CNStageIntLLROutputS7xD(250)(5);
  VNStageIntLLRInputS7xD(50)(4) <= CNStageIntLLROutputS7xD(251)(0);
  VNStageIntLLRInputS7xD(96)(4) <= CNStageIntLLROutputS7xD(251)(1);
  VNStageIntLLRInputS7xD(176)(4) <= CNStageIntLLROutputS7xD(251)(2);
  VNStageIntLLRInputS7xD(204)(4) <= CNStageIntLLROutputS7xD(251)(3);
  VNStageIntLLRInputS7xD(308)(2) <= CNStageIntLLROutputS7xD(251)(4);
  VNStageIntLLRInputS7xD(342)(3) <= CNStageIntLLROutputS7xD(251)(5);
  VNStageIntLLRInputS7xD(49)(4) <= CNStageIntLLROutputS7xD(252)(0);
  VNStageIntLLRInputS7xD(111)(4) <= CNStageIntLLROutputS7xD(252)(1);
  VNStageIntLLRInputS7xD(139)(4) <= CNStageIntLLROutputS7xD(252)(2);
  VNStageIntLLRInputS7xD(243)(4) <= CNStageIntLLROutputS7xD(252)(3);
  VNStageIntLLRInputS7xD(277)(4) <= CNStageIntLLROutputS7xD(252)(4);
  VNStageIntLLRInputS7xD(358)(3) <= CNStageIntLLROutputS7xD(252)(5);
  VNStageIntLLRInputS7xD(47)(2) <= CNStageIntLLROutputS7xD(253)(0);
  VNStageIntLLRInputS7xD(113)(4) <= CNStageIntLLROutputS7xD(253)(1);
  VNStageIntLLRInputS7xD(147)(4) <= CNStageIntLLROutputS7xD(253)(2);
  VNStageIntLLRInputS7xD(228)(4) <= CNStageIntLLROutputS7xD(253)(3);
  VNStageIntLLRInputS7xD(263)(4) <= CNStageIntLLROutputS7xD(253)(4);
  VNStageIntLLRInputS7xD(337)(4) <= CNStageIntLLROutputS7xD(253)(5);
  VNStageIntLLRInputS7xD(46)(4) <= CNStageIntLLROutputS7xD(254)(0);
  VNStageIntLLRInputS7xD(82)(4) <= CNStageIntLLROutputS7xD(254)(1);
  VNStageIntLLRInputS7xD(163)(3) <= CNStageIntLLROutputS7xD(254)(2);
  VNStageIntLLRInputS7xD(198)(4) <= CNStageIntLLROutputS7xD(254)(3);
  VNStageIntLLRInputS7xD(272)(4) <= CNStageIntLLROutputS7xD(254)(4);
  VNStageIntLLRInputS7xD(350)(4) <= CNStageIntLLROutputS7xD(254)(5);
  VNStageIntLLRInputS7xD(45)(4) <= CNStageIntLLROutputS7xD(255)(0);
  VNStageIntLLRInputS7xD(98)(3) <= CNStageIntLLROutputS7xD(255)(1);
  VNStageIntLLRInputS7xD(133)(2) <= CNStageIntLLROutputS7xD(255)(2);
  VNStageIntLLRInputS7xD(207)(3) <= CNStageIntLLROutputS7xD(255)(3);
  VNStageIntLLRInputS7xD(285)(4) <= CNStageIntLLROutputS7xD(255)(4);
  VNStageIntLLRInputS7xD(329)(4) <= CNStageIntLLROutputS7xD(255)(5);
  VNStageIntLLRInputS7xD(44)(4) <= CNStageIntLLROutputS7xD(256)(0);
  VNStageIntLLRInputS7xD(68)(3) <= CNStageIntLLROutputS7xD(256)(1);
  VNStageIntLLRInputS7xD(142)(3) <= CNStageIntLLROutputS7xD(256)(2);
  VNStageIntLLRInputS7xD(220)(4) <= CNStageIntLLROutputS7xD(256)(3);
  VNStageIntLLRInputS7xD(264)(4) <= CNStageIntLLROutputS7xD(256)(4);
  VNStageIntLLRInputS7xD(357)(4) <= CNStageIntLLROutputS7xD(256)(5);
  VNStageIntLLRInputS7xD(43)(3) <= CNStageIntLLROutputS7xD(257)(0);
  VNStageIntLLRInputS7xD(77)(2) <= CNStageIntLLROutputS7xD(257)(1);
  VNStageIntLLRInputS7xD(155)(4) <= CNStageIntLLROutputS7xD(257)(2);
  VNStageIntLLRInputS7xD(199)(4) <= CNStageIntLLROutputS7xD(257)(3);
  VNStageIntLLRInputS7xD(292)(4) <= CNStageIntLLROutputS7xD(257)(4);
  VNStageIntLLRInputS7xD(359)(4) <= CNStageIntLLROutputS7xD(257)(5);
  VNStageIntLLRInputS7xD(42)(4) <= CNStageIntLLROutputS7xD(258)(0);
  VNStageIntLLRInputS7xD(90)(4) <= CNStageIntLLROutputS7xD(258)(1);
  VNStageIntLLRInputS7xD(134)(3) <= CNStageIntLLROutputS7xD(258)(2);
  VNStageIntLLRInputS7xD(227)(4) <= CNStageIntLLROutputS7xD(258)(3);
  VNStageIntLLRInputS7xD(294)(4) <= CNStageIntLLROutputS7xD(258)(4);
  VNStageIntLLRInputS7xD(341)(4) <= CNStageIntLLROutputS7xD(258)(5);
  VNStageIntLLRInputS7xD(41)(4) <= CNStageIntLLROutputS7xD(259)(0);
  VNStageIntLLRInputS7xD(69)(4) <= CNStageIntLLROutputS7xD(259)(1);
  VNStageIntLLRInputS7xD(162)(4) <= CNStageIntLLROutputS7xD(259)(2);
  VNStageIntLLRInputS7xD(229)(3) <= CNStageIntLLROutputS7xD(259)(3);
  VNStageIntLLRInputS7xD(276)(4) <= CNStageIntLLROutputS7xD(259)(4);
  VNStageIntLLRInputS7xD(348)(4) <= CNStageIntLLROutputS7xD(259)(5);
  VNStageIntLLRInputS7xD(40)(3) <= CNStageIntLLROutputS7xD(260)(0);
  VNStageIntLLRInputS7xD(97)(4) <= CNStageIntLLROutputS7xD(260)(1);
  VNStageIntLLRInputS7xD(164)(4) <= CNStageIntLLROutputS7xD(260)(2);
  VNStageIntLLRInputS7xD(211)(4) <= CNStageIntLLROutputS7xD(260)(3);
  VNStageIntLLRInputS7xD(283)(4) <= CNStageIntLLROutputS7xD(260)(4);
  VNStageIntLLRInputS7xD(375)(3) <= CNStageIntLLROutputS7xD(260)(5);
  VNStageIntLLRInputS7xD(39)(4) <= CNStageIntLLROutputS7xD(261)(0);
  VNStageIntLLRInputS7xD(99)(4) <= CNStageIntLLROutputS7xD(261)(1);
  VNStageIntLLRInputS7xD(146)(3) <= CNStageIntLLROutputS7xD(261)(2);
  VNStageIntLLRInputS7xD(218)(4) <= CNStageIntLLROutputS7xD(261)(3);
  VNStageIntLLRInputS7xD(310)(3) <= CNStageIntLLROutputS7xD(261)(4);
  VNStageIntLLRInputS7xD(363)(3) <= CNStageIntLLROutputS7xD(261)(5);
  VNStageIntLLRInputS7xD(38)(4) <= CNStageIntLLROutputS7xD(262)(0);
  VNStageIntLLRInputS7xD(81)(3) <= CNStageIntLLROutputS7xD(262)(1);
  VNStageIntLLRInputS7xD(153)(4) <= CNStageIntLLROutputS7xD(262)(2);
  VNStageIntLLRInputS7xD(245)(4) <= CNStageIntLLROutputS7xD(262)(3);
  VNStageIntLLRInputS7xD(298)(4) <= CNStageIntLLROutputS7xD(262)(4);
  VNStageIntLLRInputS7xD(369)(3) <= CNStageIntLLROutputS7xD(262)(5);
  VNStageIntLLRInputS7xD(37)(4) <= CNStageIntLLROutputS7xD(263)(0);
  VNStageIntLLRInputS7xD(88)(4) <= CNStageIntLLROutputS7xD(263)(1);
  VNStageIntLLRInputS7xD(180)(2) <= CNStageIntLLROutputS7xD(263)(2);
  VNStageIntLLRInputS7xD(233)(3) <= CNStageIntLLROutputS7xD(263)(3);
  VNStageIntLLRInputS7xD(304)(4) <= CNStageIntLLROutputS7xD(263)(4);
  VNStageIntLLRInputS7xD(364)(4) <= CNStageIntLLROutputS7xD(263)(5);
  VNStageIntLLRInputS7xD(36)(3) <= CNStageIntLLROutputS7xD(264)(0);
  VNStageIntLLRInputS7xD(115)(4) <= CNStageIntLLROutputS7xD(264)(1);
  VNStageIntLLRInputS7xD(168)(3) <= CNStageIntLLROutputS7xD(264)(2);
  VNStageIntLLRInputS7xD(239)(4) <= CNStageIntLLROutputS7xD(264)(3);
  VNStageIntLLRInputS7xD(299)(3) <= CNStageIntLLROutputS7xD(264)(4);
  VNStageIntLLRInputS7xD(374)(4) <= CNStageIntLLROutputS7xD(264)(5);
  VNStageIntLLRInputS7xD(35)(4) <= CNStageIntLLROutputS7xD(265)(0);
  VNStageIntLLRInputS7xD(103)(4) <= CNStageIntLLROutputS7xD(265)(1);
  VNStageIntLLRInputS7xD(174)(3) <= CNStageIntLLROutputS7xD(265)(2);
  VNStageIntLLRInputS7xD(234)(4) <= CNStageIntLLROutputS7xD(265)(3);
  VNStageIntLLRInputS7xD(309)(4) <= CNStageIntLLROutputS7xD(265)(4);
  VNStageIntLLRInputS7xD(333)(3) <= CNStageIntLLROutputS7xD(265)(5);
  VNStageIntLLRInputS7xD(34)(4) <= CNStageIntLLROutputS7xD(266)(0);
  VNStageIntLLRInputS7xD(109)(4) <= CNStageIntLLROutputS7xD(266)(1);
  VNStageIntLLRInputS7xD(169)(4) <= CNStageIntLLROutputS7xD(266)(2);
  VNStageIntLLRInputS7xD(244)(1) <= CNStageIntLLROutputS7xD(266)(3);
  VNStageIntLLRInputS7xD(268)(4) <= CNStageIntLLROutputS7xD(266)(4);
  VNStageIntLLRInputS7xD(351)(3) <= CNStageIntLLROutputS7xD(266)(5);
  VNStageIntLLRInputS7xD(33)(4) <= CNStageIntLLROutputS7xD(267)(0);
  VNStageIntLLRInputS7xD(104)(4) <= CNStageIntLLROutputS7xD(267)(1);
  VNStageIntLLRInputS7xD(179)(4) <= CNStageIntLLROutputS7xD(267)(2);
  VNStageIntLLRInputS7xD(203)(4) <= CNStageIntLLROutputS7xD(267)(3);
  VNStageIntLLRInputS7xD(286)(4) <= CNStageIntLLROutputS7xD(267)(4);
  VNStageIntLLRInputS7xD(336)(3) <= CNStageIntLLROutputS7xD(267)(5);
  VNStageIntLLRInputS7xD(32)(3) <= CNStageIntLLROutputS7xD(268)(0);
  VNStageIntLLRInputS7xD(114)(4) <= CNStageIntLLROutputS7xD(268)(1);
  VNStageIntLLRInputS7xD(138)(4) <= CNStageIntLLROutputS7xD(268)(2);
  VNStageIntLLRInputS7xD(221)(4) <= CNStageIntLLROutputS7xD(268)(3);
  VNStageIntLLRInputS7xD(271)(3) <= CNStageIntLLROutputS7xD(268)(4);
  VNStageIntLLRInputS7xD(323)(3) <= CNStageIntLLROutputS7xD(268)(5);
  VNStageIntLLRInputS7xD(30)(4) <= CNStageIntLLROutputS7xD(269)(0);
  VNStageIntLLRInputS7xD(91)(4) <= CNStageIntLLROutputS7xD(269)(1);
  VNStageIntLLRInputS7xD(141)(2) <= CNStageIntLLROutputS7xD(269)(2);
  VNStageIntLLRInputS7xD(193)(3) <= CNStageIntLLROutputS7xD(269)(3);
  VNStageIntLLRInputS7xD(289)(4) <= CNStageIntLLROutputS7xD(269)(4);
  VNStageIntLLRInputS7xD(366)(4) <= CNStageIntLLROutputS7xD(269)(5);
  VNStageIntLLRInputS7xD(29)(3) <= CNStageIntLLROutputS7xD(270)(0);
  VNStageIntLLRInputS7xD(76)(4) <= CNStageIntLLROutputS7xD(270)(1);
  VNStageIntLLRInputS7xD(191)(4) <= CNStageIntLLROutputS7xD(270)(2);
  VNStageIntLLRInputS7xD(224)(4) <= CNStageIntLLROutputS7xD(270)(3);
  VNStageIntLLRInputS7xD(301)(4) <= CNStageIntLLROutputS7xD(270)(4);
  VNStageIntLLRInputS7xD(380)(3) <= CNStageIntLLROutputS7xD(270)(5);
  VNStageIntLLRInputS7xD(28)(4) <= CNStageIntLLROutputS7xD(271)(0);
  VNStageIntLLRInputS7xD(126)(3) <= CNStageIntLLROutputS7xD(271)(1);
  VNStageIntLLRInputS7xD(159)(3) <= CNStageIntLLROutputS7xD(271)(2);
  VNStageIntLLRInputS7xD(236)(4) <= CNStageIntLLROutputS7xD(271)(3);
  VNStageIntLLRInputS7xD(315)(3) <= CNStageIntLLROutputS7xD(271)(4);
  VNStageIntLLRInputS7xD(361)(4) <= CNStageIntLLROutputS7xD(271)(5);
  VNStageIntLLRInputS7xD(26)(4) <= CNStageIntLLROutputS7xD(272)(0);
  VNStageIntLLRInputS7xD(106)(3) <= CNStageIntLLROutputS7xD(272)(1);
  VNStageIntLLRInputS7xD(185)(1) <= CNStageIntLLROutputS7xD(272)(2);
  VNStageIntLLRInputS7xD(231)(3) <= CNStageIntLLROutputS7xD(272)(3);
  VNStageIntLLRInputS7xD(273)(3) <= CNStageIntLLROutputS7xD(272)(4);
  VNStageIntLLRInputS7xD(327)(4) <= CNStageIntLLROutputS7xD(272)(5);
  VNStageIntLLRInputS7xD(24)(4) <= CNStageIntLLROutputS7xD(273)(0);
  VNStageIntLLRInputS7xD(101)(4) <= CNStageIntLLROutputS7xD(273)(1);
  VNStageIntLLRInputS7xD(143)(4) <= CNStageIntLLROutputS7xD(273)(2);
  VNStageIntLLRInputS7xD(197)(4) <= CNStageIntLLROutputS7xD(273)(3);
  VNStageIntLLRInputS7xD(266)(3) <= CNStageIntLLROutputS7xD(273)(4);
  VNStageIntLLRInputS7xD(324)(4) <= CNStageIntLLROutputS7xD(273)(5);
  VNStageIntLLRInputS7xD(23)(4) <= CNStageIntLLROutputS7xD(274)(0);
  VNStageIntLLRInputS7xD(78)(4) <= CNStageIntLLROutputS7xD(274)(1);
  VNStageIntLLRInputS7xD(132)(3) <= CNStageIntLLROutputS7xD(274)(2);
  VNStageIntLLRInputS7xD(201)(4) <= CNStageIntLLROutputS7xD(274)(3);
  VNStageIntLLRInputS7xD(259)(2) <= CNStageIntLLROutputS7xD(274)(4);
  VNStageIntLLRInputS7xD(335)(4) <= CNStageIntLLROutputS7xD(274)(5);
  VNStageIntLLRInputS7xD(22)(4) <= CNStageIntLLROutputS7xD(275)(0);
  VNStageIntLLRInputS7xD(67)(1) <= CNStageIntLLROutputS7xD(275)(1);
  VNStageIntLLRInputS7xD(136)(4) <= CNStageIntLLROutputS7xD(275)(2);
  VNStageIntLLRInputS7xD(194)(4) <= CNStageIntLLROutputS7xD(275)(3);
  VNStageIntLLRInputS7xD(270)(4) <= CNStageIntLLROutputS7xD(275)(4);
  VNStageIntLLRInputS7xD(370)(3) <= CNStageIntLLROutputS7xD(275)(5);
  VNStageIntLLRInputS7xD(21)(4) <= CNStageIntLLROutputS7xD(276)(0);
  VNStageIntLLRInputS7xD(71)(3) <= CNStageIntLLROutputS7xD(276)(1);
  VNStageIntLLRInputS7xD(129)(4) <= CNStageIntLLROutputS7xD(276)(2);
  VNStageIntLLRInputS7xD(205)(1) <= CNStageIntLLROutputS7xD(276)(3);
  VNStageIntLLRInputS7xD(305)(4) <= CNStageIntLLROutputS7xD(276)(4);
  VNStageIntLLRInputS7xD(362)(4) <= CNStageIntLLROutputS7xD(276)(5);
  VNStageIntLLRInputS7xD(20)(2) <= CNStageIntLLROutputS7xD(277)(0);
  VNStageIntLLRInputS7xD(127)(4) <= CNStageIntLLROutputS7xD(277)(1);
  VNStageIntLLRInputS7xD(140)(4) <= CNStageIntLLROutputS7xD(277)(2);
  VNStageIntLLRInputS7xD(240)(4) <= CNStageIntLLROutputS7xD(277)(3);
  VNStageIntLLRInputS7xD(297)(4) <= CNStageIntLLROutputS7xD(277)(4);
  VNStageIntLLRInputS7xD(379)(2) <= CNStageIntLLROutputS7xD(277)(5);
  VNStageIntLLRInputS7xD(19)(3) <= CNStageIntLLROutputS7xD(278)(0);
  VNStageIntLLRInputS7xD(75)(4) <= CNStageIntLLROutputS7xD(278)(1);
  VNStageIntLLRInputS7xD(175)(4) <= CNStageIntLLROutputS7xD(278)(2);
  VNStageIntLLRInputS7xD(232)(3) <= CNStageIntLLROutputS7xD(278)(3);
  VNStageIntLLRInputS7xD(314)(1) <= CNStageIntLLROutputS7xD(278)(4);
  VNStageIntLLRInputS7xD(376)(3) <= CNStageIntLLROutputS7xD(278)(5);
  VNStageIntLLRInputS7xD(0)(4) <= CNStageIntLLROutputS7xD(279)(0);
  VNStageIntLLRInputS7xD(123)(3) <= CNStageIntLLROutputS7xD(279)(1);
  VNStageIntLLRInputS7xD(188)(2) <= CNStageIntLLROutputS7xD(279)(2);
  VNStageIntLLRInputS7xD(253)(3) <= CNStageIntLLROutputS7xD(279)(3);
  VNStageIntLLRInputS7xD(318)(2) <= CNStageIntLLROutputS7xD(279)(4);
  VNStageIntLLRInputS7xD(383)(4) <= CNStageIntLLROutputS7xD(279)(5);
  VNStageIntLLRInputS7xD(35)(5) <= CNStageIntLLROutputS7xD(280)(0);
  VNStageIntLLRInputS7xD(91)(5) <= CNStageIntLLROutputS7xD(280)(1);
  VNStageIntLLRInputS7xD(191)(5) <= CNStageIntLLROutputS7xD(280)(2);
  VNStageIntLLRInputS7xD(248)(5) <= CNStageIntLLROutputS7xD(280)(3);
  VNStageIntLLRInputS7xD(267)(5) <= CNStageIntLLROutputS7xD(280)(4);
  VNStageIntLLRInputS7xD(329)(5) <= CNStageIntLLROutputS7xD(280)(5);
  VNStageIntLLRInputS7xD(34)(5) <= CNStageIntLLROutputS7xD(281)(0);
  VNStageIntLLRInputS7xD(126)(4) <= CNStageIntLLROutputS7xD(281)(1);
  VNStageIntLLRInputS7xD(183)(3) <= CNStageIntLLROutputS7xD(281)(2);
  VNStageIntLLRInputS7xD(202)(4) <= CNStageIntLLROutputS7xD(281)(3);
  VNStageIntLLRInputS7xD(264)(5) <= CNStageIntLLROutputS7xD(281)(4);
  VNStageIntLLRInputS7xD(363)(4) <= CNStageIntLLROutputS7xD(281)(5);
  VNStageIntLLRInputS7xD(33)(5) <= CNStageIntLLROutputS7xD(282)(0);
  VNStageIntLLRInputS7xD(118)(4) <= CNStageIntLLROutputS7xD(282)(1);
  VNStageIntLLRInputS7xD(137)(5) <= CNStageIntLLROutputS7xD(282)(2);
  VNStageIntLLRInputS7xD(199)(5) <= CNStageIntLLROutputS7xD(282)(3);
  VNStageIntLLRInputS7xD(298)(5) <= CNStageIntLLROutputS7xD(282)(4);
  VNStageIntLLRInputS7xD(383)(5) <= CNStageIntLLROutputS7xD(282)(5);
  VNStageIntLLRInputS7xD(31)(3) <= CNStageIntLLROutputS7xD(283)(0);
  VNStageIntLLRInputS7xD(69)(5) <= CNStageIntLLROutputS7xD(283)(1);
  VNStageIntLLRInputS7xD(168)(4) <= CNStageIntLLROutputS7xD(283)(2);
  VNStageIntLLRInputS7xD(253)(4) <= CNStageIntLLROutputS7xD(283)(3);
  VNStageIntLLRInputS7xD(304)(5) <= CNStageIntLLROutputS7xD(283)(4);
  VNStageIntLLRInputS7xD(359)(5) <= CNStageIntLLROutputS7xD(283)(5);
  VNStageIntLLRInputS7xD(30)(5) <= CNStageIntLLROutputS7xD(284)(0);
  VNStageIntLLRInputS7xD(103)(5) <= CNStageIntLLROutputS7xD(284)(1);
  VNStageIntLLRInputS7xD(188)(3) <= CNStageIntLLROutputS7xD(284)(2);
  VNStageIntLLRInputS7xD(239)(5) <= CNStageIntLLROutputS7xD(284)(3);
  VNStageIntLLRInputS7xD(294)(5) <= CNStageIntLLROutputS7xD(284)(4);
  VNStageIntLLRInputS7xD(325)(5) <= CNStageIntLLROutputS7xD(284)(5);
  VNStageIntLLRInputS7xD(27)(4) <= CNStageIntLLROutputS7xD(285)(0);
  VNStageIntLLRInputS7xD(99)(5) <= CNStageIntLLROutputS7xD(285)(1);
  VNStageIntLLRInputS7xD(130)(5) <= CNStageIntLLROutputS7xD(285)(2);
  VNStageIntLLRInputS7xD(241)(4) <= CNStageIntLLROutputS7xD(285)(3);
  VNStageIntLLRInputS7xD(273)(4) <= CNStageIntLLROutputS7xD(285)(4);
  VNStageIntLLRInputS7xD(361)(5) <= CNStageIntLLROutputS7xD(285)(5);
  VNStageIntLLRInputS7xD(26)(5) <= CNStageIntLLROutputS7xD(286)(0);
  VNStageIntLLRInputS7xD(65)(4) <= CNStageIntLLROutputS7xD(286)(1);
  VNStageIntLLRInputS7xD(176)(5) <= CNStageIntLLROutputS7xD(286)(2);
  VNStageIntLLRInputS7xD(208)(4) <= CNStageIntLLROutputS7xD(286)(3);
  VNStageIntLLRInputS7xD(296)(4) <= CNStageIntLLROutputS7xD(286)(4);
  VNStageIntLLRInputS7xD(334)(3) <= CNStageIntLLROutputS7xD(286)(5);
  VNStageIntLLRInputS7xD(25)(4) <= CNStageIntLLROutputS7xD(287)(0);
  VNStageIntLLRInputS7xD(111)(5) <= CNStageIntLLROutputS7xD(287)(1);
  VNStageIntLLRInputS7xD(143)(5) <= CNStageIntLLROutputS7xD(287)(2);
  VNStageIntLLRInputS7xD(231)(4) <= CNStageIntLLROutputS7xD(287)(3);
  VNStageIntLLRInputS7xD(269)(4) <= CNStageIntLLROutputS7xD(287)(4);
  VNStageIntLLRInputS7xD(381)(4) <= CNStageIntLLROutputS7xD(287)(5);
  VNStageIntLLRInputS7xD(24)(5) <= CNStageIntLLROutputS7xD(288)(0);
  VNStageIntLLRInputS7xD(78)(5) <= CNStageIntLLROutputS7xD(288)(1);
  VNStageIntLLRInputS7xD(166)(4) <= CNStageIntLLROutputS7xD(288)(2);
  VNStageIntLLRInputS7xD(204)(5) <= CNStageIntLLROutputS7xD(288)(3);
  VNStageIntLLRInputS7xD(316)(3) <= CNStageIntLLROutputS7xD(288)(4);
  VNStageIntLLRInputS7xD(321)(5) <= CNStageIntLLROutputS7xD(288)(5);
  VNStageIntLLRInputS7xD(23)(5) <= CNStageIntLLROutputS7xD(289)(0);
  VNStageIntLLRInputS7xD(101)(5) <= CNStageIntLLROutputS7xD(289)(1);
  VNStageIntLLRInputS7xD(139)(5) <= CNStageIntLLROutputS7xD(289)(2);
  VNStageIntLLRInputS7xD(251)(3) <= CNStageIntLLROutputS7xD(289)(3);
  VNStageIntLLRInputS7xD(319)(5) <= CNStageIntLLROutputS7xD(289)(4);
  VNStageIntLLRInputS7xD(362)(5) <= CNStageIntLLROutputS7xD(289)(5);
  VNStageIntLLRInputS7xD(22)(5) <= CNStageIntLLROutputS7xD(290)(0);
  VNStageIntLLRInputS7xD(74)(4) <= CNStageIntLLROutputS7xD(290)(1);
  VNStageIntLLRInputS7xD(186)(4) <= CNStageIntLLROutputS7xD(290)(2);
  VNStageIntLLRInputS7xD(254)(3) <= CNStageIntLLROutputS7xD(290)(3);
  VNStageIntLLRInputS7xD(297)(5) <= CNStageIntLLROutputS7xD(290)(4);
  VNStageIntLLRInputS7xD(337)(5) <= CNStageIntLLROutputS7xD(290)(5);
  VNStageIntLLRInputS7xD(21)(5) <= CNStageIntLLROutputS7xD(291)(0);
  VNStageIntLLRInputS7xD(121)(4) <= CNStageIntLLROutputS7xD(291)(1);
  VNStageIntLLRInputS7xD(189)(4) <= CNStageIntLLROutputS7xD(291)(2);
  VNStageIntLLRInputS7xD(232)(4) <= CNStageIntLLROutputS7xD(291)(3);
  VNStageIntLLRInputS7xD(272)(5) <= CNStageIntLLROutputS7xD(291)(4);
  VNStageIntLLRInputS7xD(335)(5) <= CNStageIntLLROutputS7xD(291)(5);
  VNStageIntLLRInputS7xD(20)(3) <= CNStageIntLLROutputS7xD(292)(0);
  VNStageIntLLRInputS7xD(124)(3) <= CNStageIntLLROutputS7xD(292)(1);
  VNStageIntLLRInputS7xD(167)(5) <= CNStageIntLLROutputS7xD(292)(2);
  VNStageIntLLRInputS7xD(207)(4) <= CNStageIntLLROutputS7xD(292)(3);
  VNStageIntLLRInputS7xD(270)(5) <= CNStageIntLLROutputS7xD(292)(4);
  VNStageIntLLRInputS7xD(360)(5) <= CNStageIntLLROutputS7xD(292)(5);
  VNStageIntLLRInputS7xD(18)(5) <= CNStageIntLLROutputS7xD(293)(0);
  VNStageIntLLRInputS7xD(77)(3) <= CNStageIntLLROutputS7xD(293)(1);
  VNStageIntLLRInputS7xD(140)(5) <= CNStageIntLLROutputS7xD(293)(2);
  VNStageIntLLRInputS7xD(230)(4) <= CNStageIntLLROutputS7xD(293)(3);
  VNStageIntLLRInputS7xD(303)(5) <= CNStageIntLLROutputS7xD(293)(4);
  VNStageIntLLRInputS7xD(348)(5) <= CNStageIntLLROutputS7xD(293)(5);
  VNStageIntLLRInputS7xD(17)(5) <= CNStageIntLLROutputS7xD(294)(0);
  VNStageIntLLRInputS7xD(75)(5) <= CNStageIntLLROutputS7xD(294)(1);
  VNStageIntLLRInputS7xD(165)(4) <= CNStageIntLLROutputS7xD(294)(2);
  VNStageIntLLRInputS7xD(238)(5) <= CNStageIntLLROutputS7xD(294)(3);
  VNStageIntLLRInputS7xD(283)(5) <= CNStageIntLLROutputS7xD(294)(4);
  VNStageIntLLRInputS7xD(342)(4) <= CNStageIntLLROutputS7xD(294)(5);
  VNStageIntLLRInputS7xD(16)(4) <= CNStageIntLLROutputS7xD(295)(0);
  VNStageIntLLRInputS7xD(100)(5) <= CNStageIntLLROutputS7xD(295)(1);
  VNStageIntLLRInputS7xD(173)(5) <= CNStageIntLLROutputS7xD(295)(2);
  VNStageIntLLRInputS7xD(218)(5) <= CNStageIntLLROutputS7xD(295)(3);
  VNStageIntLLRInputS7xD(277)(5) <= CNStageIntLLROutputS7xD(295)(4);
  VNStageIntLLRInputS7xD(320)(3) <= CNStageIntLLROutputS7xD(295)(5);
  VNStageIntLLRInputS7xD(15)(5) <= CNStageIntLLROutputS7xD(296)(0);
  VNStageIntLLRInputS7xD(108)(5) <= CNStageIntLLROutputS7xD(296)(1);
  VNStageIntLLRInputS7xD(153)(5) <= CNStageIntLLROutputS7xD(296)(2);
  VNStageIntLLRInputS7xD(212)(4) <= CNStageIntLLROutputS7xD(296)(3);
  VNStageIntLLRInputS7xD(256)(4) <= CNStageIntLLROutputS7xD(296)(4);
  VNStageIntLLRInputS7xD(341)(5) <= CNStageIntLLROutputS7xD(296)(5);
  VNStageIntLLRInputS7xD(14)(5) <= CNStageIntLLROutputS7xD(297)(0);
  VNStageIntLLRInputS7xD(88)(5) <= CNStageIntLLROutputS7xD(297)(1);
  VNStageIntLLRInputS7xD(147)(5) <= CNStageIntLLROutputS7xD(297)(2);
  VNStageIntLLRInputS7xD(192)(5) <= CNStageIntLLROutputS7xD(297)(3);
  VNStageIntLLRInputS7xD(276)(5) <= CNStageIntLLROutputS7xD(297)(4);
  VNStageIntLLRInputS7xD(346)(5) <= CNStageIntLLROutputS7xD(297)(5);
  VNStageIntLLRInputS7xD(13)(4) <= CNStageIntLLROutputS7xD(298)(0);
  VNStageIntLLRInputS7xD(82)(5) <= CNStageIntLLROutputS7xD(298)(1);
  VNStageIntLLRInputS7xD(128)(5) <= CNStageIntLLROutputS7xD(298)(2);
  VNStageIntLLRInputS7xD(211)(5) <= CNStageIntLLROutputS7xD(298)(3);
  VNStageIntLLRInputS7xD(281)(5) <= CNStageIntLLROutputS7xD(298)(4);
  VNStageIntLLRInputS7xD(365)(5) <= CNStageIntLLROutputS7xD(298)(5);
  VNStageIntLLRInputS7xD(12)(5) <= CNStageIntLLROutputS7xD(299)(0);
  VNStageIntLLRInputS7xD(64)(4) <= CNStageIntLLROutputS7xD(299)(1);
  VNStageIntLLRInputS7xD(146)(4) <= CNStageIntLLROutputS7xD(299)(2);
  VNStageIntLLRInputS7xD(216)(5) <= CNStageIntLLROutputS7xD(299)(3);
  VNStageIntLLRInputS7xD(300)(4) <= CNStageIntLLROutputS7xD(299)(4);
  VNStageIntLLRInputS7xD(356)(4) <= CNStageIntLLROutputS7xD(299)(5);
  VNStageIntLLRInputS7xD(9)(5) <= CNStageIntLLROutputS7xD(300)(0);
  VNStageIntLLRInputS7xD(105)(4) <= CNStageIntLLROutputS7xD(300)(1);
  VNStageIntLLRInputS7xD(161)(5) <= CNStageIntLLROutputS7xD(300)(2);
  VNStageIntLLRInputS7xD(200)(5) <= CNStageIntLLROutputS7xD(300)(3);
  VNStageIntLLRInputS7xD(266)(4) <= CNStageIntLLROutputS7xD(300)(4);
  VNStageIntLLRInputS7xD(355)(5) <= CNStageIntLLROutputS7xD(300)(5);
  VNStageIntLLRInputS7xD(7)(5) <= CNStageIntLLROutputS7xD(301)(0);
  VNStageIntLLRInputS7xD(70)(5) <= CNStageIntLLROutputS7xD(301)(1);
  VNStageIntLLRInputS7xD(136)(5) <= CNStageIntLLROutputS7xD(301)(2);
  VNStageIntLLRInputS7xD(225)(5) <= CNStageIntLLROutputS7xD(301)(3);
  VNStageIntLLRInputS7xD(311)(4) <= CNStageIntLLROutputS7xD(301)(4);
  VNStageIntLLRInputS7xD(372)(4) <= CNStageIntLLROutputS7xD(301)(5);
  VNStageIntLLRInputS7xD(6)(5) <= CNStageIntLLROutputS7xD(302)(0);
  VNStageIntLLRInputS7xD(71)(4) <= CNStageIntLLROutputS7xD(302)(1);
  VNStageIntLLRInputS7xD(160)(5) <= CNStageIntLLROutputS7xD(302)(2);
  VNStageIntLLRInputS7xD(246)(5) <= CNStageIntLLROutputS7xD(302)(3);
  VNStageIntLLRInputS7xD(307)(5) <= CNStageIntLLROutputS7xD(302)(4);
  VNStageIntLLRInputS7xD(324)(5) <= CNStageIntLLROutputS7xD(302)(5);
  VNStageIntLLRInputS7xD(5)(5) <= CNStageIntLLROutputS7xD(303)(0);
  VNStageIntLLRInputS7xD(95)(5) <= CNStageIntLLROutputS7xD(303)(1);
  VNStageIntLLRInputS7xD(181)(5) <= CNStageIntLLROutputS7xD(303)(2);
  VNStageIntLLRInputS7xD(242)(5) <= CNStageIntLLROutputS7xD(303)(3);
  VNStageIntLLRInputS7xD(259)(3) <= CNStageIntLLROutputS7xD(303)(4);
  VNStageIntLLRInputS7xD(350)(5) <= CNStageIntLLROutputS7xD(303)(5);
  VNStageIntLLRInputS7xD(4)(4) <= CNStageIntLLROutputS7xD(304)(0);
  VNStageIntLLRInputS7xD(116)(4) <= CNStageIntLLROutputS7xD(304)(1);
  VNStageIntLLRInputS7xD(177)(5) <= CNStageIntLLROutputS7xD(304)(2);
  VNStageIntLLRInputS7xD(194)(5) <= CNStageIntLLROutputS7xD(304)(3);
  VNStageIntLLRInputS7xD(285)(5) <= CNStageIntLLROutputS7xD(304)(4);
  VNStageIntLLRInputS7xD(326)(4) <= CNStageIntLLROutputS7xD(304)(5);
  VNStageIntLLRInputS7xD(3)(4) <= CNStageIntLLROutputS7xD(305)(0);
  VNStageIntLLRInputS7xD(112)(5) <= CNStageIntLLROutputS7xD(305)(1);
  VNStageIntLLRInputS7xD(129)(5) <= CNStageIntLLROutputS7xD(305)(2);
  VNStageIntLLRInputS7xD(220)(5) <= CNStageIntLLROutputS7xD(305)(3);
  VNStageIntLLRInputS7xD(261)(4) <= CNStageIntLLROutputS7xD(305)(4);
  VNStageIntLLRInputS7xD(358)(4) <= CNStageIntLLROutputS7xD(305)(5);
  VNStageIntLLRInputS7xD(2)(5) <= CNStageIntLLROutputS7xD(306)(0);
  VNStageIntLLRInputS7xD(127)(5) <= CNStageIntLLROutputS7xD(306)(1);
  VNStageIntLLRInputS7xD(155)(5) <= CNStageIntLLROutputS7xD(306)(2);
  VNStageIntLLRInputS7xD(196)(5) <= CNStageIntLLROutputS7xD(306)(3);
  VNStageIntLLRInputS7xD(293)(4) <= CNStageIntLLROutputS7xD(306)(4);
  VNStageIntLLRInputS7xD(374)(5) <= CNStageIntLLROutputS7xD(306)(5);
  VNStageIntLLRInputS7xD(1)(4) <= CNStageIntLLROutputS7xD(307)(0);
  VNStageIntLLRInputS7xD(90)(5) <= CNStageIntLLROutputS7xD(307)(1);
  VNStageIntLLRInputS7xD(131)(4) <= CNStageIntLLROutputS7xD(307)(2);
  VNStageIntLLRInputS7xD(228)(5) <= CNStageIntLLROutputS7xD(307)(3);
  VNStageIntLLRInputS7xD(309)(5) <= CNStageIntLLROutputS7xD(307)(4);
  VNStageIntLLRInputS7xD(344)(5) <= CNStageIntLLROutputS7xD(307)(5);
  VNStageIntLLRInputS7xD(62)(4) <= CNStageIntLLROutputS7xD(308)(0);
  VNStageIntLLRInputS7xD(98)(4) <= CNStageIntLLROutputS7xD(308)(1);
  VNStageIntLLRInputS7xD(179)(5) <= CNStageIntLLROutputS7xD(308)(2);
  VNStageIntLLRInputS7xD(214)(5) <= CNStageIntLLROutputS7xD(308)(3);
  VNStageIntLLRInputS7xD(288)(5) <= CNStageIntLLROutputS7xD(308)(4);
  VNStageIntLLRInputS7xD(366)(5) <= CNStageIntLLROutputS7xD(308)(5);
  VNStageIntLLRInputS7xD(61)(4) <= CNStageIntLLROutputS7xD(309)(0);
  VNStageIntLLRInputS7xD(114)(5) <= CNStageIntLLROutputS7xD(309)(1);
  VNStageIntLLRInputS7xD(149)(5) <= CNStageIntLLROutputS7xD(309)(2);
  VNStageIntLLRInputS7xD(223)(5) <= CNStageIntLLROutputS7xD(309)(3);
  VNStageIntLLRInputS7xD(301)(5) <= CNStageIntLLROutputS7xD(309)(4);
  VNStageIntLLRInputS7xD(345)(4) <= CNStageIntLLROutputS7xD(309)(5);
  VNStageIntLLRInputS7xD(60)(4) <= CNStageIntLLROutputS7xD(310)(0);
  VNStageIntLLRInputS7xD(84)(4) <= CNStageIntLLROutputS7xD(310)(1);
  VNStageIntLLRInputS7xD(158)(5) <= CNStageIntLLROutputS7xD(310)(2);
  VNStageIntLLRInputS7xD(236)(5) <= CNStageIntLLROutputS7xD(310)(3);
  VNStageIntLLRInputS7xD(280)(5) <= CNStageIntLLROutputS7xD(310)(4);
  VNStageIntLLRInputS7xD(373)(3) <= CNStageIntLLROutputS7xD(310)(5);
  VNStageIntLLRInputS7xD(59)(3) <= CNStageIntLLROutputS7xD(311)(0);
  VNStageIntLLRInputS7xD(93)(5) <= CNStageIntLLROutputS7xD(311)(1);
  VNStageIntLLRInputS7xD(171)(3) <= CNStageIntLLROutputS7xD(311)(2);
  VNStageIntLLRInputS7xD(215)(5) <= CNStageIntLLROutputS7xD(311)(3);
  VNStageIntLLRInputS7xD(308)(3) <= CNStageIntLLROutputS7xD(311)(4);
  VNStageIntLLRInputS7xD(375)(4) <= CNStageIntLLROutputS7xD(311)(5);
  VNStageIntLLRInputS7xD(58)(3) <= CNStageIntLLROutputS7xD(312)(0);
  VNStageIntLLRInputS7xD(106)(4) <= CNStageIntLLROutputS7xD(312)(1);
  VNStageIntLLRInputS7xD(150)(4) <= CNStageIntLLROutputS7xD(312)(2);
  VNStageIntLLRInputS7xD(243)(5) <= CNStageIntLLROutputS7xD(312)(3);
  VNStageIntLLRInputS7xD(310)(4) <= CNStageIntLLROutputS7xD(312)(4);
  VNStageIntLLRInputS7xD(357)(5) <= CNStageIntLLROutputS7xD(312)(5);
  VNStageIntLLRInputS7xD(57)(4) <= CNStageIntLLROutputS7xD(313)(0);
  VNStageIntLLRInputS7xD(85)(4) <= CNStageIntLLROutputS7xD(313)(1);
  VNStageIntLLRInputS7xD(178)(4) <= CNStageIntLLROutputS7xD(313)(2);
  VNStageIntLLRInputS7xD(245)(5) <= CNStageIntLLROutputS7xD(313)(3);
  VNStageIntLLRInputS7xD(292)(5) <= CNStageIntLLROutputS7xD(313)(4);
  VNStageIntLLRInputS7xD(364)(5) <= CNStageIntLLROutputS7xD(313)(5);
  VNStageIntLLRInputS7xD(56)(5) <= CNStageIntLLROutputS7xD(314)(0);
  VNStageIntLLRInputS7xD(113)(5) <= CNStageIntLLROutputS7xD(314)(1);
  VNStageIntLLRInputS7xD(180)(3) <= CNStageIntLLROutputS7xD(314)(2);
  VNStageIntLLRInputS7xD(227)(5) <= CNStageIntLLROutputS7xD(314)(3);
  VNStageIntLLRInputS7xD(299)(4) <= CNStageIntLLROutputS7xD(314)(4);
  VNStageIntLLRInputS7xD(328)(3) <= CNStageIntLLROutputS7xD(314)(5);
  VNStageIntLLRInputS7xD(55)(5) <= CNStageIntLLROutputS7xD(315)(0);
  VNStageIntLLRInputS7xD(115)(5) <= CNStageIntLLROutputS7xD(315)(1);
  VNStageIntLLRInputS7xD(162)(5) <= CNStageIntLLROutputS7xD(315)(2);
  VNStageIntLLRInputS7xD(234)(5) <= CNStageIntLLROutputS7xD(315)(3);
  VNStageIntLLRInputS7xD(263)(5) <= CNStageIntLLROutputS7xD(315)(4);
  VNStageIntLLRInputS7xD(379)(3) <= CNStageIntLLROutputS7xD(315)(5);
  VNStageIntLLRInputS7xD(54)(4) <= CNStageIntLLROutputS7xD(316)(0);
  VNStageIntLLRInputS7xD(97)(5) <= CNStageIntLLROutputS7xD(316)(1);
  VNStageIntLLRInputS7xD(169)(5) <= CNStageIntLLROutputS7xD(316)(2);
  VNStageIntLLRInputS7xD(198)(5) <= CNStageIntLLROutputS7xD(316)(3);
  VNStageIntLLRInputS7xD(314)(2) <= CNStageIntLLROutputS7xD(316)(4);
  VNStageIntLLRInputS7xD(322)(4) <= CNStageIntLLROutputS7xD(316)(5);
  VNStageIntLLRInputS7xD(53)(4) <= CNStageIntLLROutputS7xD(317)(0);
  VNStageIntLLRInputS7xD(104)(5) <= CNStageIntLLROutputS7xD(317)(1);
  VNStageIntLLRInputS7xD(133)(3) <= CNStageIntLLROutputS7xD(317)(2);
  VNStageIntLLRInputS7xD(249)(3) <= CNStageIntLLROutputS7xD(317)(3);
  VNStageIntLLRInputS7xD(257)(5) <= CNStageIntLLROutputS7xD(317)(4);
  VNStageIntLLRInputS7xD(380)(4) <= CNStageIntLLROutputS7xD(317)(5);
  VNStageIntLLRInputS7xD(52)(3) <= CNStageIntLLROutputS7xD(318)(0);
  VNStageIntLLRInputS7xD(68)(4) <= CNStageIntLLROutputS7xD(318)(1);
  VNStageIntLLRInputS7xD(184)(5) <= CNStageIntLLROutputS7xD(318)(2);
  VNStageIntLLRInputS7xD(255)(5) <= CNStageIntLLROutputS7xD(318)(3);
  VNStageIntLLRInputS7xD(315)(4) <= CNStageIntLLROutputS7xD(318)(4);
  VNStageIntLLRInputS7xD(327)(5) <= CNStageIntLLROutputS7xD(318)(5);
  VNStageIntLLRInputS7xD(51)(4) <= CNStageIntLLROutputS7xD(319)(0);
  VNStageIntLLRInputS7xD(119)(4) <= CNStageIntLLROutputS7xD(319)(1);
  VNStageIntLLRInputS7xD(190)(3) <= CNStageIntLLROutputS7xD(319)(2);
  VNStageIntLLRInputS7xD(250)(3) <= CNStageIntLLROutputS7xD(319)(3);
  VNStageIntLLRInputS7xD(262)(4) <= CNStageIntLLROutputS7xD(319)(4);
  VNStageIntLLRInputS7xD(349)(4) <= CNStageIntLLROutputS7xD(319)(5);
  VNStageIntLLRInputS7xD(50)(5) <= CNStageIntLLROutputS7xD(320)(0);
  VNStageIntLLRInputS7xD(125)(2) <= CNStageIntLLROutputS7xD(320)(1);
  VNStageIntLLRInputS7xD(185)(2) <= CNStageIntLLROutputS7xD(320)(2);
  VNStageIntLLRInputS7xD(197)(5) <= CNStageIntLLROutputS7xD(320)(3);
  VNStageIntLLRInputS7xD(284)(5) <= CNStageIntLLROutputS7xD(320)(4);
  VNStageIntLLRInputS7xD(367)(5) <= CNStageIntLLROutputS7xD(320)(5);
  VNStageIntLLRInputS7xD(49)(5) <= CNStageIntLLROutputS7xD(321)(0);
  VNStageIntLLRInputS7xD(120)(2) <= CNStageIntLLROutputS7xD(321)(1);
  VNStageIntLLRInputS7xD(132)(4) <= CNStageIntLLROutputS7xD(321)(2);
  VNStageIntLLRInputS7xD(219)(4) <= CNStageIntLLROutputS7xD(321)(3);
  VNStageIntLLRInputS7xD(302)(5) <= CNStageIntLLROutputS7xD(321)(4);
  VNStageIntLLRInputS7xD(352)(5) <= CNStageIntLLROutputS7xD(321)(5);
  VNStageIntLLRInputS7xD(48)(2) <= CNStageIntLLROutputS7xD(322)(0);
  VNStageIntLLRInputS7xD(67)(2) <= CNStageIntLLROutputS7xD(322)(1);
  VNStageIntLLRInputS7xD(154)(4) <= CNStageIntLLROutputS7xD(322)(2);
  VNStageIntLLRInputS7xD(237)(4) <= CNStageIntLLROutputS7xD(322)(3);
  VNStageIntLLRInputS7xD(287)(5) <= CNStageIntLLROutputS7xD(322)(4);
  VNStageIntLLRInputS7xD(339)(5) <= CNStageIntLLROutputS7xD(322)(5);
  VNStageIntLLRInputS7xD(46)(5) <= CNStageIntLLROutputS7xD(323)(0);
  VNStageIntLLRInputS7xD(107)(4) <= CNStageIntLLROutputS7xD(323)(1);
  VNStageIntLLRInputS7xD(157)(4) <= CNStageIntLLROutputS7xD(323)(2);
  VNStageIntLLRInputS7xD(209)(4) <= CNStageIntLLROutputS7xD(323)(3);
  VNStageIntLLRInputS7xD(305)(5) <= CNStageIntLLROutputS7xD(323)(4);
  VNStageIntLLRInputS7xD(382)(4) <= CNStageIntLLROutputS7xD(323)(5);
  VNStageIntLLRInputS7xD(45)(5) <= CNStageIntLLROutputS7xD(324)(0);
  VNStageIntLLRInputS7xD(92)(5) <= CNStageIntLLROutputS7xD(324)(1);
  VNStageIntLLRInputS7xD(144)(5) <= CNStageIntLLROutputS7xD(324)(2);
  VNStageIntLLRInputS7xD(240)(5) <= CNStageIntLLROutputS7xD(324)(3);
  VNStageIntLLRInputS7xD(317)(2) <= CNStageIntLLROutputS7xD(324)(4);
  VNStageIntLLRInputS7xD(333)(4) <= CNStageIntLLROutputS7xD(324)(5);
  VNStageIntLLRInputS7xD(44)(5) <= CNStageIntLLROutputS7xD(325)(0);
  VNStageIntLLRInputS7xD(79)(4) <= CNStageIntLLROutputS7xD(325)(1);
  VNStageIntLLRInputS7xD(175)(5) <= CNStageIntLLROutputS7xD(325)(2);
  VNStageIntLLRInputS7xD(252)(4) <= CNStageIntLLROutputS7xD(325)(3);
  VNStageIntLLRInputS7xD(268)(5) <= CNStageIntLLROutputS7xD(325)(4);
  VNStageIntLLRInputS7xD(377)(3) <= CNStageIntLLROutputS7xD(325)(5);
  VNStageIntLLRInputS7xD(43)(4) <= CNStageIntLLROutputS7xD(326)(0);
  VNStageIntLLRInputS7xD(110)(5) <= CNStageIntLLROutputS7xD(326)(1);
  VNStageIntLLRInputS7xD(187)(4) <= CNStageIntLLROutputS7xD(326)(2);
  VNStageIntLLRInputS7xD(203)(5) <= CNStageIntLLROutputS7xD(326)(3);
  VNStageIntLLRInputS7xD(312)(4) <= CNStageIntLLROutputS7xD(326)(4);
  VNStageIntLLRInputS7xD(354)(4) <= CNStageIntLLROutputS7xD(326)(5);
  VNStageIntLLRInputS7xD(42)(5) <= CNStageIntLLROutputS7xD(327)(0);
  VNStageIntLLRInputS7xD(122)(4) <= CNStageIntLLROutputS7xD(327)(1);
  VNStageIntLLRInputS7xD(138)(5) <= CNStageIntLLROutputS7xD(327)(2);
  VNStageIntLLRInputS7xD(247)(5) <= CNStageIntLLROutputS7xD(327)(3);
  VNStageIntLLRInputS7xD(289)(5) <= CNStageIntLLROutputS7xD(327)(4);
  VNStageIntLLRInputS7xD(343)(5) <= CNStageIntLLROutputS7xD(327)(5);
  VNStageIntLLRInputS7xD(41)(5) <= CNStageIntLLROutputS7xD(328)(0);
  VNStageIntLLRInputS7xD(73)(4) <= CNStageIntLLROutputS7xD(328)(1);
  VNStageIntLLRInputS7xD(182)(5) <= CNStageIntLLROutputS7xD(328)(2);
  VNStageIntLLRInputS7xD(224)(5) <= CNStageIntLLROutputS7xD(328)(3);
  VNStageIntLLRInputS7xD(278)(4) <= CNStageIntLLROutputS7xD(328)(4);
  VNStageIntLLRInputS7xD(347)(5) <= CNStageIntLLROutputS7xD(328)(5);
  VNStageIntLLRInputS7xD(39)(5) <= CNStageIntLLROutputS7xD(329)(0);
  VNStageIntLLRInputS7xD(94)(3) <= CNStageIntLLROutputS7xD(329)(1);
  VNStageIntLLRInputS7xD(148)(5) <= CNStageIntLLROutputS7xD(329)(2);
  VNStageIntLLRInputS7xD(217)(5) <= CNStageIntLLROutputS7xD(329)(3);
  VNStageIntLLRInputS7xD(275)(4) <= CNStageIntLLROutputS7xD(329)(4);
  VNStageIntLLRInputS7xD(351)(4) <= CNStageIntLLROutputS7xD(329)(5);
  VNStageIntLLRInputS7xD(38)(5) <= CNStageIntLLROutputS7xD(330)(0);
  VNStageIntLLRInputS7xD(83)(5) <= CNStageIntLLROutputS7xD(330)(1);
  VNStageIntLLRInputS7xD(152)(5) <= CNStageIntLLROutputS7xD(330)(2);
  VNStageIntLLRInputS7xD(210)(5) <= CNStageIntLLROutputS7xD(330)(3);
  VNStageIntLLRInputS7xD(286)(5) <= CNStageIntLLROutputS7xD(330)(4);
  VNStageIntLLRInputS7xD(323)(4) <= CNStageIntLLROutputS7xD(330)(5);
  VNStageIntLLRInputS7xD(37)(5) <= CNStageIntLLROutputS7xD(331)(0);
  VNStageIntLLRInputS7xD(87)(5) <= CNStageIntLLROutputS7xD(331)(1);
  VNStageIntLLRInputS7xD(145)(5) <= CNStageIntLLROutputS7xD(331)(2);
  VNStageIntLLRInputS7xD(221)(5) <= CNStageIntLLROutputS7xD(331)(3);
  VNStageIntLLRInputS7xD(258)(2) <= CNStageIntLLROutputS7xD(331)(4);
  VNStageIntLLRInputS7xD(378)(4) <= CNStageIntLLROutputS7xD(331)(5);
  VNStageIntLLRInputS7xD(0)(5) <= CNStageIntLLROutputS7xD(332)(0);
  VNStageIntLLRInputS7xD(76)(5) <= CNStageIntLLROutputS7xD(332)(1);
  VNStageIntLLRInputS7xD(141)(3) <= CNStageIntLLROutputS7xD(332)(2);
  VNStageIntLLRInputS7xD(206)(3) <= CNStageIntLLROutputS7xD(332)(3);
  VNStageIntLLRInputS7xD(271)(4) <= CNStageIntLLROutputS7xD(332)(4);
  VNStageIntLLRInputS7xD(336)(4) <= CNStageIntLLROutputS7xD(332)(5);
  VNStageIntLLRInputS7xD(28)(5) <= CNStageIntLLROutputS7xD(333)(0);
  VNStageIntLLRInputS7xD(106)(5) <= CNStageIntLLROutputS7xD(333)(1);
  VNStageIntLLRInputS7xD(144)(6) <= CNStageIntLLROutputS7xD(333)(2);
  VNStageIntLLRInputS7xD(193)(4) <= CNStageIntLLROutputS7xD(333)(3);
  VNStageIntLLRInputS7xD(261)(5) <= CNStageIntLLROutputS7xD(333)(4);
  VNStageIntLLRInputS7xD(367)(6) <= CNStageIntLLROutputS7xD(333)(5);
  VNStageIntLLRInputS7xD(26)(6) <= CNStageIntLLROutputS7xD(334)(0);
  VNStageIntLLRInputS7xD(126)(5) <= CNStageIntLLROutputS7xD(334)(1);
  VNStageIntLLRInputS7xD(131)(5) <= CNStageIntLLROutputS7xD(334)(2);
  VNStageIntLLRInputS7xD(237)(5) <= CNStageIntLLROutputS7xD(334)(3);
  VNStageIntLLRInputS7xD(277)(6) <= CNStageIntLLROutputS7xD(334)(4);
  VNStageIntLLRInputS7xD(340)(5) <= CNStageIntLLROutputS7xD(334)(5);
  VNStageIntLLRInputS7xD(24)(6) <= CNStageIntLLROutputS7xD(335)(0);
  VNStageIntLLRInputS7xD(107)(5) <= CNStageIntLLROutputS7xD(335)(1);
  VNStageIntLLRInputS7xD(147)(6) <= CNStageIntLLROutputS7xD(335)(2);
  VNStageIntLLRInputS7xD(210)(6) <= CNStageIntLLROutputS7xD(335)(3);
  VNStageIntLLRInputS7xD(300)(5) <= CNStageIntLLROutputS7xD(335)(4);
  VNStageIntLLRInputS7xD(373)(4) <= CNStageIntLLROutputS7xD(335)(5);
  VNStageIntLLRInputS7xD(23)(6) <= CNStageIntLLROutputS7xD(336)(0);
  VNStageIntLLRInputS7xD(82)(6) <= CNStageIntLLROutputS7xD(336)(1);
  VNStageIntLLRInputS7xD(145)(6) <= CNStageIntLLROutputS7xD(336)(2);
  VNStageIntLLRInputS7xD(235)(4) <= CNStageIntLLROutputS7xD(336)(3);
  VNStageIntLLRInputS7xD(308)(4) <= CNStageIntLLROutputS7xD(336)(4);
  VNStageIntLLRInputS7xD(353)(5) <= CNStageIntLLROutputS7xD(336)(5);
  VNStageIntLLRInputS7xD(22)(6) <= CNStageIntLLROutputS7xD(337)(0);
  VNStageIntLLRInputS7xD(80)(5) <= CNStageIntLLROutputS7xD(337)(1);
  VNStageIntLLRInputS7xD(170)(4) <= CNStageIntLLROutputS7xD(337)(2);
  VNStageIntLLRInputS7xD(243)(6) <= CNStageIntLLROutputS7xD(337)(3);
  VNStageIntLLRInputS7xD(288)(6) <= CNStageIntLLROutputS7xD(337)(4);
  VNStageIntLLRInputS7xD(347)(6) <= CNStageIntLLROutputS7xD(337)(5);
  VNStageIntLLRInputS7xD(21)(6) <= CNStageIntLLROutputS7xD(338)(0);
  VNStageIntLLRInputS7xD(105)(5) <= CNStageIntLLROutputS7xD(338)(1);
  VNStageIntLLRInputS7xD(178)(5) <= CNStageIntLLROutputS7xD(338)(2);
  VNStageIntLLRInputS7xD(223)(6) <= CNStageIntLLROutputS7xD(338)(3);
  VNStageIntLLRInputS7xD(282)(5) <= CNStageIntLLROutputS7xD(338)(4);
  VNStageIntLLRInputS7xD(320)(4) <= CNStageIntLLROutputS7xD(338)(5);
  VNStageIntLLRInputS7xD(20)(4) <= CNStageIntLLROutputS7xD(339)(0);
  VNStageIntLLRInputS7xD(113)(6) <= CNStageIntLLROutputS7xD(339)(1);
  VNStageIntLLRInputS7xD(158)(6) <= CNStageIntLLROutputS7xD(339)(2);
  VNStageIntLLRInputS7xD(217)(6) <= CNStageIntLLROutputS7xD(339)(3);
  VNStageIntLLRInputS7xD(256)(5) <= CNStageIntLLROutputS7xD(339)(4);
  VNStageIntLLRInputS7xD(346)(6) <= CNStageIntLLROutputS7xD(339)(5);
  VNStageIntLLRInputS7xD(19)(4) <= CNStageIntLLROutputS7xD(340)(0);
  VNStageIntLLRInputS7xD(93)(6) <= CNStageIntLLROutputS7xD(340)(1);
  VNStageIntLLRInputS7xD(152)(6) <= CNStageIntLLROutputS7xD(340)(2);
  VNStageIntLLRInputS7xD(192)(6) <= CNStageIntLLROutputS7xD(340)(3);
  VNStageIntLLRInputS7xD(281)(6) <= CNStageIntLLROutputS7xD(340)(4);
  VNStageIntLLRInputS7xD(351)(5) <= CNStageIntLLROutputS7xD(340)(5);
  VNStageIntLLRInputS7xD(18)(6) <= CNStageIntLLROutputS7xD(341)(0);
  VNStageIntLLRInputS7xD(87)(6) <= CNStageIntLLROutputS7xD(341)(1);
  VNStageIntLLRInputS7xD(128)(6) <= CNStageIntLLROutputS7xD(341)(2);
  VNStageIntLLRInputS7xD(216)(6) <= CNStageIntLLROutputS7xD(341)(3);
  VNStageIntLLRInputS7xD(286)(6) <= CNStageIntLLROutputS7xD(341)(4);
  VNStageIntLLRInputS7xD(370)(4) <= CNStageIntLLROutputS7xD(341)(5);
  VNStageIntLLRInputS7xD(17)(6) <= CNStageIntLLROutputS7xD(342)(0);
  VNStageIntLLRInputS7xD(64)(5) <= CNStageIntLLROutputS7xD(342)(1);
  VNStageIntLLRInputS7xD(151)(5) <= CNStageIntLLROutputS7xD(342)(2);
  VNStageIntLLRInputS7xD(221)(6) <= CNStageIntLLROutputS7xD(342)(3);
  VNStageIntLLRInputS7xD(305)(6) <= CNStageIntLLROutputS7xD(342)(4);
  VNStageIntLLRInputS7xD(361)(6) <= CNStageIntLLROutputS7xD(342)(5);
  VNStageIntLLRInputS7xD(16)(5) <= CNStageIntLLROutputS7xD(343)(0);
  VNStageIntLLRInputS7xD(86)(3) <= CNStageIntLLROutputS7xD(343)(1);
  VNStageIntLLRInputS7xD(156)(3) <= CNStageIntLLROutputS7xD(343)(2);
  VNStageIntLLRInputS7xD(240)(6) <= CNStageIntLLROutputS7xD(343)(3);
  VNStageIntLLRInputS7xD(296)(5) <= CNStageIntLLROutputS7xD(343)(4);
  VNStageIntLLRInputS7xD(335)(6) <= CNStageIntLLROutputS7xD(343)(5);
  VNStageIntLLRInputS7xD(15)(6) <= CNStageIntLLROutputS7xD(344)(0);
  VNStageIntLLRInputS7xD(91)(6) <= CNStageIntLLROutputS7xD(344)(1);
  VNStageIntLLRInputS7xD(175)(6) <= CNStageIntLLROutputS7xD(344)(2);
  VNStageIntLLRInputS7xD(231)(5) <= CNStageIntLLROutputS7xD(344)(3);
  VNStageIntLLRInputS7xD(270)(6) <= CNStageIntLLROutputS7xD(344)(4);
  VNStageIntLLRInputS7xD(336)(5) <= CNStageIntLLROutputS7xD(344)(5);
  VNStageIntLLRInputS7xD(14)(6) <= CNStageIntLLROutputS7xD(345)(0);
  VNStageIntLLRInputS7xD(110)(6) <= CNStageIntLLROutputS7xD(345)(1);
  VNStageIntLLRInputS7xD(166)(5) <= CNStageIntLLROutputS7xD(345)(2);
  VNStageIntLLRInputS7xD(205)(2) <= CNStageIntLLROutputS7xD(345)(3);
  VNStageIntLLRInputS7xD(271)(5) <= CNStageIntLLROutputS7xD(345)(4);
  VNStageIntLLRInputS7xD(360)(6) <= CNStageIntLLROutputS7xD(345)(5);
  VNStageIntLLRInputS7xD(13)(5) <= CNStageIntLLROutputS7xD(346)(0);
  VNStageIntLLRInputS7xD(101)(6) <= CNStageIntLLROutputS7xD(346)(1);
  VNStageIntLLRInputS7xD(140)(6) <= CNStageIntLLROutputS7xD(346)(2);
  VNStageIntLLRInputS7xD(206)(4) <= CNStageIntLLROutputS7xD(346)(3);
  VNStageIntLLRInputS7xD(295)(4) <= CNStageIntLLROutputS7xD(346)(4);
  VNStageIntLLRInputS7xD(381)(5) <= CNStageIntLLROutputS7xD(346)(5);
  VNStageIntLLRInputS7xD(12)(6) <= CNStageIntLLROutputS7xD(347)(0);
  VNStageIntLLRInputS7xD(75)(6) <= CNStageIntLLROutputS7xD(347)(1);
  VNStageIntLLRInputS7xD(141)(4) <= CNStageIntLLROutputS7xD(347)(2);
  VNStageIntLLRInputS7xD(230)(5) <= CNStageIntLLROutputS7xD(347)(3);
  VNStageIntLLRInputS7xD(316)(4) <= CNStageIntLLROutputS7xD(347)(4);
  VNStageIntLLRInputS7xD(377)(4) <= CNStageIntLLROutputS7xD(347)(5);
  VNStageIntLLRInputS7xD(11)(5) <= CNStageIntLLROutputS7xD(348)(0);
  VNStageIntLLRInputS7xD(76)(6) <= CNStageIntLLROutputS7xD(348)(1);
  VNStageIntLLRInputS7xD(165)(5) <= CNStageIntLLROutputS7xD(348)(2);
  VNStageIntLLRInputS7xD(251)(4) <= CNStageIntLLROutputS7xD(348)(3);
  VNStageIntLLRInputS7xD(312)(5) <= CNStageIntLLROutputS7xD(348)(4);
  VNStageIntLLRInputS7xD(329)(6) <= CNStageIntLLROutputS7xD(348)(5);
  VNStageIntLLRInputS7xD(10)(4) <= CNStageIntLLROutputS7xD(349)(0);
  VNStageIntLLRInputS7xD(100)(6) <= CNStageIntLLROutputS7xD(349)(1);
  VNStageIntLLRInputS7xD(186)(5) <= CNStageIntLLROutputS7xD(349)(2);
  VNStageIntLLRInputS7xD(247)(6) <= CNStageIntLLROutputS7xD(349)(3);
  VNStageIntLLRInputS7xD(264)(6) <= CNStageIntLLROutputS7xD(349)(4);
  VNStageIntLLRInputS7xD(355)(6) <= CNStageIntLLROutputS7xD(349)(5);
  VNStageIntLLRInputS7xD(9)(6) <= CNStageIntLLROutputS7xD(350)(0);
  VNStageIntLLRInputS7xD(121)(5) <= CNStageIntLLROutputS7xD(350)(1);
  VNStageIntLLRInputS7xD(182)(6) <= CNStageIntLLROutputS7xD(350)(2);
  VNStageIntLLRInputS7xD(199)(6) <= CNStageIntLLROutputS7xD(350)(3);
  VNStageIntLLRInputS7xD(290)(5) <= CNStageIntLLROutputS7xD(350)(4);
  VNStageIntLLRInputS7xD(331)(4) <= CNStageIntLLROutputS7xD(350)(5);
  VNStageIntLLRInputS7xD(7)(6) <= CNStageIntLLROutputS7xD(351)(0);
  VNStageIntLLRInputS7xD(69)(6) <= CNStageIntLLROutputS7xD(351)(1);
  VNStageIntLLRInputS7xD(160)(6) <= CNStageIntLLROutputS7xD(351)(2);
  VNStageIntLLRInputS7xD(201)(5) <= CNStageIntLLROutputS7xD(351)(3);
  VNStageIntLLRInputS7xD(298)(6) <= CNStageIntLLROutputS7xD(351)(4);
  VNStageIntLLRInputS7xD(379)(4) <= CNStageIntLLROutputS7xD(351)(5);
  VNStageIntLLRInputS7xD(6)(6) <= CNStageIntLLROutputS7xD(352)(0);
  VNStageIntLLRInputS7xD(95)(6) <= CNStageIntLLROutputS7xD(352)(1);
  VNStageIntLLRInputS7xD(136)(6) <= CNStageIntLLROutputS7xD(352)(2);
  VNStageIntLLRInputS7xD(233)(4) <= CNStageIntLLROutputS7xD(352)(3);
  VNStageIntLLRInputS7xD(314)(3) <= CNStageIntLLROutputS7xD(352)(4);
  VNStageIntLLRInputS7xD(349)(5) <= CNStageIntLLROutputS7xD(352)(5);
  VNStageIntLLRInputS7xD(5)(6) <= CNStageIntLLROutputS7xD(353)(0);
  VNStageIntLLRInputS7xD(71)(5) <= CNStageIntLLROutputS7xD(353)(1);
  VNStageIntLLRInputS7xD(168)(5) <= CNStageIntLLROutputS7xD(353)(2);
  VNStageIntLLRInputS7xD(249)(4) <= CNStageIntLLROutputS7xD(353)(3);
  VNStageIntLLRInputS7xD(284)(6) <= CNStageIntLLROutputS7xD(353)(4);
  VNStageIntLLRInputS7xD(358)(5) <= CNStageIntLLROutputS7xD(353)(5);
  VNStageIntLLRInputS7xD(4)(5) <= CNStageIntLLROutputS7xD(354)(0);
  VNStageIntLLRInputS7xD(103)(6) <= CNStageIntLLROutputS7xD(354)(1);
  VNStageIntLLRInputS7xD(184)(6) <= CNStageIntLLROutputS7xD(354)(2);
  VNStageIntLLRInputS7xD(219)(5) <= CNStageIntLLROutputS7xD(354)(3);
  VNStageIntLLRInputS7xD(293)(5) <= CNStageIntLLROutputS7xD(354)(4);
  VNStageIntLLRInputS7xD(371)(4) <= CNStageIntLLROutputS7xD(354)(5);
  VNStageIntLLRInputS7xD(2)(6) <= CNStageIntLLROutputS7xD(355)(0);
  VNStageIntLLRInputS7xD(89)(5) <= CNStageIntLLROutputS7xD(355)(1);
  VNStageIntLLRInputS7xD(163)(4) <= CNStageIntLLROutputS7xD(355)(2);
  VNStageIntLLRInputS7xD(241)(5) <= CNStageIntLLROutputS7xD(355)(3);
  VNStageIntLLRInputS7xD(285)(6) <= CNStageIntLLROutputS7xD(355)(4);
  VNStageIntLLRInputS7xD(378)(5) <= CNStageIntLLROutputS7xD(355)(5);
  VNStageIntLLRInputS7xD(1)(5) <= CNStageIntLLROutputS7xD(356)(0);
  VNStageIntLLRInputS7xD(98)(5) <= CNStageIntLLROutputS7xD(356)(1);
  VNStageIntLLRInputS7xD(176)(6) <= CNStageIntLLROutputS7xD(356)(2);
  VNStageIntLLRInputS7xD(220)(6) <= CNStageIntLLROutputS7xD(356)(3);
  VNStageIntLLRInputS7xD(313)(3) <= CNStageIntLLROutputS7xD(356)(4);
  VNStageIntLLRInputS7xD(380)(5) <= CNStageIntLLROutputS7xD(356)(5);
  VNStageIntLLRInputS7xD(63)(3) <= CNStageIntLLROutputS7xD(357)(0);
  VNStageIntLLRInputS7xD(111)(6) <= CNStageIntLLROutputS7xD(357)(1);
  VNStageIntLLRInputS7xD(155)(6) <= CNStageIntLLROutputS7xD(357)(2);
  VNStageIntLLRInputS7xD(248)(6) <= CNStageIntLLROutputS7xD(357)(3);
  VNStageIntLLRInputS7xD(315)(5) <= CNStageIntLLROutputS7xD(357)(4);
  VNStageIntLLRInputS7xD(362)(6) <= CNStageIntLLROutputS7xD(357)(5);
  VNStageIntLLRInputS7xD(62)(5) <= CNStageIntLLROutputS7xD(358)(0);
  VNStageIntLLRInputS7xD(90)(6) <= CNStageIntLLROutputS7xD(358)(1);
  VNStageIntLLRInputS7xD(183)(4) <= CNStageIntLLROutputS7xD(358)(2);
  VNStageIntLLRInputS7xD(250)(4) <= CNStageIntLLROutputS7xD(358)(3);
  VNStageIntLLRInputS7xD(297)(6) <= CNStageIntLLROutputS7xD(358)(4);
  VNStageIntLLRInputS7xD(369)(4) <= CNStageIntLLROutputS7xD(358)(5);
  VNStageIntLLRInputS7xD(61)(5) <= CNStageIntLLROutputS7xD(359)(0);
  VNStageIntLLRInputS7xD(118)(5) <= CNStageIntLLROutputS7xD(359)(1);
  VNStageIntLLRInputS7xD(185)(3) <= CNStageIntLLROutputS7xD(359)(2);
  VNStageIntLLRInputS7xD(232)(5) <= CNStageIntLLROutputS7xD(359)(3);
  VNStageIntLLRInputS7xD(304)(6) <= CNStageIntLLROutputS7xD(359)(4);
  VNStageIntLLRInputS7xD(333)(5) <= CNStageIntLLROutputS7xD(359)(5);
  VNStageIntLLRInputS7xD(60)(5) <= CNStageIntLLROutputS7xD(360)(0);
  VNStageIntLLRInputS7xD(120)(3) <= CNStageIntLLROutputS7xD(360)(1);
  VNStageIntLLRInputS7xD(167)(6) <= CNStageIntLLROutputS7xD(360)(2);
  VNStageIntLLRInputS7xD(239)(6) <= CNStageIntLLROutputS7xD(360)(3);
  VNStageIntLLRInputS7xD(268)(6) <= CNStageIntLLROutputS7xD(360)(4);
  VNStageIntLLRInputS7xD(321)(6) <= CNStageIntLLROutputS7xD(360)(5);
  VNStageIntLLRInputS7xD(59)(4) <= CNStageIntLLROutputS7xD(361)(0);
  VNStageIntLLRInputS7xD(102)(5) <= CNStageIntLLROutputS7xD(361)(1);
  VNStageIntLLRInputS7xD(174)(4) <= CNStageIntLLROutputS7xD(361)(2);
  VNStageIntLLRInputS7xD(203)(6) <= CNStageIntLLROutputS7xD(361)(3);
  VNStageIntLLRInputS7xD(319)(6) <= CNStageIntLLROutputS7xD(361)(4);
  VNStageIntLLRInputS7xD(327)(6) <= CNStageIntLLROutputS7xD(361)(5);
  VNStageIntLLRInputS7xD(58)(4) <= CNStageIntLLROutputS7xD(362)(0);
  VNStageIntLLRInputS7xD(109)(5) <= CNStageIntLLROutputS7xD(362)(1);
  VNStageIntLLRInputS7xD(138)(6) <= CNStageIntLLROutputS7xD(362)(2);
  VNStageIntLLRInputS7xD(254)(4) <= CNStageIntLLROutputS7xD(362)(3);
  VNStageIntLLRInputS7xD(262)(5) <= CNStageIntLLROutputS7xD(362)(4);
  VNStageIntLLRInputS7xD(322)(5) <= CNStageIntLLROutputS7xD(362)(5);
  VNStageIntLLRInputS7xD(57)(5) <= CNStageIntLLROutputS7xD(363)(0);
  VNStageIntLLRInputS7xD(73)(5) <= CNStageIntLLROutputS7xD(363)(1);
  VNStageIntLLRInputS7xD(189)(5) <= CNStageIntLLROutputS7xD(363)(2);
  VNStageIntLLRInputS7xD(197)(6) <= CNStageIntLLROutputS7xD(363)(3);
  VNStageIntLLRInputS7xD(257)(6) <= CNStageIntLLROutputS7xD(363)(4);
  VNStageIntLLRInputS7xD(332)(5) <= CNStageIntLLROutputS7xD(363)(5);
  VNStageIntLLRInputS7xD(56)(6) <= CNStageIntLLROutputS7xD(364)(0);
  VNStageIntLLRInputS7xD(124)(4) <= CNStageIntLLROutputS7xD(364)(1);
  VNStageIntLLRInputS7xD(132)(5) <= CNStageIntLLROutputS7xD(364)(2);
  VNStageIntLLRInputS7xD(255)(6) <= CNStageIntLLROutputS7xD(364)(3);
  VNStageIntLLRInputS7xD(267)(6) <= CNStageIntLLROutputS7xD(364)(4);
  VNStageIntLLRInputS7xD(354)(5) <= CNStageIntLLROutputS7xD(364)(5);
  VNStageIntLLRInputS7xD(55)(6) <= CNStageIntLLROutputS7xD(365)(0);
  VNStageIntLLRInputS7xD(67)(3) <= CNStageIntLLROutputS7xD(365)(1);
  VNStageIntLLRInputS7xD(190)(4) <= CNStageIntLLROutputS7xD(365)(2);
  VNStageIntLLRInputS7xD(202)(5) <= CNStageIntLLROutputS7xD(365)(3);
  VNStageIntLLRInputS7xD(289)(6) <= CNStageIntLLROutputS7xD(365)(4);
  VNStageIntLLRInputS7xD(372)(5) <= CNStageIntLLROutputS7xD(365)(5);
  VNStageIntLLRInputS7xD(54)(5) <= CNStageIntLLROutputS7xD(366)(0);
  VNStageIntLLRInputS7xD(125)(3) <= CNStageIntLLROutputS7xD(366)(1);
  VNStageIntLLRInputS7xD(137)(6) <= CNStageIntLLROutputS7xD(366)(2);
  VNStageIntLLRInputS7xD(224)(6) <= CNStageIntLLROutputS7xD(366)(3);
  VNStageIntLLRInputS7xD(307)(6) <= CNStageIntLLROutputS7xD(366)(4);
  VNStageIntLLRInputS7xD(357)(6) <= CNStageIntLLROutputS7xD(366)(5);
  VNStageIntLLRInputS7xD(53)(5) <= CNStageIntLLROutputS7xD(367)(0);
  VNStageIntLLRInputS7xD(72)(5) <= CNStageIntLLROutputS7xD(367)(1);
  VNStageIntLLRInputS7xD(159)(4) <= CNStageIntLLROutputS7xD(367)(2);
  VNStageIntLLRInputS7xD(242)(6) <= CNStageIntLLROutputS7xD(367)(3);
  VNStageIntLLRInputS7xD(292)(6) <= CNStageIntLLROutputS7xD(367)(4);
  VNStageIntLLRInputS7xD(344)(6) <= CNStageIntLLROutputS7xD(367)(5);
  VNStageIntLLRInputS7xD(52)(4) <= CNStageIntLLROutputS7xD(368)(0);
  VNStageIntLLRInputS7xD(94)(4) <= CNStageIntLLROutputS7xD(368)(1);
  VNStageIntLLRInputS7xD(177)(6) <= CNStageIntLLROutputS7xD(368)(2);
  VNStageIntLLRInputS7xD(227)(6) <= CNStageIntLLROutputS7xD(368)(3);
  VNStageIntLLRInputS7xD(279)(5) <= CNStageIntLLROutputS7xD(368)(4);
  VNStageIntLLRInputS7xD(375)(5) <= CNStageIntLLROutputS7xD(368)(5);
  VNStageIntLLRInputS7xD(51)(5) <= CNStageIntLLROutputS7xD(369)(0);
  VNStageIntLLRInputS7xD(112)(6) <= CNStageIntLLROutputS7xD(369)(1);
  VNStageIntLLRInputS7xD(162)(6) <= CNStageIntLLROutputS7xD(369)(2);
  VNStageIntLLRInputS7xD(214)(6) <= CNStageIntLLROutputS7xD(369)(3);
  VNStageIntLLRInputS7xD(310)(5) <= CNStageIntLLROutputS7xD(369)(4);
  VNStageIntLLRInputS7xD(324)(6) <= CNStageIntLLROutputS7xD(369)(5);
  VNStageIntLLRInputS7xD(50)(6) <= CNStageIntLLROutputS7xD(370)(0);
  VNStageIntLLRInputS7xD(97)(6) <= CNStageIntLLROutputS7xD(370)(1);
  VNStageIntLLRInputS7xD(149)(6) <= CNStageIntLLROutputS7xD(370)(2);
  VNStageIntLLRInputS7xD(245)(6) <= CNStageIntLLROutputS7xD(370)(3);
  VNStageIntLLRInputS7xD(259)(4) <= CNStageIntLLROutputS7xD(370)(4);
  VNStageIntLLRInputS7xD(338)(4) <= CNStageIntLLROutputS7xD(370)(5);
  VNStageIntLLRInputS7xD(49)(6) <= CNStageIntLLROutputS7xD(371)(0);
  VNStageIntLLRInputS7xD(84)(5) <= CNStageIntLLROutputS7xD(371)(1);
  VNStageIntLLRInputS7xD(180)(4) <= CNStageIntLLROutputS7xD(371)(2);
  VNStageIntLLRInputS7xD(194)(6) <= CNStageIntLLROutputS7xD(371)(3);
  VNStageIntLLRInputS7xD(273)(5) <= CNStageIntLLROutputS7xD(371)(4);
  VNStageIntLLRInputS7xD(382)(5) <= CNStageIntLLROutputS7xD(371)(5);
  VNStageIntLLRInputS7xD(48)(3) <= CNStageIntLLROutputS7xD(372)(0);
  VNStageIntLLRInputS7xD(115)(6) <= CNStageIntLLROutputS7xD(372)(1);
  VNStageIntLLRInputS7xD(129)(6) <= CNStageIntLLROutputS7xD(372)(2);
  VNStageIntLLRInputS7xD(208)(5) <= CNStageIntLLROutputS7xD(372)(3);
  VNStageIntLLRInputS7xD(317)(3) <= CNStageIntLLROutputS7xD(372)(4);
  VNStageIntLLRInputS7xD(359)(6) <= CNStageIntLLROutputS7xD(372)(5);
  VNStageIntLLRInputS7xD(47)(3) <= CNStageIntLLROutputS7xD(373)(0);
  VNStageIntLLRInputS7xD(127)(6) <= CNStageIntLLROutputS7xD(373)(1);
  VNStageIntLLRInputS7xD(143)(6) <= CNStageIntLLROutputS7xD(373)(2);
  VNStageIntLLRInputS7xD(252)(5) <= CNStageIntLLROutputS7xD(373)(3);
  VNStageIntLLRInputS7xD(294)(6) <= CNStageIntLLROutputS7xD(373)(4);
  VNStageIntLLRInputS7xD(348)(6) <= CNStageIntLLROutputS7xD(373)(5);
  VNStageIntLLRInputS7xD(46)(6) <= CNStageIntLLROutputS7xD(374)(0);
  VNStageIntLLRInputS7xD(78)(6) <= CNStageIntLLROutputS7xD(374)(1);
  VNStageIntLLRInputS7xD(187)(5) <= CNStageIntLLROutputS7xD(374)(2);
  VNStageIntLLRInputS7xD(229)(4) <= CNStageIntLLROutputS7xD(374)(3);
  VNStageIntLLRInputS7xD(283)(6) <= CNStageIntLLROutputS7xD(374)(4);
  VNStageIntLLRInputS7xD(352)(6) <= CNStageIntLLROutputS7xD(374)(5);
  VNStageIntLLRInputS7xD(45)(6) <= CNStageIntLLROutputS7xD(375)(0);
  VNStageIntLLRInputS7xD(122)(5) <= CNStageIntLLROutputS7xD(375)(1);
  VNStageIntLLRInputS7xD(164)(5) <= CNStageIntLLROutputS7xD(375)(2);
  VNStageIntLLRInputS7xD(218)(6) <= CNStageIntLLROutputS7xD(375)(3);
  VNStageIntLLRInputS7xD(287)(6) <= CNStageIntLLROutputS7xD(375)(4);
  VNStageIntLLRInputS7xD(345)(5) <= CNStageIntLLROutputS7xD(375)(5);
  VNStageIntLLRInputS7xD(44)(6) <= CNStageIntLLROutputS7xD(376)(0);
  VNStageIntLLRInputS7xD(99)(6) <= CNStageIntLLROutputS7xD(376)(1);
  VNStageIntLLRInputS7xD(153)(6) <= CNStageIntLLROutputS7xD(376)(2);
  VNStageIntLLRInputS7xD(222)(3) <= CNStageIntLLROutputS7xD(376)(3);
  VNStageIntLLRInputS7xD(280)(6) <= CNStageIntLLROutputS7xD(376)(4);
  VNStageIntLLRInputS7xD(356)(5) <= CNStageIntLLROutputS7xD(376)(5);
  VNStageIntLLRInputS7xD(43)(5) <= CNStageIntLLROutputS7xD(377)(0);
  VNStageIntLLRInputS7xD(88)(6) <= CNStageIntLLROutputS7xD(377)(1);
  VNStageIntLLRInputS7xD(157)(5) <= CNStageIntLLROutputS7xD(377)(2);
  VNStageIntLLRInputS7xD(215)(6) <= CNStageIntLLROutputS7xD(377)(3);
  VNStageIntLLRInputS7xD(291)(5) <= CNStageIntLLROutputS7xD(377)(4);
  VNStageIntLLRInputS7xD(328)(4) <= CNStageIntLLROutputS7xD(377)(5);
  VNStageIntLLRInputS7xD(42)(6) <= CNStageIntLLROutputS7xD(378)(0);
  VNStageIntLLRInputS7xD(92)(6) <= CNStageIntLLROutputS7xD(378)(1);
  VNStageIntLLRInputS7xD(150)(5) <= CNStageIntLLROutputS7xD(378)(2);
  VNStageIntLLRInputS7xD(226)(2) <= CNStageIntLLROutputS7xD(378)(3);
  VNStageIntLLRInputS7xD(263)(6) <= CNStageIntLLROutputS7xD(378)(4);
  VNStageIntLLRInputS7xD(383)(6) <= CNStageIntLLROutputS7xD(378)(5);
  VNStageIntLLRInputS7xD(41)(6) <= CNStageIntLLROutputS7xD(379)(0);
  VNStageIntLLRInputS7xD(85)(5) <= CNStageIntLLROutputS7xD(379)(1);
  VNStageIntLLRInputS7xD(161)(6) <= CNStageIntLLROutputS7xD(379)(2);
  VNStageIntLLRInputS7xD(198)(6) <= CNStageIntLLROutputS7xD(379)(3);
  VNStageIntLLRInputS7xD(318)(3) <= CNStageIntLLROutputS7xD(379)(4);
  VNStageIntLLRInputS7xD(337)(6) <= CNStageIntLLROutputS7xD(379)(5);
  VNStageIntLLRInputS7xD(40)(4) <= CNStageIntLLROutputS7xD(380)(0);
  VNStageIntLLRInputS7xD(96)(5) <= CNStageIntLLROutputS7xD(380)(1);
  VNStageIntLLRInputS7xD(133)(4) <= CNStageIntLLROutputS7xD(380)(2);
  VNStageIntLLRInputS7xD(253)(5) <= CNStageIntLLROutputS7xD(380)(3);
  VNStageIntLLRInputS7xD(272)(6) <= CNStageIntLLROutputS7xD(380)(4);
  VNStageIntLLRInputS7xD(334)(4) <= CNStageIntLLROutputS7xD(380)(5);
  VNStageIntLLRInputS7xD(39)(6) <= CNStageIntLLROutputS7xD(381)(0);
  VNStageIntLLRInputS7xD(68)(5) <= CNStageIntLLROutputS7xD(381)(1);
  VNStageIntLLRInputS7xD(188)(4) <= CNStageIntLLROutputS7xD(381)(2);
  VNStageIntLLRInputS7xD(207)(5) <= CNStageIntLLROutputS7xD(381)(3);
  VNStageIntLLRInputS7xD(269)(5) <= CNStageIntLLROutputS7xD(381)(4);
  VNStageIntLLRInputS7xD(368)(2) <= CNStageIntLLROutputS7xD(381)(5);
  VNStageIntLLRInputS7xD(38)(6) <= CNStageIntLLROutputS7xD(382)(0);
  VNStageIntLLRInputS7xD(123)(4) <= CNStageIntLLROutputS7xD(382)(1);
  VNStageIntLLRInputS7xD(142)(4) <= CNStageIntLLROutputS7xD(382)(2);
  VNStageIntLLRInputS7xD(204)(6) <= CNStageIntLLROutputS7xD(382)(3);
  VNStageIntLLRInputS7xD(303)(6) <= CNStageIntLLROutputS7xD(382)(4);
  VNStageIntLLRInputS7xD(325)(6) <= CNStageIntLLROutputS7xD(382)(5);
  VNStageIntLLRInputS7xD(37)(6) <= CNStageIntLLROutputS7xD(383)(0);
  VNStageIntLLRInputS7xD(77)(4) <= CNStageIntLLROutputS7xD(383)(1);
  VNStageIntLLRInputS7xD(139)(6) <= CNStageIntLLROutputS7xD(383)(2);
  VNStageIntLLRInputS7xD(238)(6) <= CNStageIntLLROutputS7xD(383)(3);
  VNStageIntLLRInputS7xD(260)(5) <= CNStageIntLLROutputS7xD(383)(4);
  VNStageIntLLRInputS7xD(374)(6) <= CNStageIntLLROutputS7xD(383)(5);

  -- Connect output of last VN stage with top-level output
  DecodedBitsxDO <= VNStageIntLLROutputS7xD;

end arch;